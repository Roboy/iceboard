// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Tue Feb  4 18:20:54 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, INLC_c_0, INHC_c_0, 
        INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire h1, h2, h3;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(116[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(117[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(126[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(223[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(225[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(226[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(227[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(228[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(229[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(231[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(232[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(233[22:35])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(263[22:33])
    wire [7:0]data;   // verilog/TinyFPGA_B.v(326[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(350[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(358[15:20])
    
    wire pwm_setpoint_23__N_215;
    wire [23:0]pwm_setpoint_23__N_191;
    wire [23:0]pwm_setpoint_23__N_11;
    wire [7:0]commutation_state_7__N_216;
    
    wire commutation_state_7__N_224;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(222[11:28])
    
    wire n861, GHA_N_367, GLA_N_384, GHB_N_389, GLB_N_398, GHC_N_403, 
        GLC_N_412, dti_N_416, RX_N_10, n1617;
    wire [31:0]motor_state_23__N_123;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_279;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
        n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
        n1195, n39429, n516, n7, n14, n1658;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(224[11:28])
    
    wire n4;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n833, n832, n831, n830, n829, n828;
    wire [3:0]state_3__N_528;
    
    wire n4_adj_5091, n3, n39428, n2, n6935, n39427, n10, n48697, 
        n6662, n48696, n10_adj_5092, n39426, n731, n39425, n29756, 
        n4_adj_5093, n29755, n49900, n29754, n29753, n29752, n29751, 
        n39143, n29750, n29749, n29748, n39597, n39596, n39595, 
        n39594, n29747, n39593, n29746, n29745, n29744, n29743, 
        n39592, n29742, n29741, n39591, n39590, n36109, n7355, 
        n7354, n7353, n7352, n7351, n29740, n29739, n35141, n4_adj_5094, 
        n29738;
    wire [2:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n29737, n29736, n3_adj_5095, n4_adj_5096, n5, n6, n7_adj_5097, 
        n8, n9, n10_adj_5098, n11, n12, n13, n14_adj_5099, n15, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n50883;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    
    wire n12_adj_5100;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n21743, n123, n50401;
    wire [31:0]\FRAME_MATCHER.state_31__N_2660 ;
    
    wire n39142, n45257, n51286, n43275, n29735, n29734, n771, 
        n4_adj_5101, n15_adj_5102, n14_adj_5103, n44068, n39141, n39140, 
        n45167, n39075, n45172, n39139, n36411, n51252, n39138, 
        n39137, n36395, n36393, n39074, n39136, n40581, n40582, 
        n39135, n40583, n40584, n39134, n40586, n40587, n40588, 
        n40589, n36369, n40590, n39133, n36365, n39132, n40578, 
        n40574, n45246, n36407, n45183, n43841, n45214, n45252, 
        n40383, n36307, n40382, n40381, n36299, n40380, n36303, 
        n40379, n40378, n40377, n36297, n45275, n35282, n29733, 
        n40560, n40368, n40367, n2_adj_5104, n29732, n29731, n44866, 
        n29730, n29729, n27826, n40366, n3303, n40561, n40914, 
        n40365, n40562, n40913, n40364, n40363, n40563, n40912, 
        n40911, n40564, n40575, n40910, n40565, n40576, n40362, 
        n40566, n40567, n40568, n40569, n40579, n40361, n40360, 
        n40570, n40571, n40580, n40359, n40572, n40573, n39131, 
        n40358, n39371, n40357, n40356, n40355, n40354, n29728, 
        n29727, n4452, n40353, n39370, n39091, n39369, n40352, 
        n39368, n40351, n39367, n5_adj_5105, n40350, n40349, n82, 
        n40348, n40347, n40346, n40345, n40344, n40343, n39366, 
        n39365, n39364, n40342, n40341, n40340, n40339, n40338, 
        n40337, n39363, n39130, n39362, n40336, n40335, n40334, 
        n40333, n40332, n40331, n40330, n40329, n40328, n39361, 
        n39360, n39359, n39358, n40327, n40326, n36301, n39357, 
        n39356, n40325, n40324, n51668, n29724, n29723, n40323, 
        n40322, n40321, n40320, n39355, n29722, n29721, n40319, 
        n29720, n29719, \FRAME_MATCHER.i_31__N_2622 , \FRAME_MATCHER.i_31__N_2624 , 
        \FRAME_MATCHER.i_31__N_2626 , n14_adj_5106, n44859, n43061, 
        n10_adj_5107, n45250, n36235, n40318, n40317, n40316, n40315, 
        n40314, n40313, n40312, n40311, n40310, n40309, n40308, 
        n40307, n40306, n40305, n40304, n40303, n40302, n40301, 
        n40300, n40299, n40298, n40297, n40296, n40295, n40294, 
        n40293, n40292, n40291, n40290, n40289, n40288, n40287, 
        n40286, n40285, n40284, n40283, n40282, n40281, n40280, 
        n40279, n40278, n40277, n40276, n40275, n40274, n40273, 
        n40272, n40271, n40270, n40269, n40268, n40267, n40266, 
        n40265, n40264, n40263, n40262, n40261, n40260, n40259, 
        n40258, n40257, n40256, n40255, n40254, n40253, n40252, 
        n40251, n40250, n39090, n40249, n39354, n40248, n40247, 
        n40246, n39129, n652, n628, n627, n625, n623, n622, 
        n621, n30212, n40245, n40244, n40243, n30209, n40242, 
        n40241, n39353, n45643, n48576, n5_adj_5108, n30208, n30207, 
        n25_adj_5109, n24_adj_5110, n23_adj_5111, n22_adj_5112, n21_adj_5113, 
        n20_adj_5114, n19_adj_5115, n18_adj_5116, n17_adj_5117, n16_adj_5118, 
        n29718, n29717, n29716, n29715, n29714, n29713, n29712, 
        n29711, n29710, n29709, n29708, n29707, n29706, n29705, 
        n29704, n29703, n15_adj_5119, n14_adj_5120, n13_adj_5121, 
        n12_adj_5122, n11_adj_5123, n10_adj_5124, n9_adj_5125, n39352, 
        n40240, n39351, n40239, n40238, n40237, n40236, n30206, 
        n30205, n30204, n40235, n8_adj_5126, n7_adj_5127, n6_adj_5128, 
        n5_adj_5129, n4_adj_5130, n3_adj_5131, n5741, n51219, n30203, 
        n30202, n30201, n30200, n30199, n40234, n30198, n29702, 
        n30197, n30196, n30195, n40233, n30194, n40232, n40231, 
        n30193, n29701, n40230, n40229, n40228, n15_adj_5132, n30192, 
        n40227, n30191, n30190, n30189, n40226, n40225, n30188, 
        n40224, n30186, n30185, n30184, n30183, n40223, n40222, 
        n40221, n30182, n30181, n30180, n30179, n30178, n40220, 
        n30177, n30176, n30175, n30174, n30173, n30172, n30171;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n40219, n27828, n30170, n30169, n30168, n30167, 
        n30166, n30165, n40218, n30164, n40217, n4_adj_5133, n30163, 
        n30162, n30161, n30160, n30159, n40216, direction_N_3907, 
        n30158, n30157, n30156, n30155, n40215, n30154, n30153, 
        n30152, n30151, n30150, n30149, n30148, n30147, n30146, 
        n30145, n40214, n30144, n40213, n40212, n15_adj_5134, n40211, 
        n30143, n30141, n40210, n40209, n40208, n40207, n40206, 
        n39128, n40205, n30140, n40204, n30139, n30138;
    wire [1:0]a_new_adj_5265;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_5136, n40203, n40202, n30137, n30136, n30135, 
        n30134, n1910, n30133, n30132, n30131, n30130, n30129, 
        n40201, n30128, n30127, n30126, n30125, n30124, n40200, 
        n30123, n40199, n30122, n30121, direction_N_3907_adj_5137, 
        n40198, n30120, n30119, n30118, n30117, n7350, n30116, 
        n30115, n30114, n30113, n30112, n30111, n30110, n30109, 
        n40197, n30108, n30107, n30106, n30105, n43733, n30104, 
        n30103, n30102, n30101, n30100, n30099, n30098, n30097, 
        n30096, n40196, n40195, n40194, n40193, n30095, n30094, 
        n30093, n30092, n30091, n30090, n30089, n30088, n30087, 
        n30086, n4_adj_5138, n30085, n33, rw;
    wire [7:0]state_adj_5289;   // verilog/eeprom.v(23[11:16])
    
    wire n40192, n32, n31, n30, n29, n28, n27, n26, n25_adj_5141, 
        n24_adj_5142, n23_adj_5143, n22_adj_5144, n21_adj_5145, n20_adj_5146, 
        n19_adj_5147, n18_adj_5148, n17_adj_5149, n30084, n30083, 
        n30082, n30081, n30080, n30079, n40191, n30078, n30077, 
        n30076, n40190, n5_adj_5150, n30075, n30074, n30073, n30072, 
        n30071, n30070, n30069, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n40189, n16_adj_5151, n4_adj_5152, n15_adj_5153, n30068, 
        n30067, n30066, n30065, n30064, n30063, n30062, n30061, 
        n30060, n40188, n40187, n39127, n40186, n40185, n30059, 
        n30058, n40184, n40183, n40182, n14_adj_5154, n30057, n13_adj_5155, 
        n30056, n12_adj_5156, n11_adj_5157;
    wire [2:0]r_SM_Main_2__N_3542;
    
    wire n39126, n30055, n30054, n30053, n29700, n45229, n8_adj_5158, 
        n30052, n40181, n30051, n30050, n30049, n30048, n30047, 
        n30046, n30045, n30044, n30043, n30042, n30041, n30040, 
        n30039, n30038, n30037;
    wire [2:0]r_SM_Main_adj_5298;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5300;   // verilog/uart_tx.v(33[16:27])
    
    wire n40180, n40179, n40178, n40177, n40176, n40175;
    wire [2:0]r_SM_Main_2__N_3613;
    
    wire n40174, n40173, n30036, n30035, n40172, n30034, n30033, 
        n40171, n40170, n30032, n30031, n30030, n30029, n30028, 
        n30027, n30026, n30025, n30024, n30023, n30022, n30021, 
        n30020, n30019, n30018, n30017, n30016, n30015, n30014, 
        n30013, n30012, n30011, n29699;
    wire [7:0]state_adj_5307;   // verilog/i2c_controller.v(33[12:17])
    
    wire n30009, n40169, n30008;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n30007, n30006, n30005, n40168, n30004, n40167, enable_slow_N_4190, 
        n6_adj_5164, n40166, n40165, n40164, n40163, n40162, n40161, 
        n30003, n40160, n30002, n40159, n30001, n40158, n40157, 
        n40156;
    wire [7:0]state_7__N_4087;
    
    wire n30000, n29999, n29698, n6387, n29998, n29997, n29996, 
        n29995, n29994, n29993, n29992, n29991, n29990;
    wire [7:0]state_7__N_4103;
    
    wire n29989, n29988, n29987, n29986, n29985, n29984, n29983, 
        n29982, n39350, n40577, n29981, n29980, n29979, n29978, 
        n29977, n29697, n29696, n29695, n29694, n29693, n29692, 
        n10_adj_5165, n6969, n29976, n29975, n29974, n29973, n29972, 
        n29323, n29971, n29970, n28004, n29969, n29968, n29967, 
        n29966, n29965, n29964, n29963, n29962, n29961, n29960, 
        n29959, n29958, n29957, n29956, n29955, n29954, n29953, 
        n29952, n29951, n29950, n29949, n29948, n29947, n29310, 
        n9_adj_5166, n29946, n8_adj_5167, n29945, n29944, n29943, 
        n29942, n29941, n29940, n29939, n29938, n896, n897, n898, 
        n899, n900, n901, n927, n928, n929, n930, n931, n932, 
        n933, n935, n936, n937, n938, n939, n940, n941, n942, 
        n943, n944, n945, n946, n947, n948, n949, n950, n951, 
        n952, n953, n954, n955, n956, n957, n960, n995, n996, 
        n997, n998, n999, n1000, n1001, n1026, n1027, n1028, 
        n1029, n1030, n1031, n1032, n1033, n1059, n1093_adj_5168, 
        n1094_adj_5169, n1095_adj_5170, n1096_adj_5171, n1097_adj_5172, 
        n1098_adj_5173, n1099_adj_5174, n1100_adj_5175, n1101_adj_5176, 
        n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
        n1133, n1158, n1193, n1194, n1195_adj_5177, n1196, n1197, 
        n1198, n1199, n1200, n1201, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1257, n1292, 
        n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, 
        n1301, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
        n1330, n1331, n1332, n1333, n1356, n1391, n1392, n1393, 
        n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
        n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
        n1430, n1431, n1432, n1433, n1455, n1490, n1491, n1492, 
        n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
        n1501, n29937, n1521, n1522, n1523, n1524, n1525, n1526, 
        n1527, n1528, n1529, n1530, n1531, n1532, n1533, n29257, 
        n1554, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
        n1596, n1597, n1598, n1599, n1600, n1601, n1620, n1621, 
        n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
        n1630, n1631, n1632, n1633, n1653_adj_5178, n1688, n1689, 
        n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
        n1698, n1699, n1700, n1701, n29246, n1719, n1720, n1721, 
        n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
        n1730, n1731, n1732, n1733, n29936, n29234, n50892, n1752, 
        n29935, n1787, n1788, n1789, n1790, n1791, n1792, n1793, 
        n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
        n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
        n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
        n29934, n1851, n29208, n1886, n1887, n1888, n1889, n1890, 
        n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
        n1899, n1900, n1901, n29933, n1917, n1918, n1919, n1920, 
        n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
        n1929, n1930, n1931, n1932, n1933, n39125, n1950, n29932, 
        n29533, n1985, n1986, n1987, n1988, n1989, n1990, n1991, 
        n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
        n2000, n2001, n2016, n2017, n2018, n2019, n2020, n2021, 
        n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
        n2030, n2031, n2032, n2033, n29176, n2049, n29689, n2084, 
        n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
        n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, 
        n2101, n2115, n2116, n2117, n2118, n2119, n2120, n2121, 
        n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
        n2130, n2131, n2132, n2133, n2148, n25336, n2183, n2184, 
        n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
        n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, 
        n2201, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
        n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, 
        n2229, n2230, n2231, n2232, n2233, n2247, n29460, n7_adj_5179, 
        n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
        n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, 
        n2298, n2299, n2300, n2301, n2313, n2314, n2315, n2316, 
        n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
        n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
        n2333, n2346, n29125, n2381, n2382, n2383, n2384, n2385, 
        n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
        n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, 
        n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
        n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, 
        n2428, n2429, n2430, n2431, n2432, n2433, n51071, n2445, 
        n29117, n2480, n2481, n2482, n2483, n2484, n2485, n2486, 
        n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
        n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2511, 
        n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
        n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, 
        n2528, n2529, n2530, n2531, n2532, n2533, n2544, n2579, 
        n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
        n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, 
        n2596, n2597, n2598, n2599, n2600, n2601, n2610, n2611, 
        n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
        n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, 
        n2628, n2629, n2630, n2631, n2632, n2633, n2643, n2677, 
        n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, 
        n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, 
        n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
        n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, 
        n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
        n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, 
        n2733, n2742, n51594, n2777, n2778, n2779, n2780, n2781, 
        n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, 
        n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, 
        n2798, n2799, n2800, n2801, n2808, n2809, n2810, n2811, 
        n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
        n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, 
        n2828, n2829, n2830, n2831, n2832, n2833, n2841, n2876, 
        n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
        n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
        n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
        n2901, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
        n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
        n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
        n2930, n2931, n2932, n2933, n2940, n2975, n2976, n2977, 
        n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, 
        n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
        n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
        n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
        n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
        n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
        n3030, n3031, n3032, n3033, n3039, n3073, n3074, n3075, 
        n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
        n3100, n3101, n3105, n3106, n3107, n3108, n3109, n3110, 
        n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
        n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
        n3127, n3128, n3129, n3130, n3131, n3132, n3133, n51290, 
        n3138, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
        n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, 
        n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, 
        n3196, n3197, n3198, n3199, n3200, n3201, n3204, n3205, 
        n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
        n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
        n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
        n3230, n3231, n3232, n3233, n51324, n3237, n3272, n3273, 
        n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
        n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
        n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3298, 
        n3299, n3300, n3301, n6_adj_5180, n51593, n51187, n8_adj_5181, 
        n24_adj_5182, n7_adj_5183, n62, n45266, n27858, n27861, 
        n44138, n50760, n48682, n7_adj_5184, n63, n1, n27984, 
        n29684, n47744, n29679, n47736, n47730, n39073, n50863, 
        n47724, n36277, n47718, n47712, n47708, n47706, n47696, 
        n47690, n48, n49, n50, n51, n52, n53, n54, n55, n7_adj_5185, 
        n47684, n46806, n51153, n47676, n47670, n40055, n27996, 
        n47664, n40054, n47660, n6_adj_5186, n47658, n40053, n40052, 
        n40051, n40050, n40049, n29675, n29674, n29672, n29667, 
        n29664, n29663, n29662, n29661, n46745, n29658, n29657, 
        n29655, n29654, n29653, n29652, n29650, n29649, n29648, 
        n29647, n29646, n40048, n40047, n40046, n50164, n40045, 
        n51124, n48680, n40044, n29645, n29644, n46068, n40043, 
        n29633, n29631, n29630, n29629, n39124, n45319, n35422, 
        n40042, n40041, n40040, n40039, n40038, n40037, n40036, 
        n40035, n40034, n40033, n5_adj_5187, n47640, n47634, n2_adj_5188, 
        n3_adj_5189, n4_adj_5190, n5_adj_5191, n6_adj_5192, n7_adj_5193, 
        n8_adj_5194, n9_adj_5195, n10_adj_5196, n11_adj_5197, n12_adj_5198, 
        n13_adj_5199, n14_adj_5200, n15_adj_5201, n16_adj_5202, n17_adj_5203, 
        n18_adj_5204, n19_adj_5205, n20_adj_5206, n21_adj_5207, n22_adj_5208, 
        n23_adj_5209, n24_adj_5210, n25_adj_5211, n26_adj_5212, n27_adj_5213, 
        n28_adj_5214, n29_adj_5215, n30_adj_5216, n31_adj_5217, n32_adj_5218, 
        n33_adj_5219, n43957, n36379, n47628, n47626, n39123, n7_adj_5220, 
        n4_adj_5221, n50840, n36227, n47620, n39349, n36329, n39936, 
        n39935, n39934, n39933, n39932, n36223, n39931, n47616, 
        n47614, n39930, n39929, n39928, n36337, n39927, n39926, 
        n39925, n36325, n39924, n39923, n39922, n39921, n39920, 
        n39919, n39918, n39072, n39917, n39916, n39915, n39089, 
        n39088, n47602, n39903, n39122, n39902, n39901, n39900, 
        n39899, n39898, n39897, n39896, n39121, n36211, n39895, 
        n39894, n39893, n39892, n39891, n39890, n39889, n39120, 
        n47596, n47594, n10_adj_5222, n39888, n39887, n39886, n39885, 
        n39119, n39884, n36311, n39883, n35414, n47588, n36205, 
        n47582, n36203, n39872, n39871, n39870, n39869, n39868, 
        n39071, n47576, n47574, n50822, n39867, n39866, n39865, 
        n39864, n39863, n47566, n39862, n39861, n39860, n39859, 
        n47558, n39858, n39118, n39117, n39857, n39856, n39855, 
        n39854, n39853, n39852, n47552, n39851, n39850, n39849, 
        n39848, n39847, n39846, n39845, n39844, n39843, n36201, 
        n39842, n45315, n39841, n39840, n39839, n39838, n39837, 
        n39116, n47546, n39836, n39835, n39115, n39114, n47542, 
        n39834, n39833, n39832, n39831, n39113, n39830, n39112, 
        n19_adj_5223, n21_adj_5224, n23_adj_5225, n25_adj_5226, n27_adj_5227, 
        n29_adj_5228, n37, n41, n59, n61, n39829, n39828, n39827, 
        n39826, n39825, n39824, n39823, n39822, n39821, n47530, 
        n39820, n45164, n39087, n47524, n46565, n47520, n47514, 
        n39819, n47512, n39818, n39817, n39816, n39815, n47494, 
        n39814, n47488, n20400, n49702, n47482, n39813, n47478, 
        n44919, n14_adj_5229, n51067, n47474, n43483, n39812, n39811, 
        n39086, n45660, n39085, n29623, n39810, n39809, n39808, 
        n39807, n39806, n47464, n39805, n44909, n27971, n39804, 
        n47458, n47454, n39803, n44888, n44886, n50805, n44880, 
        n47440, n39802, n49682, n51039, n44868, n49681, n44865, 
        n47434, n47428, n49680, n49679, n39801, n39800, n49678, 
        n47416, n25063, n49677, n39799, n47410, n49676, n47400, 
        n47392, n47386, n47376, n4_adj_5230, n39798, n39797, n39796, 
        n39795, n47366, n47360, n47356, n39794, n39793, n39084, 
        n39111, n51013, n47350, n47348, n39792, n39791, n39790, 
        n39083, n39789, n39788, n39787, n39786, n39785, n39784, 
        n39783, n39782, n39781, n39780, n39779, n46975, n39778, 
        n39777, n39776, n39775, n39774, n39773, n39772, n39771, 
        n39770, n39769, n39768, n39767, n39766, n39765, n39764, 
        n39763, n39762, n39761, n39760, n39759, n39758, n39757, 
        n39756, n39755, n39754, n39753, n39752, n39751, n39750, 
        n39749, n39748, n39747, n39746, n39745, n39744, n39743, 
        n39742, n39741, n39740, n39739, n39738, n39737, n39736, 
        n39735, n39734, n39733, n39732, n46973, n39731, n39730, 
        n39729, n47336, n50987, n39718, n39717, n39716, n39715, 
        n39714, n39713, n39712, n39711, n39710, n39709, n39708, 
        n47326, n47320, n39707, n39706, n39705, n39704, n39082, 
        n47314, n29628, n29627, n45880, n47308, n29626, n47302, 
        n29625, n47300, n29624, n47298, n39703, n39144, n39702, 
        n49662, n50789, n46694, n47280, n47274, n39701, n39700, 
        n39699, n39698, n47268, n39697, n39696, n39695, n39694, 
        n39693, n39692, n39691, n39110, n39690, n39109, n39108, 
        n39689, n39107, n47258, n39070, n47252, n47246, n50961, 
        n47240, n47236, n47234, n39106, n47222, n39105, n39104, 
        n4_adj_5231, n47214, n27976, n39081, n27855, n39103, n47208, 
        n47206, n39102, n39080, n47200, n47198, n47188, n39079, 
        n47182, n39101, n36149, n46952, n39078, n41916, n39100, 
        n39069, n47176, n50935, n39077, n39099, n39098, n47170, 
        n39068, n47166, n47162, n39447, n36141, n47152, n39446, 
        n39445, n40585, n39444, n39443, n46788, n25135, n47146, 
        n47142, n39097, n39442, n39441, n47130, n47128, n47122, 
        n44059, n47116, n39096, n39095, n47114, n47112, n39094, 
        n47110, n47108, n47106, n47104, n47102, n36389, n39076, 
        n39093, n47100, n47096, n47094, n39092, n45192, n47090, 
        n47082, n47080, n36493, n47078, n49621, n47076, n47074, 
        n27827, n47072, n50774, n35178, n47066, n47062, n47056, 
        n39430;
    
    VCC i2 (.Y(VCC_net));
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF dir_175 (.Q(dir), .C(CLK_c), .D(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 i16553_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n25135), .I3(GND_net), .O(n30080));   // verilog/coms.v(127[12] 300[6])
    defparam i16553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16554_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n25135), .I3(GND_net), .O(n30081));   // verilog/coms.v(127[12] 300[6])
    defparam i16554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16555_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n25135), .I3(GND_net), .O(n30082));   // verilog/coms.v(127[12] 300[6])
    defparam i16555_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n39865), .I0(n2221), 
            .I1(VCC_net), .CO(n39866));
    SB_LUT4 unary_minus_10_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_DFFE dti_177 (.Q(dti), .C(CLK_c), .E(n29117), .D(dti_N_416));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n39863), .I0(n2223), 
            .I1(VCC_net), .CO(n39864));
    SB_LUT4 i16556_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n25135), .I3(GND_net), .O(n30083));   // verilog/coms.v(127[12] 300[6])
    defparam i16556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16178_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n43061), .I3(GND_net), .O(n29705));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16178_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n40157), .I0(n2632), 
            .I1(GND_net), .CO(n40158));
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n39862), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n40309), .I0(n3110), 
            .I1(VCC_net), .CO(n40310));
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n40156), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n40156), .I0(n2633), 
            .I1(VCC_net), .CO(n40157));
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n39865), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16557_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n25135), .I3(GND_net), .O(n30084));   // verilog/coms.v(127[12] 300[6])
    defparam i16557_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n39862), .I0(n2224), 
            .I1(VCC_net), .CO(n39863));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n39861), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16558_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n25135), .I3(GND_net), .O(n30085));   // verilog/coms.v(127[12] 300[6])
    defparam i16558_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n40156));
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n39861), .I0(n2225), 
            .I1(VCC_net), .CO(n39862));
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16559_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n25135), .I3(GND_net), .O(n30086));   // verilog/coms.v(127[12] 300[6])
    defparam i16559_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_23__N_11[0]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4103[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i16179_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n43061), .I3(GND_net), .O(n29706));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n39860), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_10_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n39860), .I0(n2226), 
            .I1(VCC_net), .CO(n39861));
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.GND_net(GND_net), .CLK_c(CLK_c), 
            .VCC_net(VCC_net), .\state[0] (state[0]), .\state[1] (state[1]), 
            .n43061(n43061), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .n29724(n29724), .n29723(n29723), .n29722(n29722), .n29721(n29721), 
            .n29720(n29720), .n29719(n29719), .n29718(n29718), .n29717(n29717), 
            .n29716(n29716), .n29715(n29715), .n29714(n29714), .n29713(n29713), 
            .n29712(n29712), .n29711(n29711), .n29710(n29710), .n29709(n29709), 
            .n29708(n29708), .n29707(n29707), .neopxl_color({neopxl_color}), 
            .n29706(n29706), .n29705(n29705), .\state_3__N_528[1] (state_3__N_528[1]), 
            .timer({timer}), .LED_c(LED_c), .n29323(n29323), .n29704(n29704), 
            .n29703(n29703), .n29702(n29702), .n29701(n29701), .n29700(n29700), 
            .n29699(n29699), .n29698(n29698), .n29697(n29697), .n29696(n29696), 
            .n29695(n29695), .n29694(n29694), .NEOPXL_c(NEOPXL_c), .n29633(n29633), 
            .n29623(n29623)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n39859), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n40308), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n40308), .I0(n3111), 
            .I1(VCC_net), .CO(n40309));
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n40307), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n39866), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22_adj_5144), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n947));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n40307), .I0(n3112), 
            .I1(VCC_net), .CO(n40308));
    SB_LUT4 encoder0_position_31__I_0_i1525_rep_22_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1525_rep_22_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22), 
            .I3(n39124), .O(pwm_setpoint_23__N_191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_5 (.CI(n39124), .I0(GND_net), .I1(n22), 
            .CO(n39125));
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n40306), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23), 
            .I3(n39123), .O(pwm_setpoint_23__N_191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16560_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n25135), .I3(GND_net), .O(n30087));   // verilog/coms.v(127[12] 300[6])
    defparam i16560_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n40306), .I0(n3113), 
            .I1(VCC_net), .CO(n40307));
    SB_LUT4 i16561_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n25135), .I3(GND_net), .O(n30088));   // verilog/coms.v(127[12] 300[6])
    defparam i16561_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16562_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n25135), .I3(GND_net), .O(n30089));   // verilog/coms.v(127[12] 300[6])
    defparam i16562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16563_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n25135), .I3(GND_net), .O(n30090));   // verilog/coms.v(127[12] 300[6])
    defparam i16563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16564_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n25135), .I3(GND_net), .O(n30091));   // verilog/coms.v(127[12] 300[6])
    defparam i16564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16565_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n25135), .I3(GND_net), .O(n30092));   // verilog/coms.v(127[12] 300[6])
    defparam i16565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16566_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n25135), .I3(GND_net), .O(n30093));   // verilog/coms.v(127[12] 300[6])
    defparam i16566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16567_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n25135), .I3(GND_net), .O(n30094));   // verilog/coms.v(127[12] 300[6])
    defparam i16567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16568_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n25135), .I3(GND_net), .O(n30095));   // verilog/coms.v(127[12] 300[6])
    defparam i16568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16569_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n25135), .I3(GND_net), .O(n30096));   // verilog/coms.v(127[12] 300[6])
    defparam i16569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16570_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n25135), .I3(GND_net), .O(n30097));   // verilog/coms.v(127[12] 300[6])
    defparam i16570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16571_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n25135), .I3(GND_net), .O(n30098));   // verilog/coms.v(127[12] 300[6])
    defparam i16571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16572_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n25135), .I3(GND_net), .O(n30099));   // verilog/coms.v(127[12] 300[6])
    defparam i16572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16573_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n25135), .I3(GND_net), .O(n30100));   // verilog/coms.v(127[12] 300[6])
    defparam i16573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16574_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n25135), .I3(GND_net), .O(n30101));   // verilog/coms.v(127[12] 300[6])
    defparam i16574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16575_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n25135), .I3(GND_net), .O(n30102));   // verilog/coms.v(127[12] 300[6])
    defparam i16575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16576_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n25135), .I3(GND_net), .O(n30103));   // verilog/coms.v(127[12] 300[6])
    defparam i16576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16577_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n25135), .I3(GND_net), .O(n30104));   // verilog/coms.v(127[12] 300[6])
    defparam i16577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16578_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n25135), .I3(GND_net), .O(n30105));   // verilog/coms.v(127[12] 300[6])
    defparam i16578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16579_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n25135), .I3(GND_net), .O(n30106));   // verilog/coms.v(127[12] 300[6])
    defparam i16579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16580_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n25135), .I3(GND_net), .O(n30107));   // verilog/coms.v(127[12] 300[6])
    defparam i16580_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16581_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n25135), .I3(GND_net), .O(n30108));   // verilog/coms.v(127[12] 300[6])
    defparam i16581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16582_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n25135), .I3(GND_net), .O(n30109));   // verilog/coms.v(127[12] 300[6])
    defparam i16582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16583_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n25135), .I3(GND_net), .O(n30110));   // verilog/coms.v(127[12] 300[6])
    defparam i16583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16584_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n25135), .I3(GND_net), .O(n30111));   // verilog/coms.v(127[12] 300[6])
    defparam i16584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16585_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n25135), .I3(GND_net), .O(n30112));   // verilog/coms.v(127[12] 300[6])
    defparam i16585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16586_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n25135), .I3(GND_net), .O(n30113));   // verilog/coms.v(127[12] 300[6])
    defparam i16586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16587_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n25135), .I3(GND_net), .O(n30114));   // verilog/coms.v(127[12] 300[6])
    defparam i16587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16588_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n25135), .I3(GND_net), .O(n30115));   // verilog/coms.v(127[12] 300[6])
    defparam i16588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16589_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n25135), 
            .I3(GND_net), .O(n30116));   // verilog/coms.v(127[12] 300[6])
    defparam i16589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16590_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n25135), 
            .I3(GND_net), .O(n30117));   // verilog/coms.v(127[12] 300[6])
    defparam i16590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16591_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n25135), 
            .I3(GND_net), .O(n30118));   // verilog/coms.v(127[12] 300[6])
    defparam i16591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16592_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n25135), 
            .I3(GND_net), .O(n30119));   // verilog/coms.v(127[12] 300[6])
    defparam i16592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16593_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n25135), 
            .I3(GND_net), .O(n30120));   // verilog/coms.v(127[12] 300[6])
    defparam i16593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16594_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n25135), 
            .I3(GND_net), .O(n30121));   // verilog/coms.v(127[12] 300[6])
    defparam i16594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16595_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n25135), 
            .I3(GND_net), .O(n30122));   // verilog/coms.v(127[12] 300[6])
    defparam i16595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16596_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n25135), 
            .I3(GND_net), .O(n30123));   // verilog/coms.v(127[12] 300[6])
    defparam i16596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16597_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n29176), 
            .I3(GND_net), .O(n30124));   // verilog/coms.v(127[12] 300[6])
    defparam i16597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16598_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n29176), 
            .I3(GND_net), .O(n30125));   // verilog/coms.v(127[12] 300[6])
    defparam i16598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16599_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n29176), 
            .I3(GND_net), .O(n30126));   // verilog/coms.v(127[12] 300[6])
    defparam i16599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16600_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n29176), 
            .I3(GND_net), .O(n30127));   // verilog/coms.v(127[12] 300[6])
    defparam i16600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16601_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n29176), 
            .I3(GND_net), .O(n30128));   // verilog/coms.v(127[12] 300[6])
    defparam i16601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16602_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n29176), 
            .I3(GND_net), .O(n30129));   // verilog/coms.v(127[12] 300[6])
    defparam i16602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16603_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n29176), 
            .I3(GND_net), .O(n30130));   // verilog/coms.v(127[12] 300[6])
    defparam i16603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16604_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n29176), 
            .I3(GND_net), .O(n30131));   // verilog/coms.v(127[12] 300[6])
    defparam i16604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16605_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n29176), 
            .I3(GND_net), .O(n30132));   // verilog/coms.v(127[12] 300[6])
    defparam i16605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16606_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n29176), 
            .I3(GND_net), .O(n30133));   // verilog/coms.v(127[12] 300[6])
    defparam i16606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16607_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n29176), 
            .I3(GND_net), .O(n30134));   // verilog/coms.v(127[12] 300[6])
    defparam i16607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16608_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n29176), 
            .I3(GND_net), .O(n30135));   // verilog/coms.v(127[12] 300[6])
    defparam i16608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16609_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n29176), 
            .I3(GND_net), .O(n30136));   // verilog/coms.v(127[12] 300[6])
    defparam i16609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16610_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n29176), 
            .I3(GND_net), .O(n30137));   // verilog/coms.v(127[12] 300[6])
    defparam i16610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16611_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n29176), 
            .I3(GND_net), .O(n30138));   // verilog/coms.v(127[12] 300[6])
    defparam i16611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16612_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n29176), 
            .I3(GND_net), .O(n30139));   // verilog/coms.v(127[12] 300[6])
    defparam i16612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16613_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n29176), 
            .I3(GND_net), .O(n30140));   // verilog/coms.v(127[12] 300[6])
    defparam i16613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16614_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n29176), 
            .I3(GND_net), .O(n30141));   // verilog/coms.v(127[12] 300[6])
    defparam i16614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16616_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n29176), 
            .I3(GND_net), .O(n30143));   // verilog/coms.v(127[12] 300[6])
    defparam i16616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16617_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n29176), 
            .I3(GND_net), .O(n30144));   // verilog/coms.v(127[12] 300[6])
    defparam i16617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16618_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n29176), 
            .I3(GND_net), .O(n30145));   // verilog/coms.v(127[12] 300[6])
    defparam i16618_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n39859), .I0(n2227), 
            .I1(VCC_net), .CO(n39860));
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n6662), 
            .D(n1077), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16619_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n29176), 
            .I3(GND_net), .O(n30146));   // verilog/coms.v(127[12] 300[6])
    defparam i16619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16620_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n29176), 
            .I3(GND_net), .O(n30147));   // verilog/coms.v(127[12] 300[6])
    defparam i16620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16621_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n29176), 
            .I3(GND_net), .O(n30148));   // verilog/coms.v(127[12] 300[6])
    defparam i16621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16622_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n29176), 
            .I3(GND_net), .O(n30149));   // verilog/coms.v(127[12] 300[6])
    defparam i16622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16623_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n29176), 
            .I3(GND_net), .O(n30150));   // verilog/coms.v(127[12] 300[6])
    defparam i16623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16624_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n29176), 
            .I3(GND_net), .O(n30151));   // verilog/coms.v(127[12] 300[6])
    defparam i16624_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n6662), 
            .D(n1078), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n6662), 
            .D(n1079), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n6662), 
            .D(n1080), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16625_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n29176), 
            .I3(GND_net), .O(n30152));   // verilog/coms.v(127[12] 300[6])
    defparam i16625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16626_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n29176), 
            .I3(GND_net), .O(n30153));   // verilog/coms.v(127[12] 300[6])
    defparam i16626_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n6662), 
            .D(n1081), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16627_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n29176), 
            .I3(GND_net), .O(n30154));   // verilog/coms.v(127[12] 300[6])
    defparam i16627_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n6662), 
            .D(n1082), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n6662), 
            .D(n1083), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16628_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30155));   // verilog/coms.v(127[12] 300[6])
    defparam i16628_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n6662), 
            .D(n1084), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n6662), 
            .D(n1085), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n6662), 
            .D(n1086), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16629_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30156));   // verilog/coms.v(127[12] 300[6])
    defparam i16629_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n6662), 
            .D(n1087), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n6662), 
            .D(n1088), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n6662), 
            .D(n1089), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16630_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30157));   // verilog/coms.v(127[12] 300[6])
    defparam i16630_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n6662), 
            .D(n1090), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n6662), 
            .D(n1091), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n6662), 
            .D(n1092), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n6662), 
            .D(n1093), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n6662), 
            .D(n1094), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16631_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30158));   // verilog/coms.v(127[12] 300[6])
    defparam i16631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16632_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30159));   // verilog/coms.v(127[12] 300[6])
    defparam i16632_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n6662), 
            .D(n1095), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16633_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30160));   // verilog/coms.v(127[12] 300[6])
    defparam i16633_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n6662), 
            .D(n1096), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n6662), 
            .D(n1097), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n6662), 
            .D(n1098), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n6662), 
            .D(n1099), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i16634_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30161));   // verilog/coms.v(127[12] 300[6])
    defparam i16634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16635_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30162));   // verilog/coms.v(127[12] 300[6])
    defparam i16635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16636_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30163));   // verilog/coms.v(127[12] 300[6])
    defparam i16636_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n6662), 
            .D(n1100), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n6662), 
            .D(n1101), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n6662), 
            .D(n1102), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n6662), 
            .D(n1103), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n6662), 
            .D(n1104), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n6662), 
            .D(n1105), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n6662), 
            .D(n1106), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n6662), 
            .D(n1107), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i35453_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n47066), 
            .O(n1752));
    defparam i35453_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16637_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30164));   // verilog/coms.v(127[12] 300[6])
    defparam i16637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16638_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30165));   // verilog/coms.v(127[12] 300[6])
    defparam i16638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16639_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30166));   // verilog/coms.v(127[12] 300[6])
    defparam i16639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16640_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30167));   // verilog/coms.v(127[12] 300[6])
    defparam i16640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16641_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30168));   // verilog/coms.v(127[12] 300[6])
    defparam i16641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16642_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30169));   // verilog/coms.v(127[12] 300[6])
    defparam i16642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16643_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30170));   // verilog/coms.v(127[12] 300[6])
    defparam i16643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16644_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30171));   // verilog/coms.v(127[12] 300[6])
    defparam i16644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16645_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30172));   // verilog/coms.v(127[12] 300[6])
    defparam i16645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16646_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30173));   // verilog/coms.v(127[12] 300[6])
    defparam i16646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16647_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30174));   // verilog/coms.v(127[12] 300[6])
    defparam i16647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16648_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30175));   // verilog/coms.v(127[12] 300[6])
    defparam i16648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16649_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30176));   // verilog/coms.v(127[12] 300[6])
    defparam i16649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16650_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30177));   // verilog/coms.v(127[12] 300[6])
    defparam i16650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16651_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30178));   // verilog/coms.v(127[12] 300[6])
    defparam i16651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16652_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30179));   // verilog/coms.v(127[12] 300[6])
    defparam i16652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16653_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30180));   // verilog/coms.v(127[12] 300[6])
    defparam i16653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16654_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30181));   // verilog/coms.v(127[12] 300[6])
    defparam i16654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16655_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30182));   // verilog/coms.v(127[12] 300[6])
    defparam i16655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16656_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30183));   // verilog/coms.v(127[12] 300[6])
    defparam i16656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16657_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30184));   // verilog/coms.v(127[12] 300[6])
    defparam i16657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n39858), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16658_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n30185));   // verilog/coms.v(127[12] 300[6])
    defparam i16658_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n39858), .I0(n2228), 
            .I1(VCC_net), .CO(n39859));
    SB_LUT4 i16659_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n29176), .I3(GND_net), .O(n30186));   // verilog/coms.v(127[12] 300[6])
    defparam i16659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16157_3_lut (.I0(n29257), .I1(\ID_READOUT_FSM.state [0]), .I2(n6969), 
            .I3(GND_net), .O(n29684));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16157_3_lut.LUT_INIT = 16'h4646;
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n39857), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n39857), .I0(n2229), 
            .I1(GND_net), .CO(n39858));
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n39856), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n39856), .I0(n2230), 
            .I1(GND_net), .CO(n39857));
    SB_LUT4 i16661_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n29176), .I3(GND_net), .O(n30188));   // verilog/coms.v(127[12] 300[6])
    defparam i16661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16662_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n29176), .I3(GND_net), .O(n30189));   // verilog/coms.v(127[12] 300[6])
    defparam i16662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16663_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n29176), .I3(GND_net), .O(n30190));   // verilog/coms.v(127[12] 300[6])
    defparam i16663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n39855), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16664_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n29176), .I3(GND_net), .O(n30191));   // verilog/coms.v(127[12] 300[6])
    defparam i16664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16665_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n29176), .I3(GND_net), .O(n30192));   // verilog/coms.v(127[12] 300[6])
    defparam i16665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16666_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n29176), .I3(GND_net), .O(n30193));   // verilog/coms.v(127[12] 300[6])
    defparam i16666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16667_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n29176), .I3(GND_net), .O(n30194));   // verilog/coms.v(127[12] 300[6])
    defparam i16667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16668_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n29176), .I3(GND_net), .O(n30195));   // verilog/coms.v(127[12] 300[6])
    defparam i16668_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n39855), .I0(n2231), 
            .I1(VCC_net), .CO(n39856));
    SB_LUT4 i16669_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n29176), .I3(GND_net), .O(n30196));   // verilog/coms.v(127[12] 300[6])
    defparam i16669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16670_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n29176), .I3(GND_net), .O(n30197));   // verilog/coms.v(127[12] 300[6])
    defparam i16670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n39854), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n39854), .I0(n2232), 
            .I1(GND_net), .CO(n39855));
    SB_LUT4 i16671_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n29176), .I3(GND_net), .O(n30198));   // verilog/coms.v(127[12] 300[6])
    defparam i16671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16672_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n29176), .I3(GND_net), .O(n30199));   // verilog/coms.v(127[12] 300[6])
    defparam i16672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16673_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n29176), .I3(GND_net), .O(n30200));   // verilog/coms.v(127[12] 300[6])
    defparam i16673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16674_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n29176), .I3(GND_net), .O(n30201));   // verilog/coms.v(127[12] 300[6])
    defparam i16674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16675_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n29176), .I3(GND_net), .O(n30202));   // verilog/coms.v(127[12] 300[6])
    defparam i16675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16676_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n29176), .I3(GND_net), .O(n30203));   // verilog/coms.v(127[12] 300[6])
    defparam i16676_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16677_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n29176), .I3(GND_net), .O(n30204));   // verilog/coms.v(127[12] 300[6])
    defparam i16677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16678_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n29176), .I3(GND_net), .O(n30205));   // verilog/coms.v(127[12] 300[6])
    defparam i16678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n39853), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16679_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n29176), .I3(GND_net), .O(n30206));   // verilog/coms.v(127[12] 300[6])
    defparam i16679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16680_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n29176), .I3(GND_net), .O(n30207));   // verilog/coms.v(127[12] 300[6])
    defparam i16680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16681_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n29176), .I3(GND_net), .O(n30208));   // verilog/coms.v(127[12] 300[6])
    defparam i16681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16682_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n29176), .I3(GND_net), .O(n30209));   // verilog/coms.v(127[12] 300[6])
    defparam i16682_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_10_add_3_4 (.CI(n39123), .I0(GND_net), .I1(n23), 
            .CO(n39124));
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n39853), .I0(n2233), 
            .I1(VCC_net), .CO(n39854));
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n39853));
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n50987), .I1(n2115), 
            .I2(VCC_net), .I3(n39852), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n39851), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n39851), .I0(n2116), 
            .I1(VCC_net), .CO(n39852));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n39850), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16145_4_lut (.I0(n29246), .I1(r_Bit_Index[0]), .I2(n44059), 
            .I3(r_SM_Main[1]), .O(n29672));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16145_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 i16685_4_lut (.I0(state_7__N_4103[3]), .I1(data[6]), .I2(n35422), 
            .I3(n27984), .O(n30212));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16685_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i16140_4_lut (.I0(n29234), .I1(r_Bit_Index_adj_5300[0]), .I2(n44068), 
            .I3(r_SM_Main_adj_5298[1]), .O(n29667));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i16140_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 i1_4_lut (.I0(n6969), .I1(n21743), .I2(data_ready), .I3(\ID_READOUT_FSM.state [0]), 
            .O(n44859));
    defparam i1_4_lut.LUT_INIT = 16'heaee;
    SB_LUT4 i35425_1_lut (.I0(n1653_adj_5178), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n50863));
    defparam i35425_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(n35141), .I2(\ID_READOUT_FSM.state [1]), 
            .I3(n44859), .O(n29257));
    defparam i2_4_lut.LUT_INIT = 16'h4c00;
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n6969), .I2(n29257), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n43275));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(h3), .I1(commutation_state[1]), .I2(h2), 
            .I3(h1), .O(n43957));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'hd054;
    SB_LUT4 i35445_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50883));
    defparam i35445_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34872_3_lut (.I0(n1727), .I1(n1794), .I2(n1752), .I3(GND_net), 
            .O(n1826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34872_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16180_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n43061), .I3(GND_net), .O(n29707));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16180_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34870_3_lut (.I0(n1726), .I1(n1793), .I2(n1752), .I3(GND_net), 
            .O(n1825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34870_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16181_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n43061), .I3(GND_net), .O(n29708));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16181_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n39850), .I0(n2117), 
            .I1(VCC_net), .CO(n39851));
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n39867), .I0(n2219), 
            .I1(VCC_net), .CO(n39868));
    SB_LUT4 i16182_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n43061), .I3(GND_net), .O(n29709));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16183_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n43061), .I3(GND_net), .O(n29710));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16184_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n43061), .I3(GND_net), .O(n29711));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n39849), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16185_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n43061), .I3(GND_net), .O(n29712));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16186_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n43061), .I3(GND_net), .O(n29713));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16187_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n43061), .I3(GND_net), .O(n29714));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16188_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n43061), .I3(GND_net), .O(n29715));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16189_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n43061), .I3(GND_net), .O(n29716));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16190_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n43061), .I3(GND_net), .O(n29717));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16191_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n43061), .I3(GND_net), .O(n29718));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16192_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n43061), .I3(GND_net), .O(n29719));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16193_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n43061), .I3(GND_net), .O(n29720));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16194_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n43061), .I3(GND_net), .O(n29721));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n40305), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16195_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n43061), .I3(GND_net), .O(n29722));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35454_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50892));
    defparam i35454_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16196_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n43061), .I3(GND_net), .O(n29723));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16197_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n43061), .I3(GND_net), .O(n29724));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1660 (.I0(\FRAME_MATCHER.state_31__N_2660 [2]), .I1(n7_adj_5185), 
            .I2(\FRAME_MATCHER.i_31__N_2624 ), .I3(n3303), .O(n6_adj_5186));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1660.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1661 (.I0(\FRAME_MATCHER.state_31__N_2660 [2]), .I1(\FRAME_MATCHER.i_31__N_2622 ), 
            .I2(n45880), .I3(n14_adj_5229), .O(n7_adj_5179));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1661.LUT_INIT = 16'heece;
    SB_LUT4 i4_4_lut (.I0(n7_adj_5179), .I1(n82), .I2(n6_adj_5186), .I3(n4_adj_5093), 
            .O(n51594));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut.LUT_INIT = 16'hfbfa;
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n39849), .I0(n2118), 
            .I1(VCC_net), .CO(n39850));
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n39848), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n39848), .I0(n2119), 
            .I1(VCC_net), .CO(n39849));
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n39847), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n39847), .I0(n2120), 
            .I1(VCC_net), .CO(n39848));
    SB_LUT4 i1_4_lut_adj_1662 (.I0(n14_adj_5229), .I1(n45880), .I2(\FRAME_MATCHER.i_31__N_2626 ), 
            .I3(n4452), .O(n5_adj_5187));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'hbbfb;
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n39846), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n39846), .I0(n2121), 
            .I1(VCC_net), .CO(n39847));
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n39845), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n39845), .I0(n2122), 
            .I1(VCC_net), .CO(n39846));
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n40305), .I0(n3114), 
            .I1(VCC_net), .CO(n40306));
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n39867), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n39868), .I0(n2218), 
            .I1(VCC_net), .CO(n39869));
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n39844), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n39844), .I0(n2123), 
            .I1(VCC_net), .CO(n39845));
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n39843), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n40304), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n39843), .I0(n2124), 
            .I1(VCC_net), .CO(n39844));
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n39842), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n39842), .I0(n2125), 
            .I1(VCC_net), .CO(n39843));
    SB_LUT4 i1_4_lut_adj_1663 (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(n63), 
            .I2(n3303), .I3(n123), .O(n4_adj_5221));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1663.LUT_INIT = 16'haaa2;
    SB_LUT4 i1_3_lut (.I0(n123), .I1(n5_adj_5187), .I2(n63), .I3(GND_net), 
            .O(n7_adj_5220));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut.LUT_INIT = 16'h8c8c;
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.i_31__N_2622 ), .I1(n7_adj_5220), 
            .I2(n4_adj_5221), .I3(n1), .O(n51593));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16200_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n29176), .I3(GND_net), .O(n29727));   // verilog/coms.v(127[12] 300[6])
    defparam i16200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16201_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n29176), .I3(GND_net), .O(n29728));   // verilog/coms.v(127[12] 300[6])
    defparam i16201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16202_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n29176), .I3(GND_net), .O(n29729));   // verilog/coms.v(127[12] 300[6])
    defparam i16202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16203_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n29176), .I3(GND_net), .O(n29730));   // verilog/coms.v(127[12] 300[6])
    defparam i16203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16204_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n29176), .I3(GND_net), .O(n29731));   // verilog/coms.v(127[12] 300[6])
    defparam i16204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16205_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n29176), .I3(GND_net), .O(n29732));   // verilog/coms.v(127[12] 300[6])
    defparam i16205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16206_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n29176), .I3(GND_net), .O(n29733));   // verilog/coms.v(127[12] 300[6])
    defparam i16206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16207_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n29176), .I3(GND_net), .O(n29734));   // verilog/coms.v(127[12] 300[6])
    defparam i16207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16208_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n29176), .I3(GND_net), .O(n29735));   // verilog/coms.v(127[12] 300[6])
    defparam i16208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_5097));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16209_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n29176), .I3(GND_net), .O(n29736));   // verilog/coms.v(127[12] 300[6])
    defparam i16209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16210_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n29176), .I3(GND_net), .O(n29737));   // verilog/coms.v(127[12] 300[6])
    defparam i16210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16211_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n29176), .I3(GND_net), .O(n29738));   // verilog/coms.v(127[12] 300[6])
    defparam i16211_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n40304), .I0(n3115), 
            .I1(VCC_net), .CO(n40305));
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n39841), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n39841), .I0(n2126), 
            .I1(VCC_net), .CO(n39842));
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n39840), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n39840), .I0(n2127), 
            .I1(VCC_net), .CO(n39841));
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n39839), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n39839), .I0(n2128), 
            .I1(VCC_net), .CO(n39840));
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35029_3_lut (.I0(n1628), .I1(n1695), .I2(n1653_adj_5178), 
            .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i35029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34962_3_lut (.I0(n1826), .I1(n1893), .I2(n1851), .I3(GND_net), 
            .O(n1925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35497_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50935));
    defparam i35497_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n39838), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20_adj_5146), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n945));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19_adj_5147), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n944));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18_adj_5148), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n943));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n40303), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16212_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n29176), .I3(GND_net), .O(n29739));   // verilog/coms.v(127[12] 300[6])
    defparam i16212_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n39838), .I0(n2129), 
            .I1(GND_net), .CO(n39839));
    SB_LUT4 i16213_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n29176), .I3(GND_net), .O(n29740));   // verilog/coms.v(127[12] 300[6])
    defparam i16213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n39837), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut (.I0(dti_counter[7]), .I1(dti_counter[4]), .I2(dti_counter[5]), 
            .I3(dti_counter[6]), .O(n14_adj_5106));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n39837), .I0(n2130), 
            .I1(GND_net), .CO(n39838));
    SB_LUT4 i16214_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n29176), .I3(GND_net), .O(n29741));   // verilog/coms.v(127[12] 300[6])
    defparam i16214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n39836), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16215_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n29176), .I3(GND_net), .O(n29742));   // verilog/coms.v(127[12] 300[6])
    defparam i16215_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n40303), .I0(n3116), 
            .I1(VCC_net), .CO(n40304));
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n39868), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n39836), .I0(n2131), 
            .I1(VCC_net), .CO(n39837));
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16216_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n29176), .I3(GND_net), .O(n29743));   // verilog/coms.v(127[12] 300[6])
    defparam i16216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13_adj_5155), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n938));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34874_3_lut (.I0(n1926), .I1(n1993), .I2(n1950), .I3(GND_net), 
            .O(n2025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34874_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1664 (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n46975));
    defparam i3_4_lut_adj_1664.LUT_INIT = 16'h0004;
    SB_LUT4 i16217_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n29176), .I3(GND_net), .O(n29744));   // verilog/coms.v(127[12] 300[6])
    defparam i16217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35575_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51013));
    defparam i35575_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(244[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16218_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n29176), .I3(GND_net), .O(n29745));   // verilog/coms.v(127[12] 300[6])
    defparam i16218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16219_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n29176), .I3(GND_net), .O(n29746));   // verilog/coms.v(127[12] 300[6])
    defparam i16219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35523_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50961));
    defparam i35523_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n39869), .I0(n2217), 
            .I1(VCC_net), .CO(n39870));
    SB_LUT4 unary_minus_10_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5096));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_10_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_5095));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n39835), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n40302), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1248_rep_42_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1248_rep_42_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n39835), .I0(n2132), 
            .I1(GND_net), .CO(n39836));
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n39834), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n39834), .I0(n2133), 
            .I1(VCC_net), .CO(n39835));
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n39834));
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n50961), .I1(n2016), 
            .I2(VCC_net), .I3(n39833), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n39869), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n40302), .I0(n3117), 
            .I1(VCC_net), .CO(n40303));
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n40301), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n39870), .I0(n2216), 
            .I1(VCC_net), .CO(n39871));
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n40301), .I0(n3118), 
            .I1(VCC_net), .CO(n40302));
    SB_LUT4 encoder0_position_31__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n39870), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34879_3_lut (.I0(n2126), .I1(n2193), .I2(n2148), .I3(GND_net), 
            .O(n2225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34879_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n39832), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n39832), .I0(n2017), 
            .I1(VCC_net), .CO(n39833));
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n39831), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n39831), .I0(n2018), 
            .I1(VCC_net), .CO(n39832));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n39830), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n39871), .I0(n2215), 
            .I1(VCC_net), .CO(n39872));
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n39830), .I0(n2019), 
            .I1(VCC_net), .CO(n39831));
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n39829), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n39829), .I0(n2020), 
            .I1(VCC_net), .CO(n39830));
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n39828), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n39828), .I0(n2021), 
            .I1(VCC_net), .CO(n39829));
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n39827), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n39871), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n39827), .I0(n2022), 
            .I1(VCC_net), .CO(n39828));
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n39826), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n39826), .I0(n2023), 
            .I1(VCC_net), .CO(n39827));
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n40300), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n39825), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n39825), .I0(n2024), 
            .I1(VCC_net), .CO(n39826));
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(n51013), .I1(n2214), 
            .I2(VCC_net), .I3(n39872), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i34880_3_lut (.I0(n2225), .I1(n2292), .I2(n2247), .I3(GND_net), 
            .O(n2324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34880_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n39824), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n39824), .I0(n2025), 
            .I1(VCC_net), .CO(n39825));
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n39823), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n40300), .I0(n3119), 
            .I1(VCC_net), .CO(n40301));
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n39823), .I0(n2026), 
            .I1(VCC_net), .CO(n39824));
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut (.I0(dti_counter[0]), .I1(n14_adj_5106), .I2(n10_adj_5107), 
            .I3(dti_counter[3]), .O(n25336));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n40299), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n39822), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n39822), .I0(n2027), 
            .I1(VCC_net), .CO(n39823));
    SB_LUT4 encoder0_position_31__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1665 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5231));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_4_lut_adj_1665.LUT_INIT = 16'h7bde;
    SB_LUT4 encoder0_position_31__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n39821), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n39821), .I0(n2028), 
            .I1(VCC_net), .CO(n39822));
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n39820), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n39820), .I0(n2029), 
            .I1(GND_net), .CO(n39821));
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n39819), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n39819), .I0(n2030), 
            .I1(GND_net), .CO(n39820));
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n39818), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n39818), .I0(n2031), 
            .I1(VCC_net), .CO(n39819));
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n39817), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n39817), .I0(n2032), 
            .I1(GND_net), .CO(n39818));
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n39816), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n39816), .I0(n2033), 
            .I1(VCC_net), .CO(n39817));
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n39816));
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n50935), .I1(n1917), 
            .I2(VCC_net), .I3(n39815), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n39814), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n39814), .I0(n1918), 
            .I1(VCC_net), .CO(n39815));
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n39813), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n39813), .I0(n1919), 
            .I1(VCC_net), .CO(n39814));
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n39812), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n39812), .I0(n1920), 
            .I1(VCC_net), .CO(n39813));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n39811), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n39811), .I0(n1921), 
            .I1(VCC_net), .CO(n39812));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n39810), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n39810), .I0(n1922), 
            .I1(VCC_net), .CO(n39811));
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n39809), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n39809), .I0(n1923), 
            .I1(VCC_net), .CO(n39810));
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n39808), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n39808), .I0(n1924), 
            .I1(VCC_net), .CO(n39809));
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n39807), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n39807), .I0(n1925), 
            .I1(VCC_net), .CO(n39808));
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n39806), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n40299), .I0(n3120), 
            .I1(VCC_net), .CO(n40300));
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n39806), .I0(n1926), 
            .I1(VCC_net), .CO(n39807));
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n39805), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n40298), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n39805), .I0(n1927), 
            .I1(VCC_net), .CO(n39806));
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n39804), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n40298), .I0(n3121), 
            .I1(VCC_net), .CO(n40299));
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n39804), .I0(n1928), 
            .I1(VCC_net), .CO(n39805));
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n40297), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n39803), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n39803), .I0(n1929), 
            .I1(GND_net), .CO(n39804));
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n39802), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n39802), .I0(n1930), 
            .I1(GND_net), .CO(n39803));
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n40297), .I0(n3122), 
            .I1(VCC_net), .CO(n40298));
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n39801), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n40296), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n39801), .I0(n1931), 
            .I1(VCC_net), .CO(n39802));
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n39800), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n40296), .I0(n3123), 
            .I1(VCC_net), .CO(n40297));
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n40295), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n40295), .I0(n3124), 
            .I1(VCC_net), .CO(n40296));
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n39800), .I0(n1932), 
            .I1(GND_net), .CO(n39801));
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n39799), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n39799), .I0(n1933), 
            .I1(VCC_net), .CO(n39800));
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n39799));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23_adj_5143), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n948));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n50892), .I1(n1818), 
            .I2(VCC_net), .I3(n39798), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25_adj_5141), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n950));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n39797), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n39797), .I0(n1819), 
            .I1(VCC_net), .CO(n39798));
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n39796), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n39796), .I0(n1820), 
            .I1(VCC_net), .CO(n39797));
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n39795), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n40294), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n39795), .I0(n1821), 
            .I1(VCC_net), .CO(n39796));
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n40294), .I0(n3125), 
            .I1(VCC_net), .CO(n40295));
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n40293), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n40293), .I0(n3126), 
            .I1(VCC_net), .CO(n40294));
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n39794), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n39794), .I0(n1822), 
            .I1(VCC_net), .CO(n39795));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_5156), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n937));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n39793), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n39793), .I0(n1823), 
            .I1(VCC_net), .CO(n39794));
    SB_LUT4 encoder0_position_31__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n39792), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n40292), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n39792), .I0(n1824), 
            .I1(VCC_net), .CO(n39793));
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n6662), 
            .D(n1108), .R(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35601_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51039));
    defparam i35601_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n40292), .I0(n3127), 
            .I1(VCC_net), .CO(n40293));
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n39791), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n39791), .I0(n1825), 
            .I1(VCC_net), .CO(n39792));
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n39790), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n39790), .I0(n1826), 
            .I1(VCC_net), .CO(n39791));
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n39789), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n39789), .I0(n1827), 
            .I1(VCC_net), .CO(n39790));
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n39788), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n39788), .I0(n1828), 
            .I1(VCC_net), .CO(n39789));
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n39787), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n39787), .I0(n1829), 
            .I1(GND_net), .CO(n39788));
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n39786), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n39786), .I0(n1830), 
            .I1(GND_net), .CO(n39787));
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n39785), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1180_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1180_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n39785), .I0(n1831), 
            .I1(VCC_net), .CO(n39786));
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n39784), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n39784), .I0(n1832), 
            .I1(GND_net), .CO(n39785));
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n39783), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n39783), .I0(n1833), 
            .I1(VCC_net), .CO(n39784));
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n39783));
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n40291), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n50883), .I1(n1719), 
            .I2(VCC_net), .I3(n39782), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n39781), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n39781), .I0(n1720), 
            .I1(VCC_net), .CO(n39782));
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n39780), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16220_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n29176), .I3(GND_net), .O(n29747));   // verilog/coms.v(127[12] 300[6])
    defparam i16220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34876_3_lut (.I0(n1927), .I1(n1994), .I2(n1950), .I3(GND_net), 
            .O(n2026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34876_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16221_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n29176), .I3(GND_net), .O(n29748));   // verilog/coms.v(127[12] 300[6])
    defparam i16221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16222_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n29176), .I3(GND_net), .O(n29749));   // verilog/coms.v(127[12] 300[6])
    defparam i16222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16223_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n29176), .I3(GND_net), .O(n29750));   // verilog/coms.v(127[12] 300[6])
    defparam i16223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16224_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n29176), .I3(GND_net), .O(n29751));   // verilog/coms.v(127[12] 300[6])
    defparam i16224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1380_3_lut (.I0(n48680), .I1(n1827), 
            .I2(n50164), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n39780), .I0(n1721), 
            .I1(VCC_net), .CO(n39781));
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n39779), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35633_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51071));
    defparam i35633_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16225_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n29176), .I3(GND_net), .O(n29752));   // verilog/coms.v(127[12] 300[6])
    defparam i16225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16226_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n29176), .I3(GND_net), .O(n29753));   // verilog/coms.v(127[12] 300[6])
    defparam i16226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35549_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50987));
    defparam i35549_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n39779), .I0(n1722), 
            .I1(VCC_net), .CO(n39780));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n39778), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16227_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n29176), .I3(GND_net), .O(n29754));   // verilog/coms.v(127[12] 300[6])
    defparam i16227_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n40291), .I0(n3128), 
            .I1(VCC_net), .CO(n40292));
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n39778), .I0(n1723), 
            .I1(VCC_net), .CO(n39779));
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n39777), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n39777), .I0(n1724), 
            .I1(VCC_net), .CO(n39778));
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n39776), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n39776), .I0(n1725), 
            .I1(VCC_net), .CO(n39777));
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n39775), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n39775), .I0(n1726), 
            .I1(VCC_net), .CO(n39776));
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n39774), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n39774), .I0(n1727), 
            .I1(VCC_net), .CO(n39775));
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n39773), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n39773), .I0(n1728), 
            .I1(VCC_net), .CO(n39774));
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n39772), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n39772), .I0(n1729), 
            .I1(GND_net), .CO(n39773));
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n39771), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n39771), .I0(n1730), 
            .I1(GND_net), .CO(n39772));
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n40290), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n39770), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n39770), .I0(n1731), 
            .I1(VCC_net), .CO(n39771));
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n39769), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n39769), .I0(n1732), 
            .I1(GND_net), .CO(n39770));
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n39768), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_279));   // verilog/TinyFPGA_B.v(321[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i34877_3_lut (.I0(n2125), .I1(n2192), .I2(n2148), .I3(GND_net), 
            .O(n2224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34877_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34878_3_lut (.I0(n2224), .I1(n2291), .I2(n2247), .I3(GND_net), 
            .O(n2323));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34878_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n40290), .I0(n3129), 
            .I1(GND_net), .CO(n40291));
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n39768), .I0(n1733), 
            .I1(VCC_net), .CO(n39769));
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n39768));
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n50863), .I1(n1620), 
            .I2(VCC_net), .I3(n39767), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n39766), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n39766), .I0(n1621), 
            .I1(VCC_net), .CO(n39767));
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n39765), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n39765), .I0(n1622), 
            .I1(VCC_net), .CO(n39766));
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n40289), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n39764), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n40289), .I0(n3130), 
            .I1(GND_net), .CO(n40290));
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n39764), .I0(n1623), 
            .I1(VCC_net), .CO(n39765));
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n39763), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n39763), .I0(n1624), 
            .I1(VCC_net), .CO(n39764));
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n40288), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n39762), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n39762), .I0(n1625), 
            .I1(VCC_net), .CO(n39763));
    SB_LUT4 unary_minus_10_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24), 
            .I3(n39122), .O(pwm_setpoint_23__N_191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n39761), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n40288), .I0(n3131), 
            .I1(VCC_net), .CO(n40289));
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n40287), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n40287), .I0(n3132), 
            .I1(GND_net), .CO(n40288));
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n39761), .I0(n1626), 
            .I1(VCC_net), .CO(n39762));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n39760), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n39760), .I0(n1627), 
            .I1(VCC_net), .CO(n39761));
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n39759), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n39759), .I0(n1628), 
            .I1(VCC_net), .CO(n39760));
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n39758), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n39758), .I0(n1629), 
            .I1(GND_net), .CO(n39759));
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n39757), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n39757), .I0(n1630), 
            .I1(GND_net), .CO(n39758));
    SB_LUT4 i35715_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51153));
    defparam i35715_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1773_3_lut (.I0(n2610), .I1(n2677), 
            .I2(n2643), .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n39756), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n39756), .I0(n1631), 
            .I1(VCC_net), .CO(n39757));
    SB_CARRY unary_minus_10_add_3_3 (.CI(n39122), .I0(GND_net), .I1(n24), 
            .CO(n39123));
    SB_LUT4 encoder0_position_31__I_0_i1582_rep_21_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1582_rep_21_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n39755), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n39755), .I0(n1632), 
            .I1(GND_net), .CO(n39756));
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n40286), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n25), 
            .I3(VCC_net), .O(pwm_setpoint_23__N_191[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n40286), .I0(n3133), 
            .I1(VCC_net), .CO(n40287));
    SB_CARRY unary_minus_10_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25), 
            .CO(n39122));
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n39754), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n39078), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n39754), .I0(n1633), 
            .I1(VCC_net), .CO(n39755));
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n39754));
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n50840), .I1(n1521), 
            .I2(VCC_net), .I3(n39753), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n39752), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n39752), .I0(n1522), 
            .I1(VCC_net), .CO(n39753));
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n39751), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n39751), .I0(n1523), 
            .I1(VCC_net), .CO(n39752));
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n39750), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n39750), .I0(n1524), 
            .I1(VCC_net), .CO(n39751));
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n39749), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n39749), .I0(n1525), 
            .I1(VCC_net), .CO(n39750));
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n39748), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n39748), .I0(n1526), 
            .I1(VCC_net), .CO(n39749));
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n39747), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n39747), .I0(n1527), 
            .I1(VCC_net), .CO(n39748));
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n39746), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n39746), .I0(n1528), 
            .I1(VCC_net), .CO(n39747));
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n39745), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n39745), .I0(n1529), 
            .I1(GND_net), .CO(n39746));
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n39744), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_8 (.CI(n39104), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n39105));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_5153), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n940));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n39744), .I0(n1530), 
            .I1(GND_net), .CO(n39745));
    SB_LUT4 add_224_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n39121), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n39743), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n39743), .I0(n1531), 
            .I1(VCC_net), .CO(n39744));
    SB_LUT4 add_224_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n39120), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n39742), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n39742), .I0(n1532), 
            .I1(GND_net), .CO(n39743));
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n39741), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n39741), .I0(n1533), 
            .I1(VCC_net), .CO(n39742));
    SB_CARRY add_224_24 (.CI(n39120), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n39121));
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n39741));
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(n50822), .I1(n1422), 
            .I2(VCC_net), .I3(n39740), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n39739), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n39739), .I0(n1423), 
            .I1(VCC_net), .CO(n39740));
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n40286));
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n39738), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n39738), .I0(n1424), 
            .I1(VCC_net), .CO(n39739));
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n39737), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n39737), .I0(n1425), 
            .I1(VCC_net), .CO(n39738));
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n39736), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n39736), .I0(n1426), 
            .I1(VCC_net), .CO(n39737));
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n39735), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n39735), .I0(n1427), 
            .I1(VCC_net), .CO(n39736));
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n39734), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n39734), .I0(n1428), 
            .I1(VCC_net), .CO(n39735));
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n39733), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(GND_net), .I1(n3006), 
            .I2(VCC_net), .I3(n40285), .O(n3073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n39733), .I0(n1429), 
            .I1(GND_net), .CO(n39734));
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n39732), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n39732), .I0(n1430), 
            .I1(GND_net), .CO(n39733));
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n39731), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n39731), .I0(n1431), 
            .I1(VCC_net), .CO(n39732));
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n39730), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n39730), .I0(n1432), 
            .I1(GND_net), .CO(n39731));
    SB_LUT4 add_224_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n39119), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n40284), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_23 (.CI(n39119), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n39120));
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n39729), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n40284), .I0(n3007), 
            .I1(VCC_net), .CO(n40285));
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n39729), .I0(n1433), 
            .I1(VCC_net), .CO(n39730));
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n40283), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n40283), .I0(n3008), 
            .I1(VCC_net), .CO(n40284));
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n40282), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n39070), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n39729));
    SB_CARRY add_145_13 (.CI(n39078), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n39079));
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n40282), .I0(n3009), 
            .I1(VCC_net), .CO(n40283));
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n40281), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35852_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51290));
    defparam i35852_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n40281), .I0(n3010), 
            .I1(VCC_net), .CO(n40282));
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n40280), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n40280), .I0(n3011), 
            .I1(VCC_net), .CO(n40281));
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n40279), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n40279), .I0(n3012), 
            .I1(VCC_net), .CO(n40280));
    SB_LUT4 add_224_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n39118), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n40278), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n40278), .I0(n3013), 
            .I1(VCC_net), .CO(n40279));
    SB_CARRY add_224_22 (.CI(n39118), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n39119));
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n40277), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n40277), .I0(n3014), 
            .I1(VCC_net), .CO(n40278));
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n40276), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n39103), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n40276), .I0(n3015), 
            .I1(VCC_net), .CO(n40277));
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n40275), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n39077), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n40275), .I0(n3016), 
            .I1(VCC_net), .CO(n40276));
    SB_LUT4 add_224_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n39117), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n40274), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_21 (.CI(n39117), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n39118));
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n40274), .I0(n3017), 
            .I1(VCC_net), .CO(n40275));
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n40273), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_7 (.CI(n39103), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n39104));
    SB_LUT4 add_224_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n39116), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n50805), .I1(n1323), 
            .I2(VCC_net), .I3(n39718), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n40273), .I0(n3018), 
            .I1(VCC_net), .CO(n40274));
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n39717), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n39717), .I0(n1324), 
            .I1(VCC_net), .CO(n39718));
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n40272), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n40272), .I0(n3019), 
            .I1(VCC_net), .CO(n40273));
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n39716), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n40271), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n39716), .I0(n1325), 
            .I1(VCC_net), .CO(n39717));
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n40271), .I0(n3020), 
            .I1(VCC_net), .CO(n40272));
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n39715), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n40270), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n39715), .I0(n1326), 
            .I1(VCC_net), .CO(n39716));
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n40270), .I0(n3021), 
            .I1(VCC_net), .CO(n40271));
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n40269), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n39714), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n39714), .I0(n1327), 
            .I1(VCC_net), .CO(n39715));
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n40269), .I0(n3022), 
            .I1(VCC_net), .CO(n40270));
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n39713), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n40268), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n39713), .I0(n1328), 
            .I1(VCC_net), .CO(n39714));
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n40268), .I0(n3023), 
            .I1(VCC_net), .CO(n40269));
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n39712), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35307_2_lut (.I0(n25336), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_416));
    defparam i35307_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 unary_minus_10_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n39712), .I0(n1329), 
            .I1(GND_net), .CO(n39713));
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n39711), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n39711), .I0(n1330), 
            .I1(GND_net), .CO(n39712));
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n39710), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16148_4_lut (.I0(state_7__N_4103[3]), .I1(data[7]), .I2(n35422), 
            .I3(n28004), .O(n29675));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16148_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 unary_minus_10_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n39710), .I0(n1331), 
            .I1(VCC_net), .CO(n39711));
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n39709), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n39709), .I0(n1332), 
            .I1(GND_net), .CO(n39710));
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n39708), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n39708), .I0(n1333), 
            .I1(VCC_net), .CO(n39709));
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n40267), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n39708));
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n50789), .I1(n1224), 
            .I2(VCC_net), .I3(n39707), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n39706), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n39706), .I0(n1225), 
            .I1(VCC_net), .CO(n39707));
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n39705), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n39705), .I0(n1226), 
            .I1(VCC_net), .CO(n39706));
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n39704), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n39704), .I0(n1227), 
            .I1(VCC_net), .CO(n39705));
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n39703), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n39703), .I0(n1228), 
            .I1(VCC_net), .CO(n39704));
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n39702), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n39702), .I0(n1229), 
            .I1(GND_net), .CO(n39703));
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n39701), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n39701), .I0(n1230), 
            .I1(GND_net), .CO(n39702));
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n39700), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n39700), .I0(n1231), 
            .I1(VCC_net), .CO(n39701));
    SB_LUT4 add_224_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n39105), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n39699), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35848_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51286));
    defparam i35848_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n39699), .I0(n1232), 
            .I1(GND_net), .CO(n39700));
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n39698), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n39698), .I0(n1233), 
            .I1(VCC_net), .CO(n39699));
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n40267), .I0(n3024), 
            .I1(VCC_net), .CO(n40268));
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n39698));
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n50774), .I1(n1125), 
            .I2(VCC_net), .I3(n39697), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n39696), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n39696), .I0(n1126), 
            .I1(VCC_net), .CO(n39697));
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n39695), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHC_184 (.Q(GHC), .C(CLK_c), .E(n29125), .D(GHC_N_403), 
            .R(n29460));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY add_224_20 (.CI(n39116), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n39117));
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n39695), .I0(n1127), 
            .I1(VCC_net), .CO(n39696));
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n40266), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n39694), .O(n1195_adj_5177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n39694), .I0(n1128), 
            .I1(VCC_net), .CO(n39695));
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n39693), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5109));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n39693), .I0(n1129), 
            .I1(GND_net), .CO(n39694));
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n39692), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5110));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5111));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5112));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5113));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n39692), .I0(n1130), 
            .I1(GND_net), .CO(n39693));
    SB_LUT4 add_224_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n39102), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n39691), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n40266), .I0(n3025), 
            .I1(VCC_net), .CO(n40267));
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n39691), .I0(n1131), 
            .I1(VCC_net), .CO(n39692));
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n39690), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1666 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i6_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n39690), .I0(n1132), 
            .I1(GND_net), .CO(n39691));
    SB_LUT4 i7_4_lut_adj_1667 (.I0(ID[3]), .I1(n14), .I2(n10), .I3(ID[6]), 
            .O(n27826));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i7_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5100));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1668 (.I0(delay_counter[28]), .I1(n12_adj_5100), 
            .I2(delay_counter[25]), .I3(delay_counter[30]), .O(n27858));
    defparam i6_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_DFFESR GHB_182 (.Q(GHB), .C(CLK_c), .E(n29125), .D(GHB_N_389), 
            .R(n29460));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i2_3_lut (.I0(delay_counter[17]), .I1(delay_counter[16]), .I2(delay_counter[15]), 
            .I3(GND_net), .O(n27855));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_DFFESR GHA_180 (.Q(GHA), .C(CLK_c), .E(n29125), .D(GHA_N_367), 
            .R(n29460));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 mux_238_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5114));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5115));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut (.I0(delay_counter[3]), .I1(delay_counter[5]), .I2(delay_counter[4]), 
            .I3(GND_net), .O(n14_adj_5103));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n39689), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6_4_lut_adj_1669 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_5102));
    defparam i6_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5116));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut (.I0(n15_adj_5102), .I1(delay_counter[2]), .I2(n14_adj_5103), 
            .I3(delay_counter[6]), .O(n27861));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5117));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n39689), .I0(n1133), 
            .I1(VCC_net), .CO(n39690));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n40265), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35886_1_lut (.I0(n36493), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51324));
    defparam i35886_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n40265), .I0(n3026), 
            .I1(VCC_net), .CO(n40266));
    SB_LUT4 encoder0_position_31__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2195_3_lut (.I0(n3224), .I1(n3291), 
            .I2(n3237), .I3(GND_net), .O(n23_adj_5225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n40264), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4275_4_lut (.I0(n27861), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5182));
    defparam i4275_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1670 (.I0(n24_adj_5182), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n45643));
    defparam i2_4_lut_adj_1670.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1671 (.I0(n45643), .I1(delay_counter[18]), .I2(n27855), 
            .I3(GND_net), .O(n46788));
    defparam i2_3_lut_adj_1671.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n40264), .I0(n3027), 
            .I1(VCC_net), .CO(n40265));
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n39689));
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n40263), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n40263), .I0(n3028), 
            .I1(VCC_net), .CO(n40264));
    SB_LUT4 i2_4_lut_adj_1672 (.I0(delay_counter[23]), .I1(n46788), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5184));
    defparam i2_4_lut_adj_1672.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_1673 (.I0(n7_adj_5184), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n27858), .O(n62));
    defparam i4_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 i7032_3_lut (.I0(n62), .I1(\ID_READOUT_FSM.state [0]), .I2(delay_counter[31]), 
            .I3(GND_net), .O(n21743));
    defparam i7032_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i1_2_lut (.I0(delay_counter[12]), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_5230));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1674 (.I0(delay_counter[9]), .I1(n4_adj_5230), 
            .I2(delay_counter[10]), .I3(n27861), .O(n46068));
    defparam i2_4_lut_adj_1674.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5118));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_4_lut_adj_1675 (.I0(n46068), .I1(n27855), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n46806));
    defparam i2_4_lut_adj_1675.LUT_INIT = 16'hffec;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5119));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5120));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2194_3_lut (.I0(n3223), .I1(n3290), 
            .I2(n3237), .I3(GND_net), .O(n25_adj_5226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n40262), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5121));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2192_3_lut (.I0(n3221), .I1(n3288), 
            .I2(n3237), .I3(GND_net), .O(n29_adj_5228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34881_3_lut (.I0(n2128), .I1(n2195), .I2(n2148), .I3(GND_net), 
            .O(n2227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34881_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n3220), .I1(n21_adj_5224), .I2(n3287), 
            .I3(n3237), .O(n47072));
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1677 (.I0(n3219), .I1(n23_adj_5225), .I2(n3286), 
            .I3(n3237), .O(n47074));
    defparam i1_4_lut_adj_1677.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1678 (.I0(n3229), .I1(n29_adj_5228), .I2(n3296), 
            .I3(n3237), .O(n47076));
    defparam i1_4_lut_adj_1678.LUT_INIT = 16'heefc;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5181));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_adj_1679 (.I0(n3227), .I1(n19_adj_5223), .I2(n3294), 
            .I3(n3237), .O(n47080));
    defparam i1_4_lut_adj_1679.LUT_INIT = 16'heefc;
    SB_LUT4 i2_4_lut_adj_1680 (.I0(delay_counter[22]), .I1(n46806), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5183));
    defparam i2_4_lut_adj_1680.LUT_INIT = 16'ha8a0;
    SB_LUT4 i21935_4_lut (.I0(n7_adj_5183), .I1(delay_counter[31]), .I2(n27858), 
            .I3(n8_adj_5181), .O(n1195));   // verilog/TinyFPGA_B.v(378[14:38])
    defparam i21935_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 encoder0_position_31__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n40262), .I0(n3029), 
            .I1(GND_net), .CO(n40263));
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n40261), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n40261), .I0(n3030), 
            .I1(GND_net), .CO(n40262));
    SB_LUT4 i1_4_lut_adj_1681 (.I0(n3228), .I1(n25_adj_5226), .I2(n3295), 
            .I3(n3237), .O(n47078));
    defparam i1_4_lut_adj_1681.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5122));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1682 (.I0(n3218), .I1(n27_adj_5227), .I2(n3285), 
            .I3(n3237), .O(n47082));
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5123));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2188_3_lut (.I0(n3217), .I1(n3284), 
            .I2(n3237), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16035_4_lut (.I0(n6662), .I1(n1195), .I2(n21743), .I3(n27827), 
            .O(n29533));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16035_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i34882_3_lut (.I0(n2227), .I1(n2294), .I2(n2247), .I3(GND_net), 
            .O(n2326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34882_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(n47080), .I1(n47076), .I2(n47074), 
            .I3(n47072), .O(n47090));
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i16228_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n29176), .I3(GND_net), .O(n29755));   // verilog/coms.v(127[12] 300[6])
    defparam i16228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5124));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22592_4_lut (.I0(n652), .I1(n957), .I2(n3301), .I3(n3237), 
            .O(n36109));
    defparam i22592_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i22775_4_lut (.I0(n36109), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n36297));
    defparam i22775_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n40260), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5125));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n47090), .I1(n37), .I2(n47082), .I3(n47078), 
            .O(n47094));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n49621), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5108));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 encoder0_position_31__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n3216), .I1(n47094), .I2(n3283), .I3(n3237), 
            .O(n47096));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5126));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5127));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5128));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_224_11 (.CI(n39107), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n39108));
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n40260), .I0(n3031), 
            .I1(VCC_net), .CO(n40261));
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n40259), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5129));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5130));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22873_4_lut (.I0(n36297), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n36395));
    defparam i22873_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_31__I_0_i2186_3_lut (.I0(n3215), .I1(n3282), 
            .I2(n3237), .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n41), .I1(n36395), .I2(n47096), .I3(n5_adj_5108), 
            .O(n47100));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n3214), .I1(n47100), .I2(n3281), .I3(n3237), 
            .O(n47102));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'heefc;
    SB_CARRY add_224_6 (.CI(n39102), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n39103));
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5131));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(n3213), .I1(n47102), .I2(n3280), .I3(n3237), 
            .O(n47104));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5104));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1689 (.I0(n3212), .I1(n47104), .I2(n3279), .I3(n3237), 
            .O(n47106));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n40259), .I0(n3032), 
            .I1(GND_net), .CO(n40260));
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n3211), .I1(n47106), .I2(n3278), .I3(n3237), 
            .O(n47108));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n3210), .I1(n47108), .I2(n3277), .I3(n3237), 
            .O(n47110));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n3209), .I1(n47110), .I2(n3276), .I3(n3237), 
            .O(n47112));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(n3208), .I1(n47112), .I2(n3275), .I3(n3237), 
            .O(n47114));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n3207), .I1(n47114), .I2(n3274), .I3(n3237), 
            .O(n47116));
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35889_4_lut (.I0(n61), .I1(n48576), .I2(n59), .I3(n47116), 
            .O(n36493));
    defparam i35889_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_5154), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n939));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n40258), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n40258), .I0(n3033), 
            .I1(VCC_net), .CO(n40259));
    SB_LUT4 mux_238_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_224_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n39115), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16152_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5152), 
            .I3(n27976), .O(n29679));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16152_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_adj_1695 (.I0(state_adj_5307[0]), .I1(n49702), .I2(n6387), 
            .I3(n35178), .O(n8_adj_5158));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_adj_1695.LUT_INIT = 16'h3afa;
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(CLK_c), 
            .E(n6_adj_5180), .D(commutation_state_7__N_216[0]), .S(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_5166), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i641_3_lut (.I0(n628), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100_adj_5175), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35045_3_lut (.I0(n1627), .I1(n1694), .I2(n1653_adj_5178), 
            .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i35045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34960_3_lut (.I0(n1825), .I1(n1892), .I2(n1851), .I3(GND_net), 
            .O(n1924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34960_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29517_3_lut (.I0(n4_adj_5091), .I1(n7352), .I2(n44865), .I3(GND_net), 
            .O(n44868));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29518_3_lut (.I0(encoder0_position[29]), .I1(n44868), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095_adj_5170), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22777_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n36299));
    defparam i22777_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1696 (.I0(n3225), .I1(n3221), .I2(n3224), .I3(n3219), 
            .O(n47706));
    defparam i1_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1697 (.I0(n3222), .I1(n3226), .I2(GND_net), .I3(GND_net), 
            .O(n47696));
    defparam i1_2_lut_adj_1697.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n3228), .I1(n3220), .I2(n3227), .I3(n3223), 
            .O(n47708));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n47708), .I1(n47696), .I2(n47706), 
            .I3(n3218), .O(n47712));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n3229), .I1(n36299), .I2(n3230), .I3(n3231), 
            .O(n45319));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n3215), .I1(n3216), .I2(n47712), .I3(n3217), 
            .O(n47718));
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n3213), .I1(n3214), .I2(n47718), .I3(n45319), 
            .O(n47724));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n47724), 
            .O(n47730));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n47730), 
            .O(n47736));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i35885_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n47736), 
            .O(n3237));
    defparam i35885_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n40258));
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n51219), .I1(n2907), 
            .I2(VCC_net), .I3(n40257), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1316_rep_36_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1316_rep_36_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1450_rep_23_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1450_rep_23_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1517_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n2224), .I1(n2226), .I2(n2227), .I3(n2225), 
            .O(n47542));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'hfffe;
    SB_LUT4 i22631_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n36149));
    defparam i22631_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n2222), .I1(n47542), .I2(n2223), .I3(n2228), 
            .O(n47546));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(n2229), .I1(n36149), .I2(n2230), .I3(n2231), 
            .O(n45257));
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n2220), .I1(n45257), .I2(n2221), .I3(n47546), 
            .O(n47552));
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n47552), 
            .O(n47558));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i35579_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n47558), 
            .O(n2247));
    defparam i35579_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n40256), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n40256), .I0(n2908), 
            .I1(VCC_net), .CO(n40257));
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n40255), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n40255), .I0(n2909), 
            .I1(VCC_net), .CO(n40256));
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n40254), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5099));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n40254), .I0(n2910), 
            .I1(VCC_net), .CO(n40255));
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n40253), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n40253), .I0(n2911), 
            .I1(VCC_net), .CO(n40254));
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n40252), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n40252), .I0(n2912), 
            .I1(VCC_net), .CO(n40253));
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n40251), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n40251), .I0(n2913), 
            .I1(VCC_net), .CO(n40252));
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n40250), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n40250), .I0(n2914), 
            .I1(VCC_net), .CO(n40251));
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n40249), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n40249), .I0(n2915), 
            .I1(VCC_net), .CO(n40250));
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n40248), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n40248), .I0(n2916), 
            .I1(VCC_net), .CO(n40249));
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n40247), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n40247), .I0(n2917), 
            .I1(VCC_net), .CO(n40248));
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n40246), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n40246), .I0(n2918), 
            .I1(VCC_net), .CO(n40247));
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2041_3_lut (.I0(n3006), .I1(n3073), 
            .I2(n3039), .I3(GND_net), .O(n3105));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(n3119), .I1(n3126), .I2(n3127), .I3(n3128), 
            .O(n47300));
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_10_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_224_19 (.CI(n39115), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n39116));
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n3120), .I1(n3124), .I2(n3123), .I3(n3125), 
            .O(n47298));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n47300), .I1(n3122), .I2(n3118), .I3(n3121), 
            .O(n47302));
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 i22779_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n36301));
    defparam i22779_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n3116), .I1(n47302), .I2(n3117), .I3(n47298), 
            .O(n47308));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n3129), .I1(n36301), .I2(n3130), .I3(n3131), 
            .O(n45275));
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(n3114), .I1(n3115), .I2(n45275), .I3(n47308), 
            .O(n47314));
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n40245), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n47314), 
            .O(n47320));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n40245), .I0(n2919), 
            .I1(VCC_net), .CO(n40246));
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n40244), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n40244), .I0(n2920), 
            .I1(VCC_net), .CO(n40245));
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n47320), 
            .O(n47326));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n40243), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n40243), .I0(n2921), 
            .I1(VCC_net), .CO(n40244));
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n40242), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35851_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n47326), 
            .O(n3138));
    defparam i35851_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n40242), .I0(n2922), 
            .I1(VCC_net), .CO(n40243));
    SB_LUT4 dti_counter_2056_add_4_9_lut (.I0(n49682), .I1(n35282), .I2(dti_counter[7]), 
            .I3(n40383), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 add_224_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n39101), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n40241), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 dti_counter_2056_add_4_8_lut (.I0(n49681), .I1(n35282), .I2(dti_counter[6]), 
            .I3(n40382), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2056_add_4_8 (.CI(n40382), .I0(n35282), .I1(dti_counter[6]), 
            .CO(n40383));
    SB_LUT4 dti_counter_2056_add_4_7_lut (.I0(n49680), .I1(n35282), .I2(dti_counter[5]), 
            .I3(n40381), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n40241), .I0(n2923), 
            .I1(VCC_net), .CO(n40242));
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n40240), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2056_add_4_7 (.CI(n40381), .I0(n35282), .I1(dti_counter[5]), 
            .CO(n40382));
    SB_LUT4 dti_counter_2056_add_4_6_lut (.I0(n49679), .I1(n35282), .I2(dti_counter[4]), 
            .I3(n40380), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_CARRY dti_counter_2056_add_4_6 (.CI(n40380), .I0(n35282), .I1(dti_counter[4]), 
            .CO(n40381));
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n40240), .I0(n2924), 
            .I1(VCC_net), .CO(n40241));
    SB_LUT4 dti_counter_2056_add_4_5_lut (.I0(n49678), .I1(n35282), .I2(dti_counter[3]), 
            .I3(n40379), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n40239), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n40239), .I0(n2925), 
            .I1(VCC_net), .CO(n40240));
    SB_CARRY dti_counter_2056_add_4_5 (.CI(n40379), .I0(n35282), .I1(dti_counter[3]), 
            .CO(n40380));
    SB_LUT4 i35814_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51252));
    defparam i35814_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n40238), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n40238), .I0(n2926), 
            .I1(VCC_net), .CO(n40239));
    SB_LUT4 unary_minus_10_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n40237), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n40237), .I0(n2927), 
            .I1(VCC_net), .CO(n40238));
    SB_LUT4 dti_counter_2056_add_4_4_lut (.I0(n49677), .I1(n35282), .I2(dti_counter[2]), 
            .I3(n40378), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n40236), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY dti_counter_2056_add_4_4 (.CI(n40378), .I0(n35282), .I1(dti_counter[2]), 
            .CO(n40379));
    SB_LUT4 dti_counter_2056_add_4_3_lut (.I0(n49676), .I1(n35282), .I2(dti_counter[1]), 
            .I3(n40377), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n40236), .I0(n2928), 
            .I1(VCC_net), .CO(n40237));
    SB_LUT4 encoder0_position_31__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_2056_add_4_3 (.CI(n40377), .I0(n35282), .I1(dti_counter[1]), 
            .CO(n40378));
    SB_LUT4 i35781_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51219));
    defparam i35781_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 dti_counter_2056_add_4_2_lut (.I0(n49662), .I1(n1910), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2056_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY dti_counter_2056_add_4_2 (.CI(VCC_net), .I0(n1910), .I1(dti_counter[0]), 
            .CO(n40377));
    SB_LUT4 i35749_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51187));
    defparam i35749_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n40235), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n40235), .I0(n2929), 
            .I1(GND_net), .CO(n40236));
    SB_LUT4 i35686_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51124));
    defparam i35686_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n40234), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29529_3_lut (.I0(n3), .I1(n7351), .I2(n44865), .I3(GND_net), 
            .O(n44880));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29530_3_lut (.I0(encoder0_position[30]), .I1(n44880), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i702_3_lut (.I0(n1027), .I1(n1094_adj_5169), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1313_rep_35_3_lut (.I0(n48682), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n48680));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1313_rep_35_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29515_3_lut (.I0(n5_adj_5150), .I1(n7353), .I2(n44865), .I3(GND_net), 
            .O(n44866));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n40234), .I0(n2930), 
            .I1(GND_net), .CO(n40235));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n40233), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n40233), .I0(n2931), 
            .I1(VCC_net), .CO(n40234));
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5214));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5213));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5211));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5210));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29516_3_lut (.I0(encoder0_position[28]), .I1(n44866), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5209));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096_adj_5171), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195_adj_5177), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFFESR GLA_181 (.Q(INLA_c_0), .C(CLK_c), .E(n29125), .D(GLA_N_384), 
            .R(n29460));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n40232), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5208));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5207));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dti_counter_2056__i0 (.Q(dti_counter[0]), .C(CLK_c), .D(n55));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5206));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5205));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7), .I2(encoder0_position[31]), .I3(GND_net), .O(n731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35629_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51067));
    defparam i35629_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n4_adj_5091), .I1(n5_adj_5150), .I2(n731), 
            .I3(n6_adj_5164), .O(n5_adj_5105));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'heeea;
    SB_CARRY add_224_5 (.CI(n39101), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n39102));
    SB_LUT4 i1_3_lut_adj_1719 (.I0(n3), .I1(n2), .I2(n5_adj_5105), .I3(GND_net), 
            .O(n44865));
    defparam i1_3_lut_adj_1719.LUT_INIT = 16'h8080;
    SB_LUT4 unary_minus_10_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_224_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n39114), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5204));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n40232), .I0(n2932), 
            .I1(GND_net), .CO(n40233));
    SB_CARRY add_224_18 (.CI(n39114), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n39115));
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n40231), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29537_3_lut (.I0(n6_adj_5164), .I1(n7354), .I2(n44865), .I3(GND_net), 
            .O(n44888));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2455_25_lut (.I0(n50760), .I1(n2_adj_5188), .I2(n1059), 
            .I3(n40368), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2455_24_lut (.I0(n50774), .I1(n2_adj_5188), .I2(n1158), 
            .I3(n40367), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n40231), .I0(n2933), 
            .I1(VCC_net), .CO(n40232));
    SB_CARRY add_2455_24 (.CI(n40367), .I0(n2_adj_5188), .I1(n1158), .CO(n40368));
    SB_LUT4 add_2455_23_lut (.I0(n50789), .I1(n2_adj_5188), .I2(n1257), 
            .I3(n40366), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_23 (.CI(n40366), .I0(n2_adj_5188), .I1(n1257), .CO(n40367));
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n40231));
    SB_LUT4 add_2455_22_lut (.I0(n50805), .I1(n2_adj_5188), .I2(n1356), 
            .I3(n40365), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i29538_3_lut (.I0(encoder0_position[27]), .I1(n44888), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097_adj_5172), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5203));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n51187), .I1(n2808), 
            .I2(VCC_net), .I3(n40230), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_2455_22 (.CI(n40365), .I0(n2_adj_5188), .I1(n1356), .CO(n40366));
    SB_LUT4 add_2455_21_lut (.I0(n50822), .I1(n2_adj_5188), .I2(n1455), 
            .I3(n40364), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_21 (.CI(n40364), .I0(n2_adj_5188), .I1(n1455), .CO(n40365));
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n40229), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_20_lut (.I0(n50840), .I1(n2_adj_5188), .I2(n1554), 
            .I3(n40363), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_20 (.CI(n40363), .I0(n2_adj_5188), .I1(n1554), .CO(n40364));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5202));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5201));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5200));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5199));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5198));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5197));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_2396_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n40914), 
            .O(n7350)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2396_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2396_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n40913), 
            .O(n7351)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2396_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2396_6 (.CI(n40913), .I0(n622), .I1(GND_net), .CO(n40914));
    SB_LUT4 add_2396_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n40912), 
            .O(n7352)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2396_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2396_5 (.CI(n40912), .I0(n623), .I1(VCC_net), .CO(n40913));
    SB_LUT4 add_2396_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n40911), 
            .O(n7353)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2396_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2396_4 (.CI(n40911), .I0(n516), .I1(GND_net), .CO(n40912));
    SB_LUT4 add_2396_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n40910), 
            .O(n7354)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2396_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2396_3 (.CI(n40910), .I0(n625), .I1(VCC_net), .CO(n40911));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5196));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2396_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7355)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2396_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2396_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n40910));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5195));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(CLK_c), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n2326), .I1(n2324), .I2(n2327), .I3(n2325), 
            .O(n47348));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5194));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5193));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5192));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5191));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(CLK_c), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5190));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5189));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_DFFSR pwm_setpoint_i23 (.Q(pwm_setpoint[23]), .C(CLK_c), .D(pwm_setpoint_23__N_191[23]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_23__N_11[22]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_23__N_11[21]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_23__N_11[20]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_23__N_11[19]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_23__N_11[18]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_23__N_11[17]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_23__N_11[16]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_23__N_11[15]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_23__N_11[14]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_23__N_11[13]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_23__N_11[12]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_23__N_11[11]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_23__N_11[10]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_23__N_11[9]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_23__N_11[8]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_23__N_11[7]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_23__N_11[6]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_23__N_11[5]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_23__N_11[4]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_23__N_11[3]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_23__N_11[2]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_23__N_11[1]));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 i1_3_lut_adj_1721 (.I0(n2322), .I1(n2328), .I2(n2323), .I3(GND_net), 
            .O(n47350));
    defparam i1_3_lut_adj_1721.LUT_INIT = 16'hfefe;
    SB_LUT4 i22807_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n36329));
    defparam i22807_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34673_3_lut (.I0(encoder0_position[26]), .I1(n44886), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098_adj_5173), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_adj_1722 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5107));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i2_2_lut_adj_1722.LUT_INIT = 16'heeee;
    SB_LUT4 i34966_3_lut (.I0(n2124), .I1(n2191), .I2(n2148), .I3(GND_net), 
            .O(n2223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34966_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2455_19_lut (.I0(n50863), .I1(n2_adj_5188), .I2(n1653_adj_5178), 
            .I3(n40362), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n40229), .I0(n2809), 
            .I1(VCC_net), .CO(n40230));
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n40228), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_19 (.CI(n40362), .I0(n2_adj_5188), .I1(n1653_adj_5178), 
            .CO(n40363));
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n40228), .I0(n2810), 
            .I1(VCC_net), .CO(n40229));
    SB_LUT4 add_2455_18_lut (.I0(n50883), .I1(n2_adj_5188), .I2(n1752), 
            .I3(n40361), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n40227), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_18 (.CI(n40361), .I0(n2_adj_5188), .I1(n1752), .CO(n40362));
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n40227), .I0(n2811), 
            .I1(VCC_net), .CO(n40228));
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n40226), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n40226), .I0(n2812), 
            .I1(VCC_net), .CO(n40227));
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n40225), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n40225), .I0(n2813), 
            .I1(VCC_net), .CO(n40226));
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n40224), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_17_lut (.I0(n50892), .I1(n2_adj_5188), .I2(n1851), 
            .I3(n40360), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n40224), .I0(n2814), 
            .I1(VCC_net), .CO(n40225));
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n40223), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_17 (.CI(n40360), .I0(n2_adj_5188), .I1(n1851), .CO(n40361));
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n40223), .I0(n2815), 
            .I1(VCC_net), .CO(n40224));
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n40222), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_16_lut (.I0(n50935), .I1(n2_adj_5188), .I2(n1950), 
            .I3(n40359), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_16 (.CI(n40359), .I0(n2_adj_5188), .I1(n1950), .CO(n40360));
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n40222), .I0(n2816), 
            .I1(VCC_net), .CO(n40223));
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n51067), .I1(n2412), 
            .I2(VCC_net), .I3(n39936), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2455_15_lut (.I0(n50961), .I1(n2_adj_5188), .I2(n2049), 
            .I3(n40358), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n39935), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n40221), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2455_15 (.CI(n40358), .I0(n2_adj_5188), .I1(n2049), .CO(n40359));
    SB_LUT4 add_2455_14_lut (.I0(n50987), .I1(n2_adj_5188), .I2(n2148), 
            .I3(n40357), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n40221), .I0(n2817), 
            .I1(VCC_net), .CO(n40222));
    SB_CARRY add_2455_14 (.CI(n40357), .I0(n2_adj_5188), .I1(n2148), .CO(n40358));
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n39935), .I0(n2413), 
            .I1(VCC_net), .CO(n39936));
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n39934), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n39100), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_13_lut (.I0(n51013), .I1(n2_adj_5188), .I2(n2247), 
            .I3(n40356), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_13 (.CI(n40356), .I0(n2_adj_5188), .I1(n2247), .CO(n40357));
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n39934), .I0(n2414), 
            .I1(VCC_net), .CO(n39935));
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n39933), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n39933), .I0(n2415), 
            .I1(VCC_net), .CO(n39934));
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n39932), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n39932), .I0(n2416), 
            .I1(VCC_net), .CO(n39933));
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n40220), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n39931), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n40220), .I0(n2818), 
            .I1(VCC_net), .CO(n40221));
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n40219), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n40219), .I0(n2819), 
            .I1(VCC_net), .CO(n40220));
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n40218), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n40218), .I0(n2820), 
            .I1(VCC_net), .CO(n40219));
    SB_LUT4 add_2455_12_lut (.I0(n51039), .I1(n2_adj_5188), .I2(n2346), 
            .I3(n40355), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n40217), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n39931), .I0(n2417), 
            .I1(VCC_net), .CO(n39932));
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n39930), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n39930), .I0(n2418), 
            .I1(VCC_net), .CO(n39931));
    SB_LUT4 add_224_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n39113), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n39929), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_4 (.CI(n39100), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n39101));
    SB_CARRY add_2455_12 (.CI(n40355), .I0(n2_adj_5188), .I1(n2346), .CO(n40356));
    SB_LUT4 add_2455_11_lut (.I0(n51067), .I1(n2_adj_5188), .I2(n2445), 
            .I3(n40354), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_11 (.CI(n40354), .I0(n2_adj_5188), .I1(n2445), .CO(n40355));
    SB_LUT4 add_2455_10_lut (.I0(n51071), .I1(n2_adj_5188), .I2(n2544), 
            .I3(n40353), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_10 (.CI(n40353), .I0(n2_adj_5188), .I1(n2544), .CO(n40354));
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n40217), .I0(n2821), 
            .I1(VCC_net), .CO(n40218));
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n39929), .I0(n2419), 
            .I1(VCC_net), .CO(n39930));
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n39928), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n40216), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_17 (.CI(n39113), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n39114));
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n40216), .I0(n2822), 
            .I1(VCC_net), .CO(n40217));
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n40215), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n2320), .I1(n2321), .I2(n47350), .I3(n47348), 
            .O(n47356));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n40215), .I0(n2823), 
            .I1(VCC_net), .CO(n40216));
    SB_LUT4 add_224_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n39099), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n40214), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_2455_9_lut (.I0(n51124), .I1(n2_adj_5188), .I2(n2643), 
            .I3(n40352), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_9 (.CI(n40352), .I0(n2_adj_5188), .I1(n2643), .CO(n40353));
    SB_LUT4 add_2455_8_lut (.I0(n51153), .I1(n2_adj_5188), .I2(n2742), 
            .I3(n40351), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_8 (.CI(n40351), .I0(n2_adj_5188), .I1(n2742), .CO(n40352));
    SB_LUT4 add_2455_7_lut (.I0(n51187), .I1(n2_adj_5188), .I2(n2841), 
            .I3(n40350), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_7 (.CI(n40350), .I0(n2_adj_5188), .I1(n2841), .CO(n40351));
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n40214), .I0(n2824), 
            .I1(VCC_net), .CO(n40215));
    SB_LUT4 add_2455_6_lut (.I0(n51219), .I1(n2_adj_5188), .I2(n2940), 
            .I3(n40349), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_6 (.CI(n40349), .I0(n2_adj_5188), .I1(n2940), .CO(n40350));
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n40213), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n39928), .I0(n2420), 
            .I1(VCC_net), .CO(n39929));
    SB_LUT4 add_2455_5_lut (.I0(n51252), .I1(n2_adj_5188), .I2(n3039), 
            .I3(n40348), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n40213), .I0(n2825), 
            .I1(VCC_net), .CO(n40214));
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n39927), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n40212), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n39927), .I0(n2421), 
            .I1(VCC_net), .CO(n39928));
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n39926), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n39926), .I0(n2422), 
            .I1(VCC_net), .CO(n39927));
    SB_CARRY add_2455_5 (.CI(n40348), .I0(n2_adj_5188), .I1(n3039), .CO(n40349));
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n40212), .I0(n2826), 
            .I1(VCC_net), .CO(n40213));
    SB_LUT4 i1_2_lut_adj_1724 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n47566));
    defparam i1_2_lut_adj_1724.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n39925), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_4_lut (.I0(n51286), .I1(n2_adj_5188), .I2(n3138), 
            .I3(n40347), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2455_4 (.CI(n40347), .I0(n2_adj_5188), .I1(n3138), .CO(n40348));
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n40211), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n40211), .I0(n2827), 
            .I1(VCC_net), .CO(n40212));
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n39925), .I0(n2423), 
            .I1(VCC_net), .CO(n39926));
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n39924), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n39924), .I0(n2424), 
            .I1(VCC_net), .CO(n39925));
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n39923), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n40210), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_3_lut (.I0(n51290), .I1(n2_adj_5188), .I2(n3237), 
            .I3(n40346), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n40210), .I0(n2828), 
            .I1(VCC_net), .CO(n40211));
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n1825), .I1(n1826), .I2(n1827), .I3(n1828), 
            .O(n47454));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n39597), .O(n1093_adj_5168)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n40209), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n39596), .O(n1094_adj_5169)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n39596), .I0(n1027), 
            .I1(VCC_net), .CO(n39597));
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n39595), .O(n1095_adj_5170)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n39923), .I0(n2425), 
            .I1(VCC_net), .CO(n39924));
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n39595), .I0(n1028), 
            .I1(VCC_net), .CO(n39596));
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n39594), .O(n1096_adj_5171)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n39922), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n39594), .I0(n1029), 
            .I1(GND_net), .CO(n39595));
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n39593), .O(n1097_adj_5172)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22685_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n36205));
    defparam i22685_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n39593), .I0(n1030), 
            .I1(GND_net), .CO(n39594));
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n39592), .O(n1098_adj_5173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1726 (.I0(n1823), .I1(n1824), .I2(n47454), .I3(GND_net), 
            .O(n47458));
    defparam i1_3_lut_adj_1726.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n39592), .I0(n1031), 
            .I1(VCC_net), .CO(n39593));
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n39591), .O(n1099_adj_5174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n39591), .I0(n1032), 
            .I1(GND_net), .CO(n39592));
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n1829), .I1(n36205), .I2(n1830), .I3(n1831), 
            .O(n45229));
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n39590), .O(n1100_adj_5175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n39590), .I0(n1033), 
            .I1(VCC_net), .CO(n39591));
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101_adj_5176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n39590));
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n1821), .I1(n1822), .I2(n45229), .I3(n47458), 
            .O(n47464));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_CARRY add_2455_3 (.CI(n40346), .I0(n2_adj_5188), .I1(n3237), .CO(n40347));
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n40209), .I0(n2829), 
            .I1(GND_net), .CO(n40210));
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n39922), .I0(n2426), 
            .I1(VCC_net), .CO(n39923));
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n39921), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n39112), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2455_2_lut (.I0(n51324), .I1(n2_adj_5188), .I2(n36493), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2455_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n40208), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n40208), .I0(n2830), 
            .I1(GND_net), .CO(n40209));
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n39921), .I0(n2427), 
            .I1(VCC_net), .CO(n39922));
    SB_CARRY add_224_16 (.CI(n39112), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n39113));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n39920), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n39920), .I0(n2428), 
            .I1(VCC_net), .CO(n39921));
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17_adj_5149), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n942));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16_adj_5151), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n941));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2455_2 (.CI(VCC_net), .I0(n2_adj_5188), .I1(n36493), 
            .CO(n40346));
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n40207), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n39919), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(n51290), .I1(n3204), 
            .I2(VCC_net), .I3(n40345), .O(n48576)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n40207), .I0(n2831), 
            .I1(VCC_net), .CO(n40208));
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n39919), .I0(n2429), 
            .I1(GND_net), .CO(n39920));
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n39918), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n40206), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n39111), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n40206), .I0(n2832), 
            .I1(GND_net), .CO(n40207));
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n39918), .I0(n2430), 
            .I1(GND_net), .CO(n39919));
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n39917), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_3 (.CI(n39099), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n39100));
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n39917), .I0(n2431), 
            .I1(VCC_net), .CO(n39918));
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n40344), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n40205), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n39916), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n39916), .I0(n2432), 
            .I1(GND_net), .CO(n39917));
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n40344), .I0(n3205), 
            .I1(VCC_net), .CO(n40345));
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n40205), .I0(n2833), 
            .I1(VCC_net), .CO(n40206));
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n40343), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n40343), .I0(n3206), 
            .I1(VCC_net), .CO(n40344));
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n40205));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n40342), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n39915), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n40342), .I0(n3207), 
            .I1(VCC_net), .CO(n40343));
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n39915), .I0(n2433), 
            .I1(VCC_net), .CO(n39916));
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(n51153), .I1(n2709), 
            .I2(VCC_net), .I3(n40204), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n40203), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n39915));
    SB_CARRY add_224_15 (.CI(n39111), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n39112));
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n40203), .I0(n2710), 
            .I1(VCC_net), .CO(n40204));
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n40341), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n40202), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n40341), .I0(n3208), 
            .I1(VCC_net), .CO(n40342));
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n40202), .I0(n2711), 
            .I1(VCC_net), .CO(n40203));
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n40340), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n40201), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n40201), .I0(n2712), 
            .I1(VCC_net), .CO(n40202));
    SB_LUT4 add_224_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n39110), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n47566), .I1(n2319), .I2(n47356), .I3(n36329), 
            .O(n47360));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hfefc;
    SB_LUT4 add_224_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_279), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_14 (.CI(n39110), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n39111));
    SB_CARRY add_224_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_279), 
            .CO(n39099));
    SB_LUT4 add_145_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n39098), .O(n1077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n39109), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n40340), .I0(n3209), 
            .I1(VCC_net), .CO(n40341));
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n40200), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n39097), .O(n1078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n51071), .I1(n2511), 
            .I2(VCC_net), .I3(n40055), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n40054), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n40200), .I0(n2713), 
            .I1(VCC_net), .CO(n40201));
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n40054), .I0(n2512), 
            .I1(VCC_net), .CO(n40055));
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n40339), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n40053), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n40199), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_13 (.CI(n39109), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n39110));
    SB_CARRY add_145_12 (.CI(n39077), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n39078));
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n40199), .I0(n2714), 
            .I1(VCC_net), .CO(n40200));
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n40339), .I0(n3210), 
            .I1(VCC_net), .CO(n40340));
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n40338), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n40198), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n40198), .I0(n2715), 
            .I1(VCC_net), .CO(n40199));
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n40053), .I0(n2513), 
            .I1(VCC_net), .CO(n40054));
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n40338), .I0(n3211), 
            .I1(VCC_net), .CO(n40339));
    SB_LUT4 add_224_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n39108), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n40337), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n40052), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n40052), .I0(n2514), 
            .I1(VCC_net), .CO(n40053));
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n40337), .I0(n3212), 
            .I1(VCC_net), .CO(n40338));
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n40197), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n40197), .I0(n2716), 
            .I1(VCC_net), .CO(n40198));
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n40051), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n39076), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n40051), .I0(n2515), 
            .I1(VCC_net), .CO(n40052));
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n40336), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n40050), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_32 (.CI(n39097), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n39098));
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n40336), .I0(n3213), 
            .I1(VCC_net), .CO(n40337));
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n40196), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n40050), .I0(n2516), 
            .I1(VCC_net), .CO(n40051));
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n40196), .I0(n2717), 
            .I1(VCC_net), .CO(n40197));
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n40049), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n40335), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n40195), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n40049), .I0(n2517), 
            .I1(VCC_net), .CO(n40050));
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n40195), .I0(n2718), 
            .I1(VCC_net), .CO(n40196));
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n40048), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n47360), 
            .O(n47366));
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n40048), .I0(n2518), 
            .I1(VCC_net), .CO(n40049));
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n51039), .I1(n2313), 
            .I2(VCC_net), .I3(n39903), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n40335), .I0(n3214), 
            .I1(VCC_net), .CO(n40336));
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n40194), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21632_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27826), .I3(n1195), .O(n35141));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i21632_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfbb;
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n40194), .I0(n2719), 
            .I1(VCC_net), .CO(n40195));
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n40047), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n39902), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n40334), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n39902), .I0(n2314), 
            .I1(VCC_net), .CO(n39903));
    SB_LUT4 add_145_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n39096), .O(n1079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n40334), .I0(n3215), 
            .I1(VCC_net), .CO(n40335));
    SB_CARRY add_145_31 (.CI(n39096), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n39097));
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n40193), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_12 (.CI(n39108), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n39109));
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n40333), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n40047), .I0(n2519), 
            .I1(VCC_net), .CO(n40048));
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n40333), .I0(n3216), 
            .I1(VCC_net), .CO(n40334));
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n40193), .I0(n2720), 
            .I1(VCC_net), .CO(n40194));
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n40192), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n40046), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n39901), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n39901), .I0(n2315), 
            .I1(VCC_net), .CO(n39902));
    SB_LUT4 i16096_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n43061), .I3(GND_net), .O(n29623));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16096_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n40046), .I0(n2520), 
            .I1(VCC_net), .CO(n40047));
    SB_LUT4 i16097_3_lut (.I0(h3), .I1(reg_B[0]), .I2(n46952), .I3(GND_net), 
            .O(n29624));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i16097_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n40332), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16098_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n29176), .I3(GND_net), .O(n29625));   // verilog/coms.v(127[12] 300[6])
    defparam i16098_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n40192), .I0(n2721), 
            .I1(VCC_net), .CO(n40193));
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n40045), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n39900), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27826), .I3(GND_net), .O(n27827));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 add_224_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n39107), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16099_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n29626));   // verilog/coms.v(127[12] 300[6])
    defparam i16099_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n40332), .I0(n3217), 
            .I1(VCC_net), .CO(n40333));
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n40191), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n40045), .I0(n2521), 
            .I1(VCC_net), .CO(n40046));
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n39900), .I0(n2316), 
            .I1(VCC_net), .CO(n39901));
    SB_LUT4 i16100_4_lut (.I0(state_7__N_4103[3]), .I1(data[5]), .I2(n4_adj_5133), 
            .I3(n28004), .O(n29627));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16100_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n40191), .I0(n2722), 
            .I1(VCC_net), .CO(n40192));
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n40044), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n39899), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n40044), .I0(n2522), 
            .I1(VCC_net), .CO(n40045));
    SB_CARRY add_224_9 (.CI(n39105), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n39106));
    SB_LUT4 i16101_4_lut (.I0(state_7__N_4103[3]), .I1(data[4]), .I2(n4_adj_5133), 
            .I3(n27984), .O(n29628));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16101_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n40331), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16102_4_lut (.I0(state_7__N_4103[3]), .I1(data[3]), .I2(n4), 
            .I3(n28004), .O(n29629));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16102_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n40190), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n40043), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_setpoint_23__I_0_i2_3_lut (.I0(duty[1]), .I1(pwm_setpoint_23__N_191[1]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[1]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n39899), .I0(n2317), 
            .I1(VCC_net), .CO(n39900));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27826), .I3(n1195), .O(n6969));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 add_224_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n39106), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n40331), .I0(n3218), 
            .I1(VCC_net), .CO(n40332));
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n40190), .I0(n2723), 
            .I1(VCC_net), .CO(n40191));
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n40189), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n40043), .I0(n2523), 
            .I1(VCC_net), .CO(n40044));
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n39898), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n39095), .O(n1080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35605_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n47366), 
            .O(n2346));
    defparam i35605_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 pwm_setpoint_23__I_0_i3_3_lut (.I0(duty[2]), .I1(pwm_setpoint_23__N_191[2]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[2]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16103_4_lut (.I0(state_7__N_4103[3]), .I1(data[2]), .I2(n4), 
            .I3(n27984), .O(n29630));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16103_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 pwm_setpoint_23__I_0_i4_3_lut (.I0(duty[3]), .I1(pwm_setpoint_23__N_191[3]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[3]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n27826), .I3(GND_net), .O(n6662));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n40042), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n39898), .I0(n2318), 
            .I1(VCC_net), .CO(n39899));
    SB_LUT4 pwm_setpoint_23__I_0_i5_3_lut (.I0(duty[4]), .I1(pwm_setpoint_23__N_191[4]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[4]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i6_3_lut (.I0(duty[5]), .I1(pwm_setpoint_23__N_191[5]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[5]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i7_3_lut (.I0(duty[6]), .I1(pwm_setpoint_23__N_191[6]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[6]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i8_3_lut (.I0(duty[7]), .I1(pwm_setpoint_23__N_191[7]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[7]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i9_3_lut (.I0(duty[8]), .I1(pwm_setpoint_23__N_191[8]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[8]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i10_3_lut (.I0(duty[9]), .I1(pwm_setpoint_23__N_191[9]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[9]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n40330), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_setpoint_23__I_0_i11_3_lut (.I0(duty[10]), .I1(pwm_setpoint_23__N_191[10]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[10]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n40189), .I0(n2724), 
            .I1(VCC_net), .CO(n40190));
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n40042), .I0(n2524), 
            .I1(VCC_net), .CO(n40043));
    SB_LUT4 pwm_setpoint_23__I_0_i12_3_lut (.I0(duty[11]), .I1(pwm_setpoint_23__N_191[11]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[11]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n39897), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_11 (.CI(n39076), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n39077));
    SB_LUT4 i16229_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n29176), .I3(GND_net), .O(n29756));   // verilog/coms.v(127[12] 300[6])
    defparam i16229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n40188), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n40041), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n39897), .I0(n2319), 
            .I1(VCC_net), .CO(n39898));
    SB_LUT4 add_145_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n39075), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_10 (.CI(n39106), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n39107));
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n39896), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_30 (.CI(n39095), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n39096));
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n40330), .I0(n3219), 
            .I1(VCC_net), .CO(n40331));
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n40188), .I0(n2725), 
            .I1(VCC_net), .CO(n40189));
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n40041), .I0(n2525), 
            .I1(VCC_net), .CO(n40042));
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n39896), .I0(n2320), 
            .I1(VCC_net), .CO(n39897));
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n40040), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n39895), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_10 (.CI(n39075), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n39076));
    SB_LUT4 pwm_setpoint_23__I_0_i13_3_lut (.I0(duty[12]), .I1(pwm_setpoint_23__N_191[12]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[12]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n40329), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_setpoint_23__I_0_i14_3_lut (.I0(duty[13]), .I1(pwm_setpoint_23__N_191[13]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[13]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i15_3_lut (.I0(duty[14]), .I1(pwm_setpoint_23__N_191[14]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[14]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i16_3_lut (.I0(duty[15]), .I1(pwm_setpoint_23__N_191[15]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[15]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i17_3_lut (.I0(duty[16]), .I1(pwm_setpoint_23__N_191[16]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[16]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i18_3_lut (.I0(duty[17]), .I1(pwm_setpoint_23__N_191[17]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[17]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n40329), .I0(n3220), 
            .I1(VCC_net), .CO(n40330));
    SB_LUT4 pwm_setpoint_23__I_0_i19_3_lut (.I0(duty[18]), .I1(pwm_setpoint_23__N_191[18]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[18]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_5 (.CI(n39070), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n39071));
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_setpoint_23__I_0_i20_3_lut (.I0(duty[19]), .I1(pwm_setpoint_23__N_191[19]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[19]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_145_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n39094), .O(n1081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_setpoint_23__I_0_i21_3_lut (.I0(duty[20]), .I1(pwm_setpoint_23__N_191[20]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[20]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i22_3_lut (.I0(duty[21]), .I1(pwm_setpoint_23__N_191[21]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[21]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 pwm_setpoint_23__I_0_i23_3_lut (.I0(duty[22]), .I1(pwm_setpoint_23__N_191[22]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[22]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n40187), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n40040), .I0(n2526), 
            .I1(VCC_net), .CO(n40041));
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n39895), .I0(n2321), 
            .I1(VCC_net), .CO(n39896));
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n40328), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n40187), .I0(n2726), 
            .I1(VCC_net), .CO(n40188));
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n39894), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n40186), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n40039), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n39894), .I0(n2322), 
            .I1(VCC_net), .CO(n39895));
    SB_CARRY add_145_29 (.CI(n39094), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n39095));
    SB_LUT4 add_145_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n39093), .O(n1082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16104_4_lut (.I0(state_7__N_4103[3]), .I1(data[1]), .I2(n10_adj_5222), 
            .I3(n28004), .O(n29631));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16104_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_10_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n40186), .I0(n2727), 
            .I1(VCC_net), .CO(n40187));
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n40039), .I0(n2527), 
            .I1(VCC_net), .CO(n40040));
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n39893), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n39893), .I0(n2323), 
            .I1(VCC_net), .CO(n39894));
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n40038), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n39892), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35479_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n47464), 
            .O(n1851));
    defparam i35479_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_10_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_215), 
            .I3(n39144), .O(pwm_setpoint_23__N_191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n3_adj_5095), 
            .I3(n39143), .O(pwm_setpoint_23__N_191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n39069), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n40328), .I0(n3221), 
            .I1(VCC_net), .CO(n40329));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n40185), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n40038), .I0(n2528), 
            .I1(VCC_net), .CO(n40039));
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n40037), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n40185), .I0(n2728), 
            .I1(VCC_net), .CO(n40186));
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n39892), .I0(n2324), 
            .I1(VCC_net), .CO(n39893));
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n39074), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_28 (.CI(n39093), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n39094));
    SB_CARRY add_145_4 (.CI(n39069), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n39070));
    SB_CARRY add_145_9 (.CI(n39074), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n39075));
    SB_CARRY unary_minus_10_add_3_24 (.CI(n39143), .I0(GND_net), .I1(n3_adj_5095), 
            .CO(n39144));
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n40327), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n40184), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n40037), .I0(n2529), 
            .I1(GND_net), .CO(n40038));
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n39891), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n40184), .I0(n2729), 
            .I1(GND_net), .CO(n40185));
    SB_LUT4 i22871_4_lut (.I0(n627), .I1(n831), .I2(n832), .I3(n833), 
            .O(n36393));
    defparam i22871_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 add_145_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n39092), .O(n1083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_27 (.CI(n39092), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n39093));
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n40036), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n39891), .I0(n2325), 
            .I1(VCC_net), .CO(n39892));
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n39890), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n39068), .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n39073), .O(n1102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_8 (.CI(n39073), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n39074));
    SB_LUT4 add_145_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n39091), .O(n1084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n40036), .I0(n2530), 
            .I1(GND_net), .CO(n40037));
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n39890), .I0(n2326), 
            .I1(VCC_net), .CO(n39891));
    SB_LUT4 add_145_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n39072), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n39889), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22979_4_lut (.I0(n829), .I1(n828), .I2(n36393), .I3(n830), 
            .O(n861));
    defparam i22979_4_lut.LUT_INIT = 16'heccc;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n40327), .I0(n3222), 
            .I1(VCC_net), .CO(n40328));
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n40183), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n40035), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n39889), .I0(n2327), 
            .I1(VCC_net), .CO(n39890));
    SB_CARRY add_145_26 (.CI(n39091), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n39092));
    SB_LUT4 unary_minus_10_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n4_adj_5096), 
            .I3(n39142), .O(pwm_setpoint_23__N_191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n40183), .I0(n2730), 
            .I1(GND_net), .CO(n40184));
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n40035), .I0(n2531), 
            .I1(VCC_net), .CO(n40036));
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n39888), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n39090), .O(n1085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_23 (.CI(n39142), .I0(GND_net), .I1(n4_adj_5096), 
            .CO(n39143));
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n40326), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n40182), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n40034), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n39888), .I0(n2328), 
            .I1(VCC_net), .CO(n39889));
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_25 (.CI(n39090), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n39091));
    SB_LUT4 add_145_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n39089), .O(n1086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n2424), .I1(n2427), .I2(n2422), .I3(n2425), 
            .O(n47512));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_DFFESR GLB_183 (.Q(INLB_c_0), .C(CLK_c), .E(n29125), .D(GLB_N_398), 
            .R(n29460));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFFESR GLC_185 (.Q(INLC_c_0), .C(CLK_c), .E(n29125), .D(GLC_N_412), 
            .R(n29460));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFF dti_counter_2056__i1 (.Q(dti_counter[1]), .C(CLK_c), .D(n54));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF read_189 (.Q(read), .C(CLK_c), .D(n46975));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 unary_minus_10_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n5), 
            .I3(n39141), .O(pwm_setpoint_23__N_191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n40182), .I0(n2731), 
            .I1(VCC_net), .CO(n40183));
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n40034), .I0(n2532), 
            .I1(GND_net), .CO(n40035));
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n39887), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n40326), .I0(n3223), 
            .I1(VCC_net), .CO(n40327));
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n40181), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n40033), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n39887), .I0(n2329), 
            .I1(GND_net), .CO(n39888));
    SB_CARRY add_145_3 (.CI(n39068), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n39069));
    SB_CARRY unary_minus_10_add_3_22 (.CI(n39141), .I0(GND_net), .I1(n5), 
            .CO(n39142));
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n40181), .I0(n2732), 
            .I1(GND_net), .CO(n40182));
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n40033), .I0(n2533), 
            .I1(VCC_net), .CO(n40034));
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n39886), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_24 (.CI(n39089), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n39090));
    SB_CARRY add_145_7 (.CI(n39072), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n39073));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n40325), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n40180), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n39886), .I0(n2330), 
            .I1(GND_net), .CO(n39887));
    SB_LUT4 add_145_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n39088), .O(n1087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_23 (.CI(n39088), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n39089));
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n40325), .I0(n3224), 
            .I1(VCC_net), .CO(n40326));
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n40180), .I0(n2733), 
            .I1(VCC_net), .CO(n40181));
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n40033));
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n39885), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n39087), .O(n1088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n6), 
            .I3(n39140), .O(pwm_setpoint_23__N_191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n39885), .I0(n2331), 
            .I1(VCC_net), .CO(n39886));
    SB_CARRY unary_minus_10_add_3_21 (.CI(n39140), .I0(GND_net), .I1(n6), 
            .CO(n39141));
    SB_LUT4 unary_minus_10_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n7_adj_5097), 
            .I3(n39139), .O(pwm_setpoint_23__N_191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_20 (.CI(n39139), .I0(GND_net), .I1(n7_adj_5097), 
            .CO(n39140));
    SB_LUT4 unary_minus_10_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n8), 
            .I3(n39138), .O(pwm_setpoint_23__N_191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_5167), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n1927), .I1(n1926), .I2(n1925), .I3(n1928), 
            .O(n47268));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22867_4_lut (.I0(n628), .I1(n931), .I2(n932), .I3(n933), 
            .O(n36389));
    defparam i22867_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22683_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n36203));
    defparam i22683_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1733 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n47376));
    defparam i1_2_lut_adj_1733.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(n1922), .I1(n1923), .I2(n47268), .I3(n1924), 
            .O(n47274));
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 pwm_setpoint_23__I_0_i1_3_lut (.I0(duty[0]), .I1(pwm_setpoint_23__N_191[0]), 
            .I2(duty[23]), .I3(GND_net), .O(pwm_setpoint_23__N_11[0]));   // verilog/TinyFPGA_B.v(110[13] 113[7])
    defparam pwm_setpoint_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n927), .I1(n47376), .I2(n928), .I3(n36389), 
            .O(n960));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n1929), .I1(n36203), .I2(n1930), .I3(n1931), 
            .O(n45214));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i573_3_lut (.I0(n627), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n1920), .I1(n45214), .I2(n1921), .I3(n47274), 
            .O(n47280));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i1_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i2_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i3_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i4_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i5_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i6_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i7_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22755_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n36277));
    defparam i22755_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i35503_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n47280), 
            .O(n1950));
    defparam i35503_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i8_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i9_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), .I2(motor_state_23__N_123[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n2428), .I1(n47512), .I2(n2426), .I3(n2423), 
            .O(n47514));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hfffe;
    SB_LUT4 i22803_4_lut (.I0(n949), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n36325));
    defparam i22803_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n2419), .I1(n2420), .I2(n47514), .I3(n2421), 
            .O(n47520));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1740 (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n47744));
    defparam i1_2_lut_adj_1740.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n2418), .I1(n47744), .I2(n47520), .I3(n36325), 
            .O(n47524));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n40324), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n40180));
    SB_LUT4 i1_4_lut_adj_1742 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n47524), 
            .O(n47530));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i35632_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n47530), 
            .O(n2445));
    defparam i35632_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n2528), .I1(n2525), .I2(n2526), .I3(n2523), 
            .O(n47142));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n2521), .I1(n47142), .I2(n2527), .I3(n2524), 
            .O(n47146));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'hfffe;
    SB_LUT4 i22623_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n36141));
    defparam i22623_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n2529), .I1(n36141), .I2(n2530), .I3(n2531), 
            .O(n45246));
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1746 (.I0(n2516), .I1(n45246), .I2(n2518), .I3(n2522), 
            .O(n47392));
    defparam i1_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(n2517), .I1(n2519), .I2(n2520), .I3(n47146), 
            .O(n47152));
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n2514), .I1(n2513), .I2(n2515), .I3(n47392), 
            .O(n46745));
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 i35660_4_lut (.I0(n2512), .I1(n2511), .I2(n46745), .I3(n47152), 
            .O(n2544));
    defparam i35660_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1661_rep_20_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1661_rep_20_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i10_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(GND_net), .I1(n2610), 
            .I2(VCC_net), .I3(n40179), .O(n2677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i11_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i12_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i13_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(CLK_c), .D(n43957));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n43275));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n29684));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n39884), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_19 (.CI(n39138), .I0(GND_net), .I1(n8), 
            .CO(n39139));
    SB_LUT4 encoder0_position_31__I_0_i1717_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1717_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i14_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1749 (.I0(n1029), .I1(n36277), .I2(n1030), .I3(n1031), 
            .O(n45172));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n39884), .I0(n2332), 
            .I1(GND_net), .CO(n39885));
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i15_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i16_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i17_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i18_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i19_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n40324), .I0(n3225), 
            .I1(VCC_net), .CO(n40325));
    SB_LUT4 mux_236_i20_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n40178), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1792_rep_16_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1792_rep_16_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34886_3_lut (.I0(n2827), .I1(n2894), .I2(n2841), .I3(GND_net), 
            .O(n2926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n39883), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i21_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(CLK_c), .D(n44909));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 mux_236_i22_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i23_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 unary_minus_10_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n9), 
            .I3(n39137), .O(pwm_setpoint_23__N_191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_18 (.CI(n39137), .I0(GND_net), .I1(n9), 
            .CO(n39138));
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22681_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n36201));
    defparam i22681_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1750 (.I0(n2026), .I1(n2027), .I2(GND_net), .I3(GND_net), 
            .O(n47478));
    defparam i1_2_lut_adj_1750.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n39447), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1751 (.I0(n2025), .I1(n47478), .I2(n2024), .I3(n2028), 
            .O(n47482));
    defparam i1_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n39446), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n2029), .I1(n36201), .I2(n2030), .I3(n2031), 
            .O(n45250));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n47482), 
            .O(n47488));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n2019), .I1(n2020), .I2(n47488), .I3(n45250), 
            .O(n47494));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n39446), .I0(n928), 
            .I1(VCC_net), .CO(n39447));
    SB_LUT4 i35527_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n47494), 
            .O(n2049));
    defparam i35527_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n39445), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n39445), .I0(n929), 
            .I1(GND_net), .CO(n39446));
    SB_LUT4 mux_236_i24_3_lut_4_lut (.I0(n27828), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n39444), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n39444), .I0(n930), 
            .I1(GND_net), .CO(n39445));
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n39443), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n39443), .I0(n931), 
            .I1(VCC_net), .CO(n39444));
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n39442), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n39442), .I0(n932), 
            .I1(GND_net), .CO(n39443));
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n39441), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21_adj_5145), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n946));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n39441), .I0(n933), 
            .I1(VCC_net), .CO(n39442));
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n628), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1755 (.I0(n2126), .I1(n2127), .I2(n2125), .I3(GND_net), 
            .O(n47198));
    defparam i1_3_lut_adj_1755.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n628), 
            .I1(GND_net), .CO(n39441));
    SB_LUT4 i1_3_lut_adj_1756 (.I0(n2123), .I1(n2128), .I2(n2124), .I3(GND_net), 
            .O(n47200));
    defparam i1_3_lut_adj_1756.LUT_INIT = 16'hfefe;
    SB_LUT4 i22815_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n36337));
    defparam i22815_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1757 (.I0(n2121), .I1(n2122), .I2(n47200), .I3(n47198), 
            .O(n47206));
    defparam i1_4_lut_adj_1757.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n2129), .I1(n47206), .I2(n36337), .I3(n2130), 
            .O(n47208));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n2118), .I1(n2119), .I2(n47208), .I3(n2120), 
            .O(n47214));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i35554_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n47214), 
            .O(n2148));
    defparam i35554_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6657_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_403));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6657_3_lut_4_lut.LUT_INIT = 16'haa1c;
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n39430), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n39429), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n39429), .I0(n829), 
            .I1(GND_net), .CO(n39430));
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n39428), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n39428), .I0(n830), 
            .I1(GND_net), .CO(n39429));
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n39427), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n39427), .I0(n831), 
            .I1(VCC_net), .CO(n39428));
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n39426), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n39426), .I0(n832), 
            .I1(GND_net), .CO(n39427));
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n39425), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n39425), .I0(n833), 
            .I1(VCC_net), .CO(n39426));
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n627), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n627), 
            .I1(GND_net), .CO(n39425));
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n29938));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n29937));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n29936));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n29935));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n29934));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n29933));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n40323), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i6659_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_412));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6659_3_lut_4_lut.LUT_INIT = 16'h1caa;
    SB_LUT4 i6653_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHB_N_389));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6653_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_LUT4 encoder0_position_31__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6655_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLB_N_398));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i6655_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n40178), .I0(n2611), 
            .I1(VCC_net), .CO(n40179));
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n39883), .I0(n2333), 
            .I1(VCC_net), .CO(n39884));
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n29932));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(h1), .I1(h3), .I2(h2), .I3(GND_net), 
            .O(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n40177), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n10_adj_5098), 
            .I3(n39136), .O(pwm_setpoint_23__N_191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF dti_counter_2056__i2 (.Q(dti_counter[2]), .C(CLK_c), .D(n53));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n39883));
    SB_LUT4 i35325_4_lut (.I0(n1026), .I1(n45172), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i35325_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dti_counter_2056__i3 (.Q(dti_counter[3]), .C(CLK_c), .D(n52));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i4 (.Q(dti_counter[4]), .C(CLK_c), .D(n51));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i5 (.Q(dti_counter[5]), .C(CLK_c), .D(n50));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i6 (.Q(dti_counter[6]), .C(CLK_c), .D(n49));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2056__i7 (.Q(dti_counter[7]), .C(CLK_c), .D(n48));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n29655));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(CLK_c), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n40323), .I0(n3226), 
            .I1(VCC_net), .CO(n40324));
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n40177), .I0(n2612), 
            .I1(VCC_net), .CO(n40178));
    SB_LUT4 i22857_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n36379));
    defparam i22857_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5188), .I3(n40590), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5189), .I3(n40589), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n40589), 
            .I0(GND_net), .I1(n3_adj_5189), .CO(n40590));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5190), .I3(n40588), .O(n4_adj_5091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n40588), 
            .I0(GND_net), .I1(n4_adj_5190), .CO(n40589));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5191), .I3(n40587), .O(n5_adj_5150)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n40587), 
            .I0(GND_net), .I1(n5_adj_5191), .CO(n40588));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5192), .I3(n40586), .O(n6_adj_5164)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n40586), 
            .I0(GND_net), .I1(n6_adj_5192), .CO(n40587));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5193), .I3(n40585), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n40585), 
            .I0(GND_net), .I1(n7_adj_5193), .CO(n40586));
    SB_CARRY unary_minus_10_add_3_17 (.CI(n39136), .I0(GND_net), .I1(n10_adj_5098), 
            .CO(n39137));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5194), .I3(n40584), .O(n8_adj_5167)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n40584), 
            .I0(GND_net), .I1(n8_adj_5194), .CO(n40585));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5195), .I3(n40583), .O(n9_adj_5166)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n40322), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n40583), 
            .I0(GND_net), .I1(n9_adj_5195), .CO(n40584));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5196), .I3(n40582), .O(n10_adj_5165)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n40582), 
            .I0(GND_net), .I1(n10_adj_5196), .CO(n40583));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5197), .I3(n40581), .O(n11_adj_5157)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n40581), 
            .I0(GND_net), .I1(n11_adj_5197), .CO(n40582));
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n40322), .I0(n3227), 
            .I1(VCC_net), .CO(n40323));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5198), .I3(n40580), .O(n12_adj_5156)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n40176), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n40580), 
            .I0(GND_net), .I1(n12_adj_5198), .CO(n40581));
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n40176), .I0(n2613), 
            .I1(VCC_net), .CO(n40177));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5199), .I3(n40579), .O(n13_adj_5155)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n40579), 
            .I0(GND_net), .I1(n13_adj_5199), .CO(n40580));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5200), .I3(n40578), .O(n14_adj_5154)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n40578), 
            .I0(GND_net), .I1(n14_adj_5200), .CO(n40579));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5201), .I3(n40577), .O(n15_adj_5153)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n40321), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n40577), 
            .I0(GND_net), .I1(n15_adj_5201), .CO(n40578));
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n40175), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5202), .I3(n40576), .O(n16_adj_5151)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n40576), 
            .I0(GND_net), .I1(n16_adj_5202), .CO(n40577));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5203), .I3(n40575), .O(n17_adj_5149)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n40575), 
            .I0(GND_net), .I1(n17_adj_5203), .CO(n40576));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5204), .I3(n40574), .O(n18_adj_5148)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11), 
            .I3(n39135), .O(pwm_setpoint_23__N_191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n40574), 
            .I0(GND_net), .I1(n18_adj_5204), .CO(n40575));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5205), .I3(n40573), .O(n19_adj_5147)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n40573), 
            .I0(GND_net), .I1(n19_adj_5205), .CO(n40574));
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5206), .I3(n40572), .O(n20_adj_5146)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n40572), 
            .I0(GND_net), .I1(n20_adj_5206), .CO(n40573));
    SB_CARRY add_145_22 (.CI(n39087), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n39088));
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n40175), .I0(n2614), 
            .I1(VCC_net), .CO(n40176));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5207), .I3(n40571), .O(n21_adj_5145)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n40321), .I0(n3228), 
            .I1(VCC_net), .CO(n40322));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n40571), 
            .I0(GND_net), .I1(n21_adj_5207), .CO(n40572));
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n40174), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5208), .I3(n40570), .O(n22_adj_5144)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n40570), 
            .I0(GND_net), .I1(n22_adj_5208), .CO(n40571));
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5209), .I3(n40569), .O(n23_adj_5143)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n40569), 
            .I0(GND_net), .I1(n23_adj_5209), .CO(n40570));
    SB_LUT4 encoder0_position_31__I_0_i1790_rep_15_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1790_rep_15_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5210), .I3(n40568), .O(n24_adj_5142)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n40568), 
            .I0(GND_net), .I1(n24_adj_5210), .CO(n40569));
    SB_LUT4 i34884_3_lut (.I0(n2825), .I1(n2892), .I2(n2841), .I3(GND_net), 
            .O(n2924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5211), .I3(n40567), .O(n25_adj_5141)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n40567), 
            .I0(GND_net), .I1(n25_adj_5211), .CO(n40568));
    SB_LUT4 encoder0_position_31__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5212), .I3(n40566), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n40566), 
            .I0(GND_net), .I1(n26_adj_5212), .CO(n40567));
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n40174), .I0(n2615), 
            .I1(VCC_net), .CO(n40175));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5213), .I3(n40565), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n40565), 
            .I0(GND_net), .I1(n27_adj_5213), .CO(n40566));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5214), .I3(n40564), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n40320), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n40173), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n40564), 
            .I0(GND_net), .I1(n28_adj_5214), .CO(n40565));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5215), .I3(n40563), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n40563), 
            .I0(GND_net), .I1(n29_adj_5215), .CO(n40564));
    SB_LUT4 encoder0_position_31__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_16 (.CI(n39135), .I0(GND_net), .I1(n11), 
            .CO(n39136));
    SB_LUT4 encoder0_position_31__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5216), .I3(n40562), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n40562), 
            .I0(GND_net), .I1(n30_adj_5216), .CO(n40563));
    SB_LUT4 add_145_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n39086), .O(n1089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5217), .I3(n40561), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n40561), 
            .I0(GND_net), .I1(n31_adj_5217), .CO(n40562));
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n40320), .I0(n3229), 
            .I1(GND_net), .CO(n40321));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5218), .I3(n40560), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n40173), .I0(n2616), 
            .I1(VCC_net), .CO(n40174));
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n40560), 
            .I0(GND_net), .I1(n32_adj_5218), .CO(n40561));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5219), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5219), .CO(n40560));
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12), 
            .I3(n39134), .O(pwm_setpoint_23__N_191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n40319), .O(n49621)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n39071), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n40172), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1760 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n47222));
    defparam i1_3_lut_adj_1760.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n39863), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_21 (.CI(n39086), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n39087));
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n40319), .I0(n3230), 
            .I1(GND_net), .CO(n40320));
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n40172), .I0(n2617), 
            .I1(VCC_net), .CO(n40173));
    SB_LUT4 add_145_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n39085), .O(n1090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1761 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n47386));
    defparam i1_2_lut_adj_1761.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n40318), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n40171), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_15 (.CI(n39134), .I0(GND_net), .I1(n12), 
            .CO(n39135));
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n40171), .I0(n2618), 
            .I1(VCC_net), .CO(n40172));
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_20 (.CI(n39085), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n39086));
    SB_LUT4 unary_minus_10_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n13), 
            .I3(n39133), .O(pwm_setpoint_23__N_191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_14 (.CI(n39133), .I0(GND_net), .I1(n13), 
            .CO(n39134));
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n40318), .I0(n3231), 
            .I1(VCC_net), .CO(n40319));
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n40170), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n40317), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n40170), .I0(n2619), 
            .I1(VCC_net), .CO(n40171));
    SB_LUT4 i22889_4_lut (.I0(n951), .I1(n2631), .I2(n2632), .I3(n2633), 
            .O(n36411));
    defparam i22889_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i35339_4_lut (.I0(n47386), .I1(n1125), .I2(n47222), .I3(n36379), 
            .O(n1158));
    defparam i35339_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n2619), .I1(n2627), .I2(n2625), .I3(n2623), 
            .O(n47574));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n40169), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5099), 
            .I3(n39132), .O(pwm_setpoint_23__N_191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n39084), .O(n1091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n2629), .I1(n47574), .I2(n36411), .I3(n2630), 
            .O(n47576));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'heccc;
    SB_CARRY add_145_19 (.CI(n39084), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n39085));
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n2615), .I1(n2616), .I2(n2617), .I3(n47576), 
            .O(n47582));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1765 (.I0(n2624), .I1(n2622), .I2(GND_net), .I3(GND_net), 
            .O(n47594));
    defparam i1_2_lut_adj_1765.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1766 (.I0(n2626), .I1(n2621), .I2(n2628), .I3(GND_net), 
            .O(n47596));
    defparam i1_3_lut_adj_1766.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n2612), .I1(n2613), .I2(n2614), .I3(n47582), 
            .O(n47588));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 add_145_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n39083), .O(n1092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n2618), .I1(n2620), .I2(n47596), .I3(n47594), 
            .O(n47602));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'hfffe;
    SB_CARRY add_145_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n39068));
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n40317), .I0(n3232), 
            .I1(GND_net), .CO(n40318));
    SB_LUT4 i35689_4_lut (.I0(n2610), .I1(n47602), .I2(n47588), .I3(n2611), 
            .O(n2643));
    defparam i35689_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n40169), .I0(n2620), 
            .I1(VCC_net), .CO(n40170));
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22789_3_lut (.I0(n952), .I1(n2732), .I2(n2733), .I3(GND_net), 
            .O(n36311));
    defparam i22789_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1769 (.I0(n2725), .I1(n2720), .I2(n2727), .I3(GND_net), 
            .O(n47234));
    defparam i1_3_lut_adj_1769.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(n2723), .I1(n2721), .I2(n2726), .I3(n2728), 
            .O(n47236));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(n47236), .I1(n47234), .I2(n2722), .I3(n2724), 
            .O(n47240));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n40316), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n40168), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_13 (.CI(n39132), .I0(GND_net), .I1(n14_adj_5099), 
            .CO(n39133));
    SB_CARRY add_145_18 (.CI(n39083), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n39084));
    SB_LUT4 add_145_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n39082), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n40168), .I0(n2621), 
            .I1(VCC_net), .CO(n40169));
    SB_CARRY add_145_6 (.CI(n39071), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n39072));
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n2729), .I1(n36311), .I2(n2730), .I3(n2731), 
            .O(n45252));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'ha080;
    SB_LUT4 unary_minus_10_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15), 
            .I3(n39131), .O(pwm_setpoint_23__N_191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_17 (.CI(n39082), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n39083));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_5164), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5_adj_5150), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n516));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_5091), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3), .I2(encoder0_position[31]), .I3(GND_net), .O(n622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2_adj_5104), .I3(n39371), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4895_2_lut (.I0(n2), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4895_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n2717), .I1(n2718), .I2(n47240), .I3(n2719), 
            .O(n47246));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5131), .I3(n39370), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n39370), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5131), .CO(n39371));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5130), .I3(n39369), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n40316), .I0(n3233), 
            .I1(VCC_net), .CO(n40317));
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n40167), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n39081), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n39369), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5130), .CO(n39370));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5129), .I3(n39368), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n39368), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5129), .CO(n39369));
    SB_CARRY add_145_16 (.CI(n39081), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n39082));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5128), .I3(n39367), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n39367), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5128), .CO(n39368));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5127), .I3(n39366), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n39366), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5127), .CO(n39367));
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n2715), .I1(n2716), .I2(n47246), .I3(n45252), 
            .O(n47252));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099_adj_5174), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n47252), 
            .O(n47258));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 i35721_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n47258), 
            .O(n2742));
    defparam i35721_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5126), .I3(n39365), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n39365), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5126), .CO(n39366));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5125), .I3(n39364), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n39364), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5125), .CO(n39365));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5124), .I3(n39363), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_12 (.CI(n39131), .I0(GND_net), .I1(n15), 
            .CO(n39132));
    SB_LUT4 unary_minus_10_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16), 
            .I3(n39130), .O(pwm_setpoint_23__N_191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_11_lut.LUT_INIT = 16'hC33C;
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.n1653(CLK_c), .ENCODER0_B_N_keep(ENCODER0_B_N), 
            .ENCODER0_A_N_keep(ENCODER0_A_N), .\a_new[1] (a_new[1]), .b_prev(b_prev), 
            .n29689(n29689), .n1617(n1617), .direction_N_3907(direction_N_3907), 
            .encoder0_position({encoder0_position}), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(285[57] 292[6])
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n39363), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5124), .CO(n39364));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5123), .I3(n39362), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n39362), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5123), .CO(n39363));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5122), .I3(n39361), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n39361), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5122), .CO(n39362));
    SB_LUT4 i1_3_lut_adj_1776 (.I0(n2822), .I1(n2820), .I2(n2826), .I3(GND_net), 
            .O(n47614));
    defparam i1_3_lut_adj_1776.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5121), .I3(n39360), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n2828), .I1(n2823), .I2(n2825), .I3(n2827), 
            .O(n47616));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_CARRY unary_minus_10_add_3_11 (.CI(n39130), .I0(GND_net), .I1(n16), 
            .CO(n39131));
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n47616), .I1(n47614), .I2(n2824), .I3(n2821), 
            .O(n47620));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_10_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17), 
            .I3(n39129), .O(pwm_setpoint_23__N_191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n39360), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5121), .CO(n39361));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5120), .I3(n39359), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n39359), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5120), .CO(n39360));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5119), .I3(n39358), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n39358), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5119), .CO(n39359));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5118), .I3(n39357), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n39357), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5118), .CO(n39358));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5117), .I3(n39356), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n40315), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n39356), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5117), .CO(n39357));
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n40167), .I0(n2622), 
            .I1(VCC_net), .CO(n40168));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5116), .I3(n39355), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n39355), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5116), .CO(n39356));
    SB_LUT4 i22885_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n36407));
    defparam i22885_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n2817), .I1(n2818), .I2(n47620), .I3(n2819), 
            .O(n47626));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5115), .I3(n39354), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n47626), .I1(n2829), .I2(n36407), .I3(n2830), 
            .O(n47628));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'heaaa;
    SB_CARRY unary_minus_10_add_3_10 (.CI(n39129), .I0(GND_net), .I1(n17), 
            .CO(n39130));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n39354), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5115), .CO(n39355));
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n47628), 
            .O(n47634));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n47634), 
            .O(n47640));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'hfffe;
    SB_LUT4 i35752_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n47640), 
            .O(n2841));
    defparam i35752_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n40315), .I0(n957), 
            .I1(GND_net), .CO(n40316));
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5114), .I3(n39353), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n39353), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5114), .CO(n39354));
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n40166), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18), 
            .I3(n39128), .O(pwm_setpoint_23__N_191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5113), .I3(n39352), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n39352), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5113), .CO(n39353));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5112), .I3(n39351), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n40166), .I0(n2623), 
            .I1(VCC_net), .CO(n40167));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n39351), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5112), .CO(n39352));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5111), .I3(n39350), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n39080), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n39350), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5111), .CO(n39351));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5110), .I3(n39349), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n39349), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5110), .CO(n39350));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5109), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5109), .CO(n39349));
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n40165), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_15 (.CI(n39080), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n39081));
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n652), 
            .I1(VCC_net), .CO(n40315));
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n51286), .I1(n3105), 
            .I2(VCC_net), .I3(n40314), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n40165), .I0(n2624), 
            .I1(VCC_net), .CO(n40166));
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n40164), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35402_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50840));
    defparam i35402_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n40164), .I0(n2625), 
            .I1(VCC_net), .CO(n40165));
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n40163), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n39079), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n40313), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_9 (.CI(n39128), .I0(GND_net), .I1(n18), 
            .CO(n39129));
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n40163), .I0(n2626), 
            .I1(VCC_net), .CO(n40164));
    SB_CARRY add_145_14 (.CI(n39079), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n39080));
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1783 (.I0(n2922), .I1(n2926), .I2(GND_net), .I3(GND_net), 
            .O(n47162));
    defparam i1_2_lut_adj_1783.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n2928), .I1(n2925), .I2(n2927), .I3(n2920), 
            .O(n47166));
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 i22785_3_lut (.I0(n954), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n36307));
    defparam i22785_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n40313), .I0(n3106), 
            .I1(VCC_net), .CO(n40314));
    SB_LUT4 i1_4_lut_adj_1785 (.I0(n2919), .I1(n47166), .I2(n47162), .I3(n2924), 
            .O(n47170));
    defparam i1_4_lut_adj_1785.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n2929), .I1(n36307), .I2(n2930), .I3(n2931), 
            .O(n45266));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n2916), .I1(n2917), .I2(n2918), .I3(n47170), 
            .O(n47176));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n2913), .I1(n2915), .I2(n47176), .I3(n45266), 
            .O(n47182));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n2914), .I1(n2912), .I2(n2923), .I3(n2921), 
            .O(n46565));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n2910), .I1(n46565), .I2(n2911), .I3(n47182), 
            .O(n47188));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hfffe;
    SB_LUT4 i35784_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n47188), 
            .O(n2940));
    defparam i35784_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n40162), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19), 
            .I3(n39127), .O(pwm_setpoint_23__N_191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n40162), .I0(n2627), 
            .I1(VCC_net), .CO(n40163));
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n39104), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n39866), .I0(n2220), 
            .I1(VCC_net), .CO(n39867));
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22714_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n36235));
    defparam i22714_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY unary_minus_10_add_3_8 (.CI(n39127), .I0(GND_net), .I1(n19), 
            .CO(n39128));
    SB_LUT4 unary_minus_10_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20), 
            .I3(n39126), .O(pwm_setpoint_23__N_191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n3020), .I1(n3021), .I2(n3024), .I3(n3022), 
            .O(n47660));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n40161), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n40161), .I0(n2628), 
            .I1(VCC_net), .CO(n40162));
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n40312), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1792 (.I0(n3028), .I1(n3019), .I2(n3023), .I3(GND_net), 
            .O(n47658));
    defparam i1_3_lut_adj_1792.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(n3016), .I1(n3017), .I2(n3018), .I3(n3026), 
            .O(n47684));
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n40160), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1794 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n47400));
    defparam i1_3_lut_adj_1794.LUT_INIT = 16'hfefe;
    SB_LUT4 i22781_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n36303));
    defparam i22781_3_lut.LUT_INIT = 16'hc8c8;
    GND i1 (.Y(GND_net));
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n47658), .I1(n47660), .I2(n3027), .I3(n3025), 
            .O(n47664));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n3029), .I1(n36303), .I2(n3030), .I3(n3031), 
            .O(n45315));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n40312), .I0(n3107), 
            .I1(VCC_net), .CO(n40313));
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n40311), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n40160), .I0(n2629), 
            .I1(GND_net), .CO(n40161));
    SB_CARRY unary_minus_10_add_3_7 (.CI(n39126), .I0(GND_net), .I1(n20), 
            .CO(n39127));
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n40311), .I0(n3108), 
            .I1(VCC_net), .CO(n40312));
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n40159), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21), 
            .I3(n39125), .O(pwm_setpoint_23__N_191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n40159), .I0(n2630), 
            .I1(GND_net), .CO(n40160));
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n40158), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n39864), .I0(n2222), 
            .I1(VCC_net), .CO(n39865));
    SB_CARRY unary_minus_10_add_3_6 (.CI(n39125), .I0(GND_net), .I1(n21), 
            .CO(n39126));
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n40310), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n39864), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n40158), .I0(n2631), 
            .I1(VCC_net), .CO(n40159));
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n40310), .I0(n3109), 
            .I1(VCC_net), .CO(n40311));
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n40157), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n40309), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n3013), .I1(n3015), .I2(n45315), .I3(n47664), 
            .O(n47670));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(n3008), .I1(n3010), .I2(n3014), .I3(n47684), 
            .O(n47690));
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n3009), .I1(n3011), .I2(n3012), .I3(n47670), 
            .O(n47676));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 i35817_4_lut (.I0(n3006), .I1(n47676), .I2(n47690), .I3(n3007), 
            .O(n3039));
    defparam i35817_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24_adj_5142), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n949));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_5165), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n935));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i709_3_lut (.I0(n935), .I1(n1101_adj_5176), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n1229), .I1(n36235), .I2(n1230), .I3(n1231), 
            .O(n45167));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16117_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5152), 
            .I3(n27971), .O(n29644));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16117_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35354_4_lut (.I0(n1225), .I1(n1224), .I2(n45167), .I3(n47400), 
            .O(n1257));
    defparam i35354_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1111_rep_52_3_lut (.I0(n1695), .I1(n1794), 
            .I2(n1752), .I3(GND_net), .O(n48697));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1111_rep_52_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34463_2_lut (.I0(n1752), .I1(n1653_adj_5178), .I2(GND_net), 
            .I3(GND_net), .O(n49900));
    defparam i34463_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_31__I_0_i1178_rep_51_3_lut (.I0(n48697), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n48696));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1178_rep_51_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34963_4_lut (.I0(n48696), .I1(n1628), .I2(n1851), .I3(n49900), 
            .O(n50401));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34963_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i16118_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5138), 
            .I3(n27976), .O(n29645));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16118_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34964_3_lut (.I0(n50401), .I1(n1992), .I2(n1950), .I3(GND_net), 
            .O(n2024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i34964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16119_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5138), 
            .I3(n27971), .O(n29646));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16119_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16120_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_5094), 
            .I3(n27976), .O(n29647));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16120_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16121_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_5094), 
            .I3(n27971), .O(n29648));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16121_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i16122_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n35414), 
            .I3(n27976), .O(n29649));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16122_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16123_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n35414), 
            .I3(n27971), .O(n29650));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16123_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16125_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n29176), 
            .I3(GND_net), .O(n29652));   // verilog/coms.v(127[12] 300[6])
    defparam i16125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16126_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n29176), 
            .I3(GND_net), .O(n29653));   // verilog/coms.v(127[12] 300[6])
    defparam i16126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16127_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n45660), .I3(GND_net), .O(n29654));   // verilog/coms.v(127[12] 300[6])
    defparam i16127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16128_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n46973), .I3(GND_net), 
            .O(n29655));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16130_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n29176), .I3(GND_net), .O(n29657));   // verilog/coms.v(127[12] 300[6])
    defparam i16130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16131_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n29176), .I3(GND_net), .O(n29658));   // verilog/coms.v(127[12] 300[6])
    defparam i16131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29565_2_lut (.I0(n82), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n44919));
    defparam i29565_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i22707_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n36227));
    defparam i22707_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i3_4_lut_adj_1801 (.I0(n5_adj_5187), .I1(n44919), .I2(\FRAME_MATCHER.i_31__N_2624 ), 
            .I3(n3303), .O(n46694));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1801.LUT_INIT = 16'hbbfb;
    SB_LUT4 i1_4_lut_adj_1802 (.I0(\FRAME_MATCHER.i_31__N_2622 ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n46694), .I3(n25063), .O(n43483));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1802.LUT_INIT = 16'heafa;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(enable_slow_N_4190), .I1(data_ready), 
            .I2(state_adj_5289[1]), .I3(state_adj_5289[0]), .O(n43841));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'hccd0;
    SB_LUT4 i1_4_lut_adj_1804 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n47336));
    defparam i1_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i16134_4_lut (.I0(rw), .I1(state_adj_5289[0]), .I2(state_adj_5289[1]), 
            .I3(n5741), .O(n29661));   // verilog/eeprom.v(26[8] 58[4])
    defparam i16134_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i16135_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5298[1]), .I2(n20400), 
            .I3(n4_adj_5101), .O(n29662));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i16135_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i16136_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4087[0]), 
            .I3(enable_slow_N_4190), .O(n29663));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16136_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i16137_4_lut (.I0(state_7__N_4103[3]), .I1(data[0]), .I2(n10_adj_5222), 
            .I3(n27984), .O(n29664));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16137_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n1329), .I1(n36227), .I2(n1330), .I3(n1331), 
            .O(n45164));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'ha080;
    SB_LUT4 i35370_4_lut (.I0(n45164), .I1(n1323), .I2(n1324), .I3(n47336), 
            .O(n1356));
    defparam i35370_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut_4_lut (.I0(n2), .I1(encoder0_position[31]), 
            .I2(n47474), .I3(n7350), .O(n828));
    defparam encoder0_position_31__I_0_i500_4_lut_4_lut.LUT_INIT = 16'ha808;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653_adj_5178), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5098));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35384_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50822));
    defparam i35384_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35367_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50805));
    defparam i35367_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35351_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50789));
    defparam i35351_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35336_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50774));
    defparam i35336_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35322_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50760));
    defparam i35322_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22703_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n36223));
    defparam i22703_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5188));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1806 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n47410));
    defparam i1_2_lut_adj_1806.LUT_INIT = 16'heeee;
    SB_LUT4 i16405_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n46973), .I3(GND_net), 
            .O(n29932));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(n1429), .I1(n36223), .I2(n1430), .I3(n1431), 
            .O(n45183));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'ha080;
    SB_LUT4 i16406_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n46973), .I3(GND_net), 
            .O(n29933));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16407_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n46973), .I3(GND_net), 
            .O(n29934));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16408_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n46973), .I3(GND_net), 
            .O(n29935));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16409_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n46973), .I3(GND_net), 
            .O(n29936));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n47410), 
            .O(n47416));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 i35387_4_lut (.I0(n1423), .I1(n1422), .I2(n47416), .I3(n45183), 
            .O(n1455));
    defparam i35387_4_lut.LUT_INIT = 16'h0001;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 i16410_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n46973), .I3(GND_net), 
            .O(n29937));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1809 (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(\ID_READOUT_FSM.state [0]), .I3(GND_net), .O(n46973));
    defparam i2_3_lut_adj_1809.LUT_INIT = 16'hdfdf;
    SB_LUT4 i16411_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n46973), .I3(GND_net), 
            .O(n29938));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i16411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16412_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n45660), .I3(GND_net), .O(n29939));   // verilog/coms.v(127[12] 300[6])
    defparam i16412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_5092), .I3(control_mode[2]), .O(n27828));   // verilog/TinyFPGA_B.v(268[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16165_3_lut (.I0(h1), .I1(reg_B[2]), .I2(n46952), .I3(GND_net), 
            .O(n29692));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i16165_3_lut.LUT_INIT = 16'hacac;
    motorControl control (.\Kp[10] (Kp[10]), .GND_net(GND_net), .IntegralLimit({IntegralLimit}), 
            .\Kp[11] (Kp[11]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[12] (Kp[12]), 
            .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .\Kp[15] (Kp[15]), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Kp[4] (Kp[4]), 
            .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Ki[2] (Ki[2]), 
            .\Kp[8] (Kp[8]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Kp[9] (Kp[9]), 
            .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), 
            .\Ki[13] (Ki[13]), .PWMLimit({PWMLimit}), .duty({duty}), .clk32MHz(clk32MHz), 
            .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .VCC_net(VCC_net), .setpoint({setpoint}), 
            .motor_state({motor_state})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(271[16] 283[4])
    SB_LUT4 i16166_3_lut (.I0(h2), .I1(reg_B[1]), .I2(n46952), .I3(GND_net), 
            .O(n29693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i16166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16167_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n43061), .I3(GND_net), .O(n29694));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16413_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n45660), .I3(GND_net), .O(n29940));   // verilog/coms.v(127[12] 300[6])
    defparam i16413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16414_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n45660), .I3(GND_net), .O(n29941));   // verilog/coms.v(127[12] 300[6])
    defparam i16414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16168_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n43061), .I3(GND_net), .O(n29695));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16169_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n43061), .I3(GND_net), .O(n29696));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16170_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n43061), .I3(GND_net), .O(n29697));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16171_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n43061), .I3(GND_net), .O(n29698));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16415_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n45660), .I3(GND_net), .O(n29942));   // verilog/coms.v(127[12] 300[6])
    defparam i16415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16172_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n43061), .I3(GND_net), .O(n29699));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16416_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n45660), .I3(GND_net), .O(n29943));   // verilog/coms.v(127[12] 300[6])
    defparam i16416_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16417_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n45660), .I3(GND_net), .O(n29944));   // verilog/coms.v(127[12] 300[6])
    defparam i16417_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16173_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n43061), .I3(GND_net), .O(n29700));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16174_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n43061), .I3(GND_net), .O(n29701));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16418_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n45660), .I3(GND_net), .O(n29945));   // verilog/coms.v(127[12] 300[6])
    defparam i16418_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16175_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n43061), .I3(GND_net), .O(n29702));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16419_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n45660), .I3(GND_net), .O(n29946));   // verilog/coms.v(127[12] 300[6])
    defparam i16419_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16420_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n45660), .I3(GND_net), .O(n29947));   // verilog/coms.v(127[12] 300[6])
    defparam i16420_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16421_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n45660), .I3(GND_net), .O(n29948));   // verilog/coms.v(127[12] 300[6])
    defparam i16421_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16422_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n45660), .I3(GND_net), .O(n29949));   // verilog/coms.v(127[12] 300[6])
    defparam i16422_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16423_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n45660), .I3(GND_net), .O(n29950));   // verilog/coms.v(127[12] 300[6])
    defparam i16423_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16424_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n45660), .I3(GND_net), .O(n29951));   // verilog/coms.v(127[12] 300[6])
    defparam i16424_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16425_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n45660), .I3(GND_net), .O(n29952));   // verilog/coms.v(127[12] 300[6])
    defparam i16425_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16176_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n43061), .I3(GND_net), .O(n29703));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34727_3_lut (.I0(n2049), .I1(n1950), .I2(n1851), .I3(GND_net), 
            .O(n50164));
    defparam i34727_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 i21773_1_lut_2_lut (.I0(n25336), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n1910));
    defparam i21773_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i16162_3_lut_4_lut (.I0(n1617), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_3907), .O(n29689));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16162_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5298[1]), .I1(r_SM_Main_adj_5298[0]), 
            .I2(r_SM_Main_2__N_3613[1]), .I3(r_SM_Main_adj_5298[2]), .O(n51668));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i34420_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n49662));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34420_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i29555_4_lut_4_lut_4_lut (.I0(h1), .I1(h3), .I2(h2), .I3(commutation_state[2]), 
            .O(n44909));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i29555_4_lut_4_lut_4_lut.LUT_INIT = 16'hc544;
    SB_LUT4 i34377_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n49676));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34377_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i6649_3_lut_4_lut_4_lut (.I0(commutation_state[1]), .I1(commutation_state[2]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_367));
    defparam i6649_3_lut_4_lut_4_lut.LUT_INIT = 16'h1a14;
    SB_LUT4 i6651_3_lut_4_lut_4_lut (.I0(commutation_state[1]), .I1(commutation_state[2]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_384));
    defparam i6651_3_lut_4_lut_4_lut.LUT_INIT = 16'ha141;
    SB_LUT4 i16426_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n45660), .I3(GND_net), .O(n29953));   // verilog/coms.v(127[12] 300[6])
    defparam i16426_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16427_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n45660), .I3(GND_net), .O(n29954));   // verilog/coms.v(127[12] 300[6])
    defparam i16427_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16428_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n45660), .I3(GND_net), .O(n29955));   // verilog/coms.v(127[12] 300[6])
    defparam i16428_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16429_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n45660), .I3(GND_net), .O(n29956));   // verilog/coms.v(127[12] 300[6])
    defparam i16429_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34430_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n49677));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34430_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i16430_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n45660), .I3(GND_net), .O(n29957));   // verilog/coms.v(127[12] 300[6])
    defparam i16430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16431_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n45660), .I3(GND_net), .O(n29958));   // verilog/coms.v(127[12] 300[6])
    defparam i16431_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16432_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n45660), .I3(GND_net), .O(n29959));   // verilog/coms.v(127[12] 300[6])
    defparam i16432_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34429_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n49678));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34429_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i16433_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n45660), .I3(GND_net), .O(n29960));   // verilog/coms.v(127[12] 300[6])
    defparam i16433_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34428_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n49679));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34428_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i21772_2_lut (.I0(n25336), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n35282));
    defparam i21772_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_238_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16434_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n45660), .I3(GND_net), .O(n29961));   // verilog/coms.v(127[12] 300[6])
    defparam i16434_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16435_3_lut (.I0(\data_out_frame[27] [1]), .I1(n41916), .I2(n29310), 
            .I3(GND_net), .O(n29962));   // verilog/coms.v(127[12] 300[6])
    defparam i16435_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i16436_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n25135), .I3(GND_net), .O(n29963));   // verilog/coms.v(127[12] 300[6])
    defparam i16436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16437_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n25135), .I3(GND_net), .O(n29964));   // verilog/coms.v(127[12] 300[6])
    defparam i16437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34427_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n49680));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34427_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i16438_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n25135), .I3(GND_net), .O(n29965));   // verilog/coms.v(127[12] 300[6])
    defparam i16438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i34426_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n49681));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34426_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 mux_238_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16439_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n25135), .I3(GND_net), .O(n29966));   // verilog/coms.v(127[12] 300[6])
    defparam i16439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16440_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n25135), .I3(GND_net), .O(n29967));   // verilog/coms.v(127[12] 300[6])
    defparam i16440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34425_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n49682));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i34425_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i29535_3_lut (.I0(n7), .I1(n7355), .I2(n44865), .I3(GND_net), 
            .O(n44886));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i29535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1810 (.I0(commutation_state[0]), .I1(n4_adj_5231), 
            .I2(commutation_state_prev[0]), .I3(dti_N_416), .O(n29117));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_2_lut_4_lut_adj_1810.LUT_INIT = 16'hdeff;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n29208), 
            .I3(rx_data_ready), .O(n43733));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i16441_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n25135), .I3(GND_net), .O(n29968));   // verilog/coms.v(127[12] 300[6])
    defparam i16441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1811 (.I0(n5_adj_5105), .I1(n3), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n47474));
    defparam i1_3_lut_adj_1811.LUT_INIT = 16'h8080;
    SB_LUT4 mux_238_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16442_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n25135), .I3(GND_net), .O(n29969));   // verilog/coms.v(127[12] 300[6])
    defparam i16442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1812 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n47122));
    defparam i1_2_lut_adj_1812.LUT_INIT = 16'heeee;
    SB_LUT4 i16443_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n25135), .I3(GND_net), .O(n29970));   // verilog/coms.v(127[12] 300[6])
    defparam i16443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16444_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n25135), .I3(GND_net), .O(n29971));   // verilog/coms.v(127[12] 300[6])
    defparam i16444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22847_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n36369));
    defparam i22847_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1813 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n47122), 
            .O(n47128));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n1529), .I1(n47128), .I2(n36369), .I3(n1530), 
            .O(n47130));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'heccc;
    SB_LUT4 i16445_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n25135), .I3(GND_net), .O(n29972));   // verilog/coms.v(127[12] 300[6])
    defparam i16445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16446_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n25135), .I3(GND_net), .O(n29973));   // verilog/coms.v(127[12] 300[6])
    defparam i16446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16447_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n25135), .I3(GND_net), .O(n29974));   // verilog/coms.v(127[12] 300[6])
    defparam i16447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16448_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n25135), .I3(GND_net), .O(n29975));   // verilog/coms.v(127[12] 300[6])
    defparam i16448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16449_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n25135), .I3(GND_net), .O(n29976));   // verilog/coms.v(127[12] 300[6])
    defparam i16449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21617_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(84[16:31])
    defparam i21617_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16450_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n25135), .I3(GND_net), .O(n29977));   // verilog/coms.v(127[12] 300[6])
    defparam i16450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16451_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n25135), .I3(GND_net), .O(n29978));   // verilog/coms.v(127[12] 300[6])
    defparam i16451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21616_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(82[16:31])
    defparam i21616_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21999_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(80[16:31])
    defparam i21999_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i16452_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n25135), .I3(GND_net), .O(n29979));   // verilog/coms.v(127[12] 300[6])
    defparam i16452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16106_4_lut_4_lut (.I0(state[1]), .I1(state[0]), .I2(n29323), 
            .I3(state_3__N_528[1]), .O(n29633));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16106_4_lut_4_lut.LUT_INIT = 16'hfa7a;
    SB_LUT4 i16453_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n25135), .I3(GND_net), .O(n29980));   // verilog/coms.v(127[12] 300[6])
    defparam i16453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16454_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n25135), .I3(GND_net), .O(n29981));   // verilog/coms.v(127[12] 300[6])
    defparam i16454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_3_lut (.I0(h2), .I1(h3), .I2(h1), .I3(GND_net), .O(n6_adj_5180));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1815 (.I0(h3), .I1(h2), .I2(h1), .I3(GND_net), 
            .O(commutation_state_7__N_216[0]));   // verilog/TinyFPGA_B.v(148[4] 150[7])
    defparam i1_3_lut_adj_1815.LUT_INIT = 16'h1414;
    SB_LUT4 i16455_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n25135), .I3(GND_net), .O(n29982));   // verilog/coms.v(127[12] 300[6])
    defparam i16455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16456_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n25135), .I3(GND_net), .O(n29983));   // verilog/coms.v(127[12] 300[6])
    defparam i16456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16457_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n25135), .I3(GND_net), .O(n29984));   // verilog/coms.v(127[12] 300[6])
    defparam i16457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16458_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n25135), .I3(GND_net), .O(n29985));   // verilog/coms.v(127[12] 300[6])
    defparam i16458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16459_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n25135), .I3(GND_net), .O(n29986));   // verilog/coms.v(127[12] 300[6])
    defparam i16459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16460_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n25135), .I3(GND_net), .O(n29987));   // verilog/coms.v(127[12] 300[6])
    defparam i16460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16461_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n25135), .I3(GND_net), .O(n29988));   // verilog/coms.v(127[12] 300[6])
    defparam i16461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16462_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n25135), .I3(GND_net), .O(n29989));   // verilog/coms.v(127[12] 300[6])
    defparam i16462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16463_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n25135), .I3(GND_net), .O(n29990));   // verilog/coms.v(127[12] 300[6])
    defparam i16463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i35405_4_lut (.I0(n1522), .I1(n1521), .I2(n47130), .I3(n1523), 
            .O(n1554));
    defparam i35405_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22691_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n36211));
    defparam i22691_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n47428));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(n1629), .I1(n36211), .I2(n1630), .I3(n1631), 
            .O(n45192));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'ha080;
    SB_LUT4 i16464_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n25135), .I3(GND_net), .O(n29991));   // verilog/coms.v(127[12] 300[6])
    defparam i16464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16465_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n25135), .I3(GND_net), .O(n29992));   // verilog/coms.v(127[12] 300[6])
    defparam i16465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16466_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n25135), .I3(GND_net), .O(n29993));   // verilog/coms.v(127[12] 300[6])
    defparam i16466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16467_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n25135), .I3(GND_net), .O(n29994));   // verilog/coms.v(127[12] 300[6])
    defparam i16467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16468_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n25135), .I3(GND_net), .O(n29995));   // verilog/coms.v(127[12] 300[6])
    defparam i16468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16469_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n25135), .I3(GND_net), .O(n29996));   // verilog/coms.v(127[12] 300[6])
    defparam i16469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16470_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n25135), .I3(GND_net), .O(n29997));   // verilog/coms.v(127[12] 300[6])
    defparam i16470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16471_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n25135), .I3(GND_net), .O(n29998));   // verilog/coms.v(127[12] 300[6])
    defparam i16471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16472_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n25135), .I3(GND_net), .O(n29999));   // verilog/coms.v(127[12] 300[6])
    defparam i16472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16473_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n25135), .I3(GND_net), .O(n30000));   // verilog/coms.v(127[12] 300[6])
    defparam i16473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16474_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n25135), .I3(GND_net), .O(n30001));   // verilog/coms.v(127[12] 300[6])
    defparam i16474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16475_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n25135), .I3(GND_net), .O(n30002));   // verilog/coms.v(127[12] 300[6])
    defparam i16475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16476_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n25135), .I3(GND_net), .O(n30003));   // verilog/coms.v(127[12] 300[6])
    defparam i16476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16477_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n25135), .I3(GND_net), .O(n30004));   // verilog/coms.v(127[12] 300[6])
    defparam i16477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15927_2_lut (.I0(n29125), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n29460));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i15927_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35174_4_lut (.I0(commutation_state[1]), .I1(n25336), .I2(dti), 
            .I3(commutation_state[2]), .O(n29125));
    defparam i35174_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n1623), .I1(n45192), .I2(n1624), .I3(n47428), 
            .O(n47434));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093_adj_5168), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1819 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5092));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i4_4_lut_adj_1819.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1820 (.I0(control_mode[6]), .I1(n10_adj_5092), 
            .I2(control_mode[2]), .I3(GND_net), .O(n27996));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i5_3_lut_adj_1820.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1821 (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n44138));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut_adj_1821.LUT_INIT = 16'h4000;
    SB_LUT4 i1_2_lut_adj_1822 (.I0(n27828), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5132));   // verilog/TinyFPGA_B.v(268[5:22])
    defparam i1_2_lut_adj_1822.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut_adj_1823 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n27996), .I3(GND_net), .O(n15_adj_5134));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i2_3_lut_adj_1823.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_238_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5134), .I3(n15_adj_5132), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i16177_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n43061), .I3(GND_net), .O(n29704));   // verilog/neopixel.v(35[12] 117[6])
    defparam i16177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i24_1_lut (.I0(duty[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16478_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n25135), .I3(GND_net), .O(n30005));   // verilog/coms.v(127[12] 300[6])
    defparam i16478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16479_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n25135), .I3(GND_net), .O(n30006));   // verilog/coms.v(127[12] 300[6])
    defparam i16479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16480_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n25135), .I3(GND_net), .O(n30007));   // verilog/coms.v(127[12] 300[6])
    defparam i16480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16481_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n25135), .I3(GND_net), .O(n30008));   // verilog/coms.v(127[12] 300[6])
    defparam i16481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16482_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n25135), .I3(GND_net), .O(n30009));   // verilog/coms.v(127[12] 300[6])
    defparam i16482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16484_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n25135), .I3(GND_net), .O(n30011));   // verilog/coms.v(127[12] 300[6])
    defparam i16484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1246_rep_37_3_lut (.I0(n1894), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n48682));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1246_rep_37_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16485_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n25135), 
            .I3(GND_net), .O(n30012));   // verilog/coms.v(127[12] 300[6])
    defparam i16485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35429_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n47434), 
            .O(n1653_adj_5178));
    defparam i35429_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i16486_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n25135), 
            .I3(GND_net), .O(n30013));   // verilog/coms.v(127[12] 300[6])
    defparam i16486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16487_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n25135), 
            .I3(GND_net), .O(n30014));   // verilog/coms.v(127[12] 300[6])
    defparam i16487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16488_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n25135), 
            .I3(GND_net), .O(n30015));   // verilog/coms.v(127[12] 300[6])
    defparam i16488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16489_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n25135), 
            .I3(GND_net), .O(n30016));   // verilog/coms.v(127[12] 300[6])
    defparam i16489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16490_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n25135), 
            .I3(GND_net), .O(n30017));   // verilog/coms.v(127[12] 300[6])
    defparam i16490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16491_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n25135), 
            .I3(GND_net), .O(n30018));   // verilog/coms.v(127[12] 300[6])
    defparam i16491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16492_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n25135), 
            .I3(GND_net), .O(n30019));   // verilog/coms.v(127[12] 300[6])
    defparam i16492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16493_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n25135), 
            .I3(GND_net), .O(n30020));   // verilog/coms.v(127[12] 300[6])
    defparam i16493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16494_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n25135), 
            .I3(GND_net), .O(n30021));   // verilog/coms.v(127[12] 300[6])
    defparam i16494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16495_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n25135), 
            .I3(GND_net), .O(n30022));   // verilog/coms.v(127[12] 300[6])
    defparam i16495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16496_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n25135), 
            .I3(GND_net), .O(n30023));   // verilog/coms.v(127[12] 300[6])
    defparam i16496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16497_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n25135), 
            .I3(GND_net), .O(n30024));   // verilog/coms.v(127[12] 300[6])
    defparam i16497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16498_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n25135), 
            .I3(GND_net), .O(n30025));   // verilog/coms.v(127[12] 300[6])
    defparam i16498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16499_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n25135), 
            .I3(GND_net), .O(n30026));   // verilog/coms.v(127[12] 300[6])
    defparam i16499_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16500_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n25135), 
            .I3(GND_net), .O(n30027));   // verilog/coms.v(127[12] 300[6])
    defparam i16500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16501_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n25135), 
            .I3(GND_net), .O(n30028));   // verilog/coms.v(127[12] 300[6])
    defparam i16501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16502_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n25135), 
            .I3(GND_net), .O(n30029));   // verilog/coms.v(127[12] 300[6])
    defparam i16502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16503_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n25135), 
            .I3(GND_net), .O(n30030));   // verilog/coms.v(127[12] 300[6])
    defparam i16503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16504_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n25135), 
            .I3(GND_net), .O(n30031));   // verilog/coms.v(127[12] 300[6])
    defparam i16504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16505_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n25135), 
            .I3(GND_net), .O(n30032));   // verilog/coms.v(127[12] 300[6])
    defparam i16505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16506_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n25135), 
            .I3(GND_net), .O(n30033));   // verilog/coms.v(127[12] 300[6])
    defparam i16506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16507_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n25135), 
            .I3(GND_net), .O(n30034));   // verilog/coms.v(127[12] 300[6])
    defparam i16507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16508_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n25135), 
            .I3(GND_net), .O(n30035));   // verilog/coms.v(127[12] 300[6])
    defparam i16508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16509_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n25135), .I3(GND_net), .O(n30036));   // verilog/coms.v(127[12] 300[6])
    defparam i16509_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16510_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n25135), .I3(GND_net), .O(n30037));   // verilog/coms.v(127[12] 300[6])
    defparam i16510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16511_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n25135), .I3(GND_net), .O(n30038));   // verilog/coms.v(127[12] 300[6])
    defparam i16511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16512_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n25135), .I3(GND_net), .O(n30039));   // verilog/coms.v(127[12] 300[6])
    defparam i16512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16513_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n25135), .I3(GND_net), .O(n30040));   // verilog/coms.v(127[12] 300[6])
    defparam i16513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16514_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n25135), .I3(GND_net), .O(n30041));   // verilog/coms.v(127[12] 300[6])
    defparam i16514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16515_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n25135), .I3(GND_net), .O(n30042));   // verilog/coms.v(127[12] 300[6])
    defparam i16515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16516_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n25135), .I3(GND_net), .O(n30043));   // verilog/coms.v(127[12] 300[6])
    defparam i16516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16517_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n25135), .I3(GND_net), .O(n30044));   // verilog/coms.v(127[12] 300[6])
    defparam i16517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16518_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n25135), .I3(GND_net), .O(n30045));   // verilog/coms.v(127[12] 300[6])
    defparam i16518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16519_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n25135), .I3(GND_net), .O(n30046));   // verilog/coms.v(127[12] 300[6])
    defparam i16519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16520_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n25135), .I3(GND_net), .O(n30047));   // verilog/coms.v(127[12] 300[6])
    defparam i16520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_5157), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n936));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16521_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n25135), .I3(GND_net), .O(n30048));   // verilog/coms.v(127[12] 300[6])
    defparam i16521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16522_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n25135), .I3(GND_net), .O(n30049));   // verilog/coms.v(127[12] 300[6])
    defparam i16522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16523_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n25135), .I3(GND_net), .O(n30050));   // verilog/coms.v(127[12] 300[6])
    defparam i16523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16524_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n25135), .I3(GND_net), .O(n30051));   // verilog/coms.v(127[12] 300[6])
    defparam i16524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16525_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n25135), .I3(GND_net), .O(n30052));   // verilog/coms.v(127[12] 300[6])
    defparam i16525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16526_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n25135), .I3(GND_net), .O(n30053));   // verilog/coms.v(127[12] 300[6])
    defparam i16526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16527_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n25135), .I3(GND_net), .O(n30054));   // verilog/coms.v(127[12] 300[6])
    defparam i16527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16528_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n25135), .I3(GND_net), .O(n30055));   // verilog/coms.v(127[12] 300[6])
    defparam i16528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16529_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n25135), .I3(GND_net), .O(n30056));   // verilog/coms.v(127[12] 300[6])
    defparam i16529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16530_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n25135), .I3(GND_net), .O(n30057));   // verilog/coms.v(127[12] 300[6])
    defparam i16530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16531_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n25135), .I3(GND_net), .O(n30058));   // verilog/coms.v(127[12] 300[6])
    defparam i16531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16532_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n25135), .I3(GND_net), .O(n30059));   // verilog/coms.v(127[12] 300[6])
    defparam i16532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16533_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n25135), .I3(GND_net), .O(n30060));   // verilog/coms.v(127[12] 300[6])
    defparam i16533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16534_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n25135), .I3(GND_net), .O(n30061));   // verilog/coms.v(127[12] 300[6])
    defparam i16534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16535_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n25135), .I3(GND_net), .O(n30062));   // verilog/coms.v(127[12] 300[6])
    defparam i16535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16536_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n25135), .I3(GND_net), .O(n30063));   // verilog/coms.v(127[12] 300[6])
    defparam i16536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16537_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n25135), .I3(GND_net), .O(n30064));   // verilog/coms.v(127[12] 300[6])
    defparam i16537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16538_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n25135), .I3(GND_net), .O(n30065));   // verilog/coms.v(127[12] 300[6])
    defparam i16538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16539_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n25135), .I3(GND_net), .O(n30066));   // verilog/coms.v(127[12] 300[6])
    defparam i16539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16540_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n25135), .I3(GND_net), .O(n30067));   // verilog/coms.v(127[12] 300[6])
    defparam i16540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16541_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n25135), .I3(GND_net), .O(n30068));   // verilog/coms.v(127[12] 300[6])
    defparam i16541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16542_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n25135), .I3(GND_net), .O(n30069));   // verilog/coms.v(127[12] 300[6])
    defparam i16542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16543_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n25135), .I3(GND_net), .O(n30070));   // verilog/coms.v(127[12] 300[6])
    defparam i16543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16544_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n25135), .I3(GND_net), .O(n30071));   // verilog/coms.v(127[12] 300[6])
    defparam i16544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16545_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n25135), .I3(GND_net), .O(n30072));   // verilog/coms.v(127[12] 300[6])
    defparam i16545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16546_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n25135), .I3(GND_net), .O(n30073));   // verilog/coms.v(127[12] 300[6])
    defparam i16546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16547_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n25135), .I3(GND_net), .O(n30074));   // verilog/coms.v(127[12] 300[6])
    defparam i16547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16548_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n25135), .I3(GND_net), .O(n30075));   // verilog/coms.v(127[12] 300[6])
    defparam i16548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16549_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n25135), .I3(GND_net), .O(n30076));   // verilog/coms.v(127[12] 300[6])
    defparam i16549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16550_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n25135), .I3(GND_net), .O(n30077));   // verilog/coms.v(127[12] 300[6])
    defparam i16550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16551_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n25135), .I3(GND_net), .O(n30078));   // verilog/coms.v(127[12] 300[6])
    defparam i16551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16552_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n25135), .I3(GND_net), .O(n30079));   // verilog/coms.v(127[12] 300[6])
    defparam i16552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n29208));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h4303;
    SB_LUT4 i1_3_lut_adj_1824 (.I0(n1726), .I1(n1728), .I2(n1727), .I3(GND_net), 
            .O(n47056));
    defparam i1_3_lut_adj_1824.LUT_INIT = 16'hfefe;
    SB_LUT4 i22843_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n36365));
    defparam i22843_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i16147_3_lut_4_lut (.I0(n1658), .I1(b_prev_adj_5136), .I2(a_new_adj_5265[1]), 
            .I3(direction_N_3907_adj_5137), .O(n29674));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16147_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_4_lut_adj_1825 (.I0(n1723), .I1(n1724), .I2(n47056), .I3(n1725), 
            .O(n47062));
    defparam i1_4_lut_adj_1825.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1826 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n47440));
    defparam i1_2_lut_adj_1826.LUT_INIT = 16'h8888;
    coms neopxl_color_23__I_0 (.\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .CLK_c(CLK_c), .GND_net(GND_net), 
         .n29756(n29756), .control_mode({control_mode}), .n25135(n25135), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n29755(n29755), 
         .\FRAME_MATCHER.i_31__N_2622 (\FRAME_MATCHER.i_31__N_2622 ), .n29754(n29754), 
         .\FRAME_MATCHER.state_31__N_2660[2] (\FRAME_MATCHER.state_31__N_2660 [2]), 
         .\FRAME_MATCHER.i_31__N_2626 (\FRAME_MATCHER.i_31__N_2626 ), .n4452(n4452), 
         .n7(n7_adj_5185), .rx_data({rx_data}), .n771(n771), .n29753(n29753), 
         .n29752(n29752), .n45880(n45880), .n3303(n3303), .\data_in[2] ({\data_in[2] }), 
         .\data_in[0] ({\data_in[0] }), .\data_in[3] ({\data_in[3] }), .\data_in[1] ({\data_in[1] }), 
         .n63(n63), .\data_out_frame[8] ({\data_out_frame[8] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .n29751(n29751), .n29750(n29750), .n29749(n29749), .PWMLimit({PWMLimit}), 
         .n29748(n29748), .\data_in_frame[8] ({\data_in_frame[8] }), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n29747(n29747), .rx_data_ready(rx_data_ready), .setpoint({setpoint}), 
         .n29746(n29746), .\data_in_frame[10] ({\data_in_frame[10] }), .n29745(n29745), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .n29744(n29744), .n29743(n29743), .n29742(n29742), .n29741(n29741), 
         .n29740(n29740), .n29739(n29739), .n29738(n29738), .n29737(n29737), 
         .n29736(n29736), .n29735(n29735), .n29734(n29734), .n29733(n29733), 
         .n29732(n29732), .n29731(n29731), .n29730(n29730), .n29729(n29729), 
         .n29728(n29728), .n29727(n29727), .n51593(n51593), .n51594(n51594), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .n14(n14_adj_5229), 
         .tx_active(tx_active), .DE_c(DE_c), .LED_c(LED_c), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .n25063(n25063), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[6] ({\data_in_frame[6] }), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .n29310(n29310), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .\data_out_frame[27][1] (\data_out_frame[27] [1]), 
         .ID({ID}), .n4(n4_adj_5093), .n29176(n29176), .n41916(n41916), 
         .n30209(n30209), .IntegralLimit({IntegralLimit}), .n30208(n30208), 
         .n30207(n30207), .n30206(n30206), .n30205(n30205), .n30204(n30204), 
         .n30203(n30203), .n30202(n30202), .n30201(n30201), .n30200(n30200), 
         .n30199(n30199), .n30198(n30198), .n30197(n30197), .n30196(n30196), 
         .n30195(n30195), .n30194(n30194), .n30193(n30193), .n30192(n30192), 
         .n30191(n30191), .n30190(n30190), .n30189(n30189), .n30188(n30188), 
         .n30186(n30186), .n30185(n30185), .n30184(n30184), .n30183(n30183), 
         .n30182(n30182), .n30181(n30181), .n30180(n30180), .n30179(n30179), 
         .n30178(n30178), .n30177(n30177), .n30176(n30176), .n30175(n30175), 
         .n30174(n30174), .n30173(n30173), .n30172(n30172), .n30171(n30171), 
         .n30170(n30170), .n30169(n30169), .n30168(n30168), .n30167(n30167), 
         .n30166(n30166), .n30165(n30165), .n30164(n30164), .n30163(n30163), 
         .n30162(n30162), .n30161(n30161), .n30160(n30160), .n30159(n30159), 
         .n30158(n30158), .n30157(n30157), .n30156(n30156), .n30155(n30155), 
         .n30154(n30154), .\Kp[1] (Kp[1]), .n30153(n30153), .\Kp[2] (Kp[2]), 
         .n30152(n30152), .\Kp[3] (Kp[3]), .n30151(n30151), .\Kp[4] (Kp[4]), 
         .n30150(n30150), .\Kp[5] (Kp[5]), .n30149(n30149), .\Kp[6] (Kp[6]), 
         .n30148(n30148), .\Kp[7] (Kp[7]), .n30147(n30147), .\Kp[8] (Kp[8]), 
         .n30146(n30146), .\Kp[9] (Kp[9]), .n30145(n30145), .\Kp[10] (Kp[10]), 
         .n30144(n30144), .\Kp[11] (Kp[11]), .n30143(n30143), .\Kp[12] (Kp[12]), 
         .n30141(n30141), .\Kp[13] (Kp[13]), .n30140(n30140), .\Kp[14] (Kp[14]), 
         .n30139(n30139), .\Kp[15] (Kp[15]), .n30138(n30138), .\Ki[1] (Ki[1]), 
         .n30137(n30137), .\Ki[2] (Ki[2]), .n30136(n30136), .\Ki[3] (Ki[3]), 
         .n30135(n30135), .\Ki[4] (Ki[4]), .n30134(n30134), .\Ki[5] (Ki[5]), 
         .n30133(n30133), .\Ki[6] (Ki[6]), .n30132(n30132), .\Ki[7] (Ki[7]), 
         .n30131(n30131), .\Ki[8] (Ki[8]), .n30130(n30130), .\Ki[9] (Ki[9]), 
         .n30129(n30129), .\Ki[10] (Ki[10]), .n30128(n30128), .\Ki[11] (Ki[11]), 
         .n30127(n30127), .\Ki[12] (Ki[12]), .n30126(n30126), .\Ki[13] (Ki[13]), 
         .n30125(n30125), .\Ki[14] (Ki[14]), .n30124(n30124), .\Ki[15] (Ki[15]), 
         .n30123(n30123), .n30122(n30122), .n30121(n30121), .n30120(n30120), 
         .n30119(n30119), .n30118(n30118), .n30117(n30117), .n30116(n30116), 
         .n30115(n30115), .n30114(n30114), .n30113(n30113), .n30112(n30112), 
         .n30111(n30111), .n30110(n30110), .n30109(n30109), .n30108(n30108), 
         .n30107(n30107), .n30106(n30106), .n30105(n30105), .n30104(n30104), 
         .n30103(n30103), .n30102(n30102), .n30101(n30101), .n30100(n30100), 
         .n30099(n30099), .n30098(n30098), .n30097(n30097), .n30096(n30096), 
         .n30095(n30095), .n30094(n30094), .n30093(n30093), .n30092(n30092), 
         .n30091(n30091), .n30090(n30090), .n30089(n30089), .n30088(n30088), 
         .n30087(n30087), .n30086(n30086), .n30085(n30085), .n30084(n30084), 
         .n30083(n30083), .n30082(n30082), .n30081(n30081), .n30080(n30080), 
         .n30079(n30079), .n30078(n30078), .n30077(n30077), .n30076(n30076), 
         .n30075(n30075), .n30074(n30074), .n30073(n30073), .n30072(n30072), 
         .n30071(n30071), .n30070(n30070), .n30069(n30069), .n30068(n30068), 
         .n30067(n30067), .n30066(n30066), .n30065(n30065), .n30064(n30064), 
         .n30063(n30063), .n30062(n30062), .n30061(n30061), .n30060(n30060), 
         .n30059(n30059), .n30058(n30058), .n30057(n30057), .n30056(n30056), 
         .n30055(n30055), .n30054(n30054), .n30053(n30053), .n30052(n30052), 
         .n30051(n30051), .n30050(n30050), .n30049(n30049), .n30048(n30048), 
         .n30047(n30047), .n30046(n30046), .n30045(n30045), .n30044(n30044), 
         .n30043(n30043), .n30042(n30042), .n30041(n30041), .n30040(n30040), 
         .n30039(n30039), .n30038(n30038), .n30037(n30037), .n30036(n30036), 
         .n30035(n30035), .n30034(n30034), .n30033(n30033), .n30032(n30032), 
         .n30031(n30031), .n30030(n30030), .n30029(n30029), .n30028(n30028), 
         .n30027(n30027), .n30026(n30026), .n30025(n30025), .n30024(n30024), 
         .n30023(n30023), .n30022(n30022), .n30021(n30021), .n30020(n30020), 
         .n30019(n30019), .n30018(n30018), .n30017(n30017), .n30016(n30016), 
         .n30015(n30015), .n30014(n30014), .n30013(n30013), .n30012(n30012), 
         .n30011(n30011), .n30009(n30009), .n30008(n30008), .n30007(n30007), 
         .n30006(n30006), .n30005(n30005), .n30004(n30004), .n30003(n30003), 
         .n30002(n30002), .n30001(n30001), .n30000(n30000), .n29999(n29999), 
         .n29998(n29998), .n29997(n29997), .n29996(n29996), .n29995(n29995), 
         .n29994(n29994), .n29993(n29993), .n29992(n29992), .n29991(n29991), 
         .n29990(n29990), .n29989(n29989), .n29988(n29988), .n29987(n29987), 
         .n29986(n29986), .n29985(n29985), .n29984(n29984), .n29983(n29983), 
         .n29982(n29982), .n29981(n29981), .n29980(n29980), .n29979(n29979), 
         .n29978(n29978), .n29977(n29977), .n29976(n29976), .n29975(n29975), 
         .n29974(n29974), .n29973(n29973), .n29972(n29972), .n29971(n29971), 
         .n29970(n29970), .n29969(n29969), .n29968(n29968), .n29967(n29967), 
         .n29966(n29966), .n29965(n29965), .n29964(n29964), .n29963(n29963), 
         .n29962(n29962), .n29961(n29961), .neopxl_color({neopxl_color}), 
         .n29960(n29960), .n29959(n29959), .n29958(n29958), .n29957(n29957), 
         .n29956(n29956), .n29955(n29955), .n29954(n29954), .n29953(n29953), 
         .n29952(n29952), .n29951(n29951), .n29950(n29950), .n29949(n29949), 
         .n29948(n29948), .n29947(n29947), .n29946(n29946), .n29945(n29945), 
         .n29944(n29944), .n29943(n29943), .n29942(n29942), .n29941(n29941), 
         .n29940(n29940), .n29939(n29939), .n43483(n43483), .n29658(n29658), 
         .n29657(n29657), .n29654(n29654), .n29653(n29653), .\Ki[0] (Ki[0]), 
         .n29652(n29652), .\Kp[0] (Kp[0]), .n29626(n29626), .n29625(n29625), 
         .n82(n82), .\FRAME_MATCHER.i_31__N_2624 (\FRAME_MATCHER.i_31__N_2624 ), 
         .n45660(n45660), .\state[0] (state_adj_5307[0]), .\state[2] (state_adj_5307[2]), 
         .\state[3] (state_adj_5307[3]), .n6935(n6935), .n123(n123), .n1(n1), 
         .n29234(n29234), .\r_SM_Main_2__N_3613[1] (r_SM_Main_2__N_3613[1]), 
         .r_SM_Main({r_SM_Main_adj_5298}), .\r_Bit_Index[0] (r_Bit_Index_adj_5300[0]), 
         .tx_o(tx_o), .n44068(n44068), .n29667(n29667), .n29662(n29662), 
         .n51668(n51668), .VCC_net(VCC_net), .n20400(n20400), .n4_adj_6(n4_adj_5101), 
         .tx_enable(tx_enable), .n29246(n29246), .r_Rx_Data(r_Rx_Data), 
         .r_SM_Main_adj_14({r_SM_Main}), .RX_N_10(RX_N_10), .\r_Bit_Index[0]_adj_10 (r_Bit_Index[0]), 
         .n44059(n44059), .\r_SM_Main_2__N_3542[2] (r_SM_Main_2__N_3542[2]), 
         .n27976(n27976), .n4_adj_11(n4_adj_5152), .n29679(n29679), .n29672(n29672), 
         .n43733(n43733), .n29650(n29650), .n29649(n29649), .n29648(n29648), 
         .n29647(n29647), .n29646(n29646), .n29645(n29645), .n29644(n29644), 
         .n44138(n44138), .n4_adj_12(n4_adj_5138), .n4_adj_13(n4_adj_5094), 
         .n27971(n27971), .n35414(n35414)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(238[8] 261[4])
    SB_LUT4 encoder0_position_31__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n47440), .I1(n1722), .I2(n47062), .I3(n36365), 
            .O(n47066));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'hfefc;
    EEPROM eeprom (.GND_net(GND_net), .enable_slow_N_4190(enable_slow_N_4190), 
           .\state[1] (state_adj_5289[1]), .CLK_c(CLK_c), .\state[0] (state_adj_5289[0]), 
           .\state[3] (state_adj_5307[3]), .\state[0]_adj_2 (state_adj_5307[0]), 
           .read(read), .n5740({n5741}), .\state[2] (state_adj_5307[2]), 
           .n29661(n29661), .rw(rw), .n43841(n43841), .data_ready(data_ready), 
           .n6387(n6387), .sda_enable(sda_enable), .\state_7__N_4087[0] (state_7__N_4087[0]), 
           .\saved_addr[0] (saved_addr[0]), .\state_7__N_4103[3] (state_7__N_4103[3]), 
           .n6935(n6935), .scl_enable(scl_enable), .n10(n10_adj_5222), 
           .n35178(n35178), .n35422(n35422), .n8(n8_adj_5158), .VCC_net(VCC_net), 
           .n29675(n29675), .data({data}), .n4(n4_adj_5133), .n4_adj_3(n4), 
           .scl(scl), .sda_out(sda_out), .n30212(n30212), .n29664(n29664), 
           .n29663(n29663), .n29631(n29631), .n29630(n29630), .n29629(n29629), 
           .n29628(n29628), .n29627(n29627), .n49702(n49702), .n27984(n27984), 
           .n28004(n28004)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(387[10] 398[6])
    \quadrature_decoder(1,500000)  quad_counter1 (.\a_new[1] (a_new_adj_5265[1]), 
            .b_prev(b_prev_adj_5136), .GND_net(GND_net), .ENCODER1_B_N_keep(ENCODER1_B_N), 
            .n1653(CLK_c), .ENCODER1_A_N_keep(ENCODER1_A_N), .direction_N_3907(direction_N_3907_adj_5137), 
            .encoder1_position({encoder1_position}), .n29674(n29674), .n1658(n1658), 
            .VCC_net(VCC_net)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(294[57] 301[6])
    \grp_debouncer(3,1000)  debounce (.reg_B({reg_B}), .CLK_c(CLK_c), .n29693(n29693), 
            .data_o({h1, h2, h3}), .n29692(n29692), .data_i({hall1, 
            hall2, hall3}), .n46952(n46952), .n29624(n29624), .GND_net(GND_net), 
            .VCC_net(VCC_net));   // verilog/TinyFPGA_B.v(98[26] 102[3])
    pwm PWM (.GND_net(GND_net), .pwm_out(pwm_out), .clk32MHz(clk32MHz), 
        .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (GND_net, CLK_c, VCC_net, \state[0] , 
            \state[1] , n43061, \neo_pixel_transmitter.t0 , n29724, 
            n29723, n29722, n29721, n29720, n29719, n29718, n29717, 
            n29716, n29715, n29714, n29713, n29712, n29711, n29710, 
            n29709, n29708, n29707, neopxl_color, n29706, n29705, 
            \state_3__N_528[1] , timer, LED_c, n29323, n29704, n29703, 
            n29702, n29701, n29700, n29699, n29698, n29697, n29696, 
            n29695, n29694, NEOPXL_c, n29633, n29623) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output \state[0] ;
    output \state[1] ;
    output n43061;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input n29724;
    input n29723;
    input n29722;
    input n29721;
    input n29720;
    input n29719;
    input n29718;
    input n29717;
    input n29716;
    input n29715;
    input n29714;
    input n29713;
    input n29712;
    input n29711;
    input n29710;
    input n29709;
    input n29708;
    input n29707;
    input [23:0]neopxl_color;
    input n29706;
    input n29705;
    output \state_3__N_528[1] ;
    output [31:0]timer;
    input LED_c;
    output n29323;
    input n29704;
    input n29703;
    input n29702;
    input n29701;
    input n29700;
    input n29699;
    input n29698;
    input n29697;
    input n29696;
    input n29695;
    input n29694;
    output NEOPXL_c;
    input n29633;
    input n29623;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n2791;
    wire [31:0]n2852;
    
    wire n2819, n2890, n2789, n2888, n2790, n2889, n2788, n2887, 
        n2802, n2901, n2800, n2899, n2795, n2894, n2793, n2892, 
        n2794, n2893, n2792, n2891, n2807, n2906, n2804, n2903, 
        n2787, n2886, n2801, n2900, n2805, n2904, n2803, n2902, 
        n2806, n2905, n2798, n2897;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n2909, n2799, n2898, n2809, n2908, n2808, n2907, n2797, 
        n2896, \neo_pixel_transmitter.done_N_736 , n51572, \neo_pixel_transmitter.done , 
        n2796, n2895, start_N_727, n7, start, n33, n41, n2885, 
        n38, n43, n40, n46, n39, n47, n2918;
    wire [31:0]n971;
    
    wire n39233, n1007, n2, n8;
    wire [31:0]n133;
    
    wire n6801, n29524, n39232, n2702;
    wire [31:0]n2753;
    
    wire n2720, n2708, n2698, n2700, n2688, n2701, n2706, n2703, 
        n2709, n2694, n2692, n2693, n2691, n2697, n2707, n2699, 
        n2704, n2696, n2695, n2690, n2689, n2705, n32, n39_adj_4930, 
        n27833, n4, n41104, n45044, n7_adj_4931, n27992, n45055, 
        n26, n38_adj_4932, n44, n42, n2786, n43_adj_4933, n41_adj_4934, 
        n50168, n49673, n36377, n45052, n50169, n45124, \neo_pixel_transmitter.done_N_742 , 
        n29447, n39231;
    wire [31:0]n1;
    
    wire n2589;
    wire [31:0]n2654;
    
    wire n2621, n2603, n2609, n1205;
    wire [31:0]n1268;
    
    wire n1235, n1304, n1204, n1303, n1207, n1306, n1206, n1305, 
        n40445, n1309, n1209, n1308, n1108;
    wire [31:0]n1169;
    
    wire n1136, n1107, n1106, n1109, n1208, n36229, n1105, n12, 
        n1104, n8_adj_4935, n2606, n2601, n2604, n2600, n2608, 
        n2607, n2602, n2597, n1203, n10, n14, n1202, n2599, 
        n2591, n1302, n1307, n1301, n14_adj_4936, n12_adj_4937, 
        n16, n2593, n1334, n2592, n2590, n2596, n2594, n2598, 
        n2595, n2605, n40444, n30, n37, n36, n42_adj_4938, n40_adj_4939, 
        n2687, n41_adj_4940, n40443, n39_adj_4941, n40442, n2502;
    wire [31:0]n2555;
    
    wire n2522, n2498, n2499, n2503, n2501, n2507, n2500, n2508, 
        n2505, n2504, n2497, n2506, n2492, n2491, n2490, n2496, 
        n2494, n2495, n2493, n2509, n28, n35, n2588, n34, n40_adj_4943, 
        n38_adj_4944, n39_adj_4945, n37_adj_4946, n40441, n2402;
    wire [31:0]n2456;
    
    wire n2423, n2400, n2406, n2408, n2407, n2395, n2393, n2394, 
        n2392, n2399, n2397, n2398, n2396, n2405, n2404, n2409, 
        n2403, n2401, n2391, n2489, n22, n28_adj_4948, n36_adj_4949, 
        n34_adj_4950, n33_adj_4951, n37_adj_4952, n39_adj_4953, n40440, 
        n29401, n39230, n26374, n39229, n40439, n2300;
    wire [31:0]n2357;
    
    wire n2324, n2299, n2308, n2307, n2304, n2302, n2294, n2293, 
        n2292, n2309, n2296, n2297, n2295, n2298, n2306, n40438, 
        n40437, n40436, n40435, n2301, n2305, n40434, n2303, n34_adj_4956, 
        n1400, n39999;
    wire [31:0]n1367;
    
    wire n39998, n25, n32_adj_4957, n40433, n2390, n31, n35_adj_4958, 
        n37_adj_4959, n39997, n39996, n2199;
    wire [31:0]n2258;
    
    wire n2225, n2200, n2198, n2202, n2205, n39995, n2209, n2204, 
        n2207, n2203, n2201, n2206, n2193, n2208, n40432, n2197, 
        n2195, n2196, n2194, n30_adj_4961, n36169, n2291, n34_adj_4962, 
        n32_adj_4963, n33_adj_4964, n31_adj_4965, n39994, n39993, 
        n2100;
    wire [31:0]n2159;
    
    wire n2126, n2107, n2104, n2103, n2099, n2098, n2102, n40431, 
        n2097, n2106, n2105, n2108, n2101, n2109, n2096, n2095, 
        n2094, n2192, n28_adj_4966, n24, n32_adj_4967, n30_adj_4968, 
        n31_adj_4969, n29, n39992, n40430, n48737, n48738, n48879, 
        n48878, n39991, n40429, n40428, n40427, n1999;
    wire [31:0]n2060;
    
    wire n2027, n1997, n1998, n1996, n2004, n2002, n2003, n2005, 
        n2008, n2001, n2000, n2006, n2007, n2009, n40426, n40425, 
        n40424, n1995, n2093, n18_adj_4972, n36165, n40423, n30_adj_4973, 
        n28_adj_4974, n29_adj_4975, n27, n40422, n40421, n1499, 
        n39728, n1433;
    wire [31:0]n1466;
    
    wire n1401, n39727, n1402, n39726, n1403, n39725, n40420, 
        n40419, n1404, n39724, n36085, n48, n46_adj_4977, n47_adj_4978, 
        n45, n40418, n44_adj_4979, n43_adj_4980, n54, n40417, n1405, 
        n39723, n1406, n39722, n40416, n1407, n39721, n1408, n39720, 
        n40415, n1409, n39719, n49;
    wire [31:0]n133_adj_5090;
    
    wire n40414, n40413, n40412, n40411, n40410, n40409, n1923, 
        n40408, n40407;
    wire [3:0]state_3__N_528;
    
    wire n29462, n40406, n49666, n6_adj_4990, n49686, n1900;
    wire [31:0]n1961;
    
    wire n1928, n1901, n1899, n1898, n1897, n1896, n1907, n1902, 
        n1908, n1909, n1905, n1903, n40405, n1904, n1906, n40404, 
        n36163, n28_adj_4993, n40403, n26_adj_4995, n27_adj_4996, 
        n1994, n25_adj_4997, n40402, n40401, n40400, n40399, n40398, 
        n40397, n40396, n40395, n48860, n40394, n48861, n48867, 
        n48866, n40393, n40392, n40391, n40390, n40389, n40388, 
        n40387, n40386, n40385, n40384, n40376, n1805;
    wire [31:0]n1862;
    
    wire n1829, n1803, n1807, n1802, n1801, n1799, n1800, n1798, 
        n1797, n1809, n40375, n40374, n1804, n40373, n1808, n1806, 
        n26_adj_5028, n19_adj_5029, n1895, n16_adj_5030, n24_adj_5031, 
        n28_adj_5032, n40372, n40371, n40370, n40369, n50683, n1037, 
        n40920, n50665, n40919, n1006, n40918, n50661, n40917, 
        n50662, n1008, n40916, n1009, n51353, n40915, n40909, 
        n40908, n40907, n40906, n40905, n40904, n40903, n1697, 
        n1598, n1631, n40902, n1698, n1599, n40901, n1699, n1600, 
        n40900, n1700, n1601, n40899, n1701, n1602, n40898, n1702, 
        n1603, n40897, n1703, n1604, n40896, n1704, n1605, n40895, 
        n1705, n1606, n40894, n1706, n1607, n40893, n1707, n1608, 
        n40892, n1708, n1609, n51354, n40891, n1709, n1796, n40890, 
        n1730;
    wire [31:0]n1763;
    
    wire n40889, n40888, n40887, n40886, n40885, n40884, n40883, 
        n40882, n40881, n40880, n40879, n40878, n40877, n40876, 
        n40875, n40874, n40873, n40872, n40871, n40870, n40869, 
        n40868, n40867, n40866, n40865, n40864, n40863, n40862, 
        n40861, n40860, n40859, n40858, n40857, n40856, n40855, 
        n40854, n40853, n40852, n40851, n40850, n40849, n40848, 
        n40847, n40846, n40845, n40844, n40843, n40842, n40841, 
        n40840, n40839, n40838, n27999, n39279, n48490, n39278, 
        n48488, n40837, n40836, n40835, n40834, n40833, n40832, 
        n40831, n40830, n40829, n40828, n40827, n40826, n40825, 
        n40824, n40823, n40822, n39277, n48486, n40821, n40820, 
        n40819, n39276, n48484, n40818, n39275, n48482, n18_adj_5034, 
        n24_adj_5035, n22_adj_5036, n26_adj_5037, n39274, n48480, 
        n40817, n40816, n40815, n40814, n40813, n40812, n40811, 
        n17_adj_5038, n40810, n21_adj_5039, n20, n24_adj_5040, n40809, 
        n40808, n40807, n40806, n40805, n40804, n40803, n40802, 
        n40801, n40800, n40799, n40798, n40797, n40796, n39273, 
        n48478, n40795, n40794, n40793, n40792, n40791, n39272, 
        n48476, n40790, n40789, n40788, n40787, n40786, n40785, 
        n40784, n40783, n40782, n40781, n40780, n40779, n40778, 
        n40777, n40776, n40775, n40774, n40773, n40772, n40771, 
        n40770, n40769, n39271, n48474, n40768, n40767, n40766, 
        n40765, n40764, n40763, n40762, n39270, n48472, n40761, 
        n40760, n39269, n48470, n40759, n1502;
    wire [31:0]n1565;
    
    wire n1532, n40758, n1501, n40757, n1506, n1500, n39268, n48468, 
        n40756, n40755, n1509, n1507, n1508, n40754, n40753, n40752, 
        n1505, n1503, n1504, n18_adj_5041, n20_adj_5042, n15_adj_5043, 
        n40751, n40750, n40749, n40748, n40747, n40746, n40745, 
        n39267, n48466, n15_adj_5044, n19_adj_5045, n18_adj_5046, 
        n22_adj_5047, n40744, n40743, n40742, n40741, n40740, n40739, 
        n39266, n48464, n40738, n40737, n40736, n39265, n48462, 
        n40735, n40734, n40733, n40732, n40731, n40730, n40729, 
        n40728, n40727, n39264, n48460, n40726, n40725, n40724, 
        n40723, n40722, n40721, n40720, n40719, n40718, n40717, 
        n40716, n39263, n48458, n40715, n40714, n40713, n40712, 
        n40711, n40710, n40709, n40708, n40707, n40706, n40705, 
        n40704, n40703, n40702, n40701, n40700, n40699, n40698, 
        n40697, n39262, n48456;
    wire [31:0]one_wire_N_679;
    
    wire n44921, n48440, n48446, n49688, n45056, n44939, n44187, 
        n103, n16_adj_5048, n6_adj_5049, n40696, n40695, n40694, 
        n40693, n46958, n40692, n40691, n40690, n40689, n40688, 
        n40687, n40686, n40685, n40684, n40683, n40682, n40681, 
        n40680, n40679, n40678, n40677, n40676, n40675, n40674, 
        n40673, n40672, n40671, n40670, n40669, n2984, n40668;
    wire [31:0]n2951;
    
    wire n40667, n40666, n40665, n40664, n40663, n40662, n40661, 
        n40660, n40659, n40658, n40657, n40656, n40655, n40654, 
        n40653, n40652, n40651, n40650, n40649, n40648, n40647, 
        n40646, n40645, n40644, n3083, n40643, n3017;
    wire [31:0]n3050;
    
    wire n2985, n40642, n2986, n40641, n2987, n40640, n2988, n40639, 
        n2989, n40638, n2990, n40637, n2991, n40636, n2992, n40635, 
        n2993, n40634, n2994, n40633, n2995, n40632, n2996, n40631, 
        n2997, n40630, n2998, n40629, n2999, n40628, n3000, n40627, 
        n3001, n40626, n3002, n40625, n3003, n40624, n3004, n40623, 
        n3005, n40622, n3006, n40621, n3007, n40620, n3008, n40619, 
        n32241, n40618, n63, n3116, n40617, n61, n3084, n40616, 
        n59, n3085, n40615, n57, n3086, n40614, n55, n3087, 
        n40613, n53, n3088, n40612, n51, n3089, n40611, n49_adj_5050, 
        n3090, n40610, n47_adj_5051, n3091, n40609, n45_adj_5052, 
        n3092, n40608, n43_adj_5053, n3093, n40607, n39261, n48454, 
        n41_adj_5055, n3094, n40606, n39_adj_5056, n3095, n40605, 
        n37_adj_5057, n3096, n40604, n35_adj_5058, n3097, n40603, 
        n33_adj_5059, n3098, n40602, n31_adj_5060, n3099, n40601, 
        n29_adj_5061, n3100, n40600, n27_adj_5062, n3101, n40599, 
        n25_adj_5063, n3102, n40598, n23_adj_5064, n3103, n40597, 
        n21_adj_5065, n3104, n40596, n19_adj_5066, n3105, n40595, 
        n17_adj_5067, n3106, n40594, n15_adj_5068, n3107, n40593, 
        n13_adj_5069, n3108, n40592, n11_adj_5070, n3109, n51355, 
        n40591, n3209, n48887, n48888, n51417, n48828, n48827, 
        n51420, n39260, n39259, n39258, n39257, n39256, n39255, 
        n39254, n39253, n39252, n51411, n51414, n39251, n39250, 
        n39382, n39381, n39380, n39379, n39378, n39249, n39377, 
        n39376, n39375, n39374, n39373, n39372, n7_adj_5071, n36_adj_5072, 
        n46_adj_5073, n42_adj_5074, n34_adj_5075, n43_adj_5076, n50, 
        n48_adj_5077, n49_adj_5078, n47_adj_5079, n29408, n26382, 
        n35_adj_5080, n43_adj_5081, n40_adj_5082, n45_adj_5083, n42_adj_5084, 
        n48_adj_5085, n41_adj_5086, n49_adj_5087, n48048, n48050, 
        n48052, n48054, n36185, n48062, n48066, n48072, n48078, 
        n41260, n45525;
    wire [4:0]color_bit_N_722;
    
    wire n49685, n51360, n50555, n36189, n16_adj_5088, n17_adj_5089, 
        n51357;
    
    SB_LUT4 mod_5_i1949_3_lut (.I0(n2791), .I1(n2852[26]), .I2(n2819), 
            .I3(GND_net), .O(n2890));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1947_3_lut (.I0(n2789), .I1(n2852[28]), .I2(n2819), 
            .I3(GND_net), .O(n2888));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1948_3_lut (.I0(n2790), .I1(n2852[27]), .I2(n2819), 
            .I3(GND_net), .O(n2889));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1946_3_lut (.I0(n2788), .I1(n2852[29]), .I2(n2819), 
            .I3(GND_net), .O(n2887));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1960_3_lut (.I0(n2802), .I1(n2852[15]), .I2(n2819), 
            .I3(GND_net), .O(n2901));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1958_3_lut (.I0(n2800), .I1(n2852[17]), .I2(n2819), 
            .I3(GND_net), .O(n2899));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1953_3_lut (.I0(n2795), .I1(n2852[22]), .I2(n2819), 
            .I3(GND_net), .O(n2894));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1951_3_lut (.I0(n2793), .I1(n2852[24]), .I2(n2819), 
            .I3(GND_net), .O(n2892));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1952_3_lut (.I0(n2794), .I1(n2852[23]), .I2(n2819), 
            .I3(GND_net), .O(n2893));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1950_3_lut (.I0(n2792), .I1(n2852[25]), .I2(n2819), 
            .I3(GND_net), .O(n2891));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1965_3_lut (.I0(n2807), .I1(n2852[10]), .I2(n2819), 
            .I3(GND_net), .O(n2906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1962_3_lut (.I0(n2804), .I1(n2852[13]), .I2(n2819), 
            .I3(GND_net), .O(n2903));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1945_3_lut (.I0(n2787), .I1(n2852[30]), .I2(n2819), 
            .I3(GND_net), .O(n2886));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1959_3_lut (.I0(n2801), .I1(n2852[16]), .I2(n2819), 
            .I3(GND_net), .O(n2900));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1963_3_lut (.I0(n2805), .I1(n2852[12]), .I2(n2819), 
            .I3(GND_net), .O(n2904));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1961_3_lut (.I0(n2803), .I1(n2852[14]), .I2(n2819), 
            .I3(GND_net), .O(n2902));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1964_3_lut (.I0(n2806), .I1(n2852[11]), .I2(n2819), 
            .I3(GND_net), .O(n2905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1956_3_lut (.I0(n2798), .I1(n2852[19]), .I2(n2819), 
            .I3(GND_net), .O(n2897));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1968_3_lut (.I0(bit_ctr[7]), .I1(n2852[7]), .I2(n2819), 
            .I3(GND_net), .O(n2909));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1957_3_lut (.I0(n2799), .I1(n2852[18]), .I2(n2819), 
            .I3(GND_net), .O(n2898));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1967_3_lut (.I0(n2809), .I1(n2852[8]), .I2(n2819), 
            .I3(GND_net), .O(n2908));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1966_3_lut (.I0(n2808), .I1(n2852[9]), .I2(n2819), 
            .I3(GND_net), .O(n2907));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1955_3_lut (.I0(n2797), .I1(n2852[20]), .I2(n2819), 
            .I3(GND_net), .O(n2896));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1955_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n51572), .D(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1954_3_lut (.I0(n2796), .I1(n2852[21]), .I2(n2819), 
            .I3(GND_net), .O(n2895));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1954_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE start_103 (.Q(start), .C(CLK_c), .E(n7), .D(start_N_727));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2898), .I2(n2909), .I3(GND_net), 
            .O(n33));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut (.I0(n2895), .I1(n2896), .I2(n2907), .I3(n2908), 
            .O(n41));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2900), .I1(n2886), .I2(n2885), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut (.I0(n2897), .I1(n2905), .I2(n2902), .I3(n2904), 
            .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n2891), .I1(n2893), .I2(n2892), .I3(n2894), 
            .O(n40));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n41), .I1(n33), .I2(n2903), .I3(n2906), .O(n46));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2887), .I1(n2889), .I2(n2888), .I3(n2890), 
            .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43), .I1(n2899), .I2(n38), .I3(n2901), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39), .I2(n46), .I3(n40), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n39233), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_3_lut (.I0(n1007), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n8));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_DFFESR bit_ctr_2058__i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n6801), 
            .D(n133[31]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n6801), 
            .D(n133[0]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n6801), 
            .D(n133[30]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n6801), 
            .D(n133[29]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n6801), 
            .D(n133[28]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n6801), 
            .D(n133[27]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n6801), 
            .D(n133[26]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n6801), 
            .D(n133[25]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n6801), 
            .D(n133[24]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n6801), 
            .D(n133[23]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n6801), 
            .D(n133[22]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n39232), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n39232), .I0(GND_net), .I1(VCC_net), 
            .CO(n39233));
    SB_LUT4 mod_5_i1892_3_lut (.I0(n2702), .I1(n2753[16]), .I2(n2720), 
            .I3(GND_net), .O(n2801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1898_3_lut (.I0(n2708), .I1(n2753[10]), .I2(n2720), 
            .I3(GND_net), .O(n2807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1888_3_lut (.I0(n2698), .I1(n2753[20]), .I2(n2720), 
            .I3(GND_net), .O(n2797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1890_3_lut (.I0(n2700), .I1(n2753[18]), .I2(n2720), 
            .I3(GND_net), .O(n2799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1878_3_lut (.I0(n2688), .I1(n2753[30]), .I2(n2720), 
            .I3(GND_net), .O(n2787));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1891_3_lut (.I0(n2701), .I1(n2753[17]), .I2(n2720), 
            .I3(GND_net), .O(n2800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1896_3_lut (.I0(n2706), .I1(n2753[12]), .I2(n2720), 
            .I3(GND_net), .O(n2805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1893_3_lut (.I0(n2703), .I1(n2753[15]), .I2(n2720), 
            .I3(GND_net), .O(n2802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1899_3_lut (.I0(n2709), .I1(n2753[9]), .I2(n2720), 
            .I3(GND_net), .O(n2808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1884_3_lut (.I0(n2694), .I1(n2753[24]), .I2(n2720), 
            .I3(GND_net), .O(n2793));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1882_3_lut (.I0(n2692), .I1(n2753[26]), .I2(n2720), 
            .I3(GND_net), .O(n2791));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1883_3_lut (.I0(n2693), .I1(n2753[25]), .I2(n2720), 
            .I3(GND_net), .O(n2792));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1881_3_lut (.I0(n2691), .I1(n2753[27]), .I2(n2720), 
            .I3(GND_net), .O(n2790));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1887_3_lut (.I0(n2697), .I1(n2753[21]), .I2(n2720), 
            .I3(GND_net), .O(n2796));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1897_3_lut (.I0(n2707), .I1(n2753[11]), .I2(n2720), 
            .I3(GND_net), .O(n2806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1889_3_lut (.I0(n2699), .I1(n2753[19]), .I2(n2720), 
            .I3(GND_net), .O(n2798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1894_3_lut (.I0(n2704), .I1(n2753[14]), .I2(n2720), 
            .I3(GND_net), .O(n2803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1886_3_lut (.I0(n2696), .I1(n2753[22]), .I2(n2720), 
            .I3(GND_net), .O(n2795));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1885_3_lut (.I0(n2695), .I1(n2753[23]), .I2(n2720), 
            .I3(GND_net), .O(n2794));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1880_3_lut (.I0(n2690), .I1(n2753[28]), .I2(n2720), 
            .I3(GND_net), .O(n2789));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1879_3_lut (.I0(n2689), .I1(n2753[29]), .I2(n2720), 
            .I3(GND_net), .O(n2788));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1900_3_lut (.I0(bit_ctr[8]), .I1(n2753[8]), .I2(n2720), 
            .I3(GND_net), .O(n2809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1895_3_lut (.I0(n2705), .I1(n2753[13]), .I2(n2720), 
            .I3(GND_net), .O(n2804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_3_lut_adj_1535 (.I0(n2804), .I1(bit_ctr[7]), .I2(n2809), 
            .I3(GND_net), .O(n32));   // verilog/neopixel.v(22[26:36])
    defparam i8_3_lut_adj_1535.LUT_INIT = 16'heaea;
    SB_LUT4 i15_4_lut_adj_1536 (.I0(n2794), .I1(n2795), .I2(n2803), .I3(n2798), 
            .O(n39_adj_4930));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i29686_4_lut (.I0(n27833), .I1(n4), .I2(n41104), .I3(\state[0] ), 
            .O(n45044));
    defparam i29686_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[1] ), 
            .I2(start), .I3(n45044), .O(n7_adj_4931));
    defparam i20_4_lut.LUT_INIT = 16'hcecf;
    SB_LUT4 i1_4_lut (.I0(n27992), .I1(n7_adj_4931), .I2(n45055), .I3(\state[1] ), 
            .O(n43061));
    defparam i1_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 i2_2_lut (.I0(n2788), .I1(n2789), .I2(GND_net), .I3(GND_net), 
            .O(n26));   // verilog/neopixel.v(22[26:36])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1537 (.I0(n2790), .I1(n2792), .I2(n2791), .I3(n2793), 
            .O(n38_adj_4932));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1538 (.I0(n39_adj_4930), .I1(n2806), .I2(n32), 
            .I3(n2796), .O(n44));   // verilog/neopixel.v(22[26:36])
    defparam i20_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1539 (.I0(n2808), .I1(n2802), .I2(n2805), .I3(n2800), 
            .O(n42));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n2787), .I1(n38_adj_4932), .I2(n26), .I3(n2786), 
            .O(n43_adj_4933));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n2799), .I1(n2797), .I2(n2807), .I3(n2801), 
            .O(n41_adj_4934));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n41_adj_4934), .I1(n43_adj_4933), .I2(n42), 
            .I3(n44), .O(n2819));   // verilog/neopixel.v(22[26:36])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34896_4_lut (.I0(n41104), .I1(n4), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n50168));
    defparam i34896_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n49673), .I1(n36377), .I2(\state[1] ), .I3(n27833), 
            .O(n45052));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n45052), .I1(n50169), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n45124));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i42_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_742 ));
    defparam i42_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n29447), .I2(VCC_net), 
            .I3(n39231), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1811_3_lut (.I0(n2589), .I1(n2654[30]), .I2(n2621), 
            .I3(GND_net), .O(n2688));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1825_3_lut (.I0(n2603), .I1(n2654[16]), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1825_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n6801), 
            .D(n133[21]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1831_3_lut (.I0(n2609), .I1(n2654[10]), .I2(n2621), 
            .I3(GND_net), .O(n2708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i875_3_lut (.I0(n1205), .I1(n1268[28]), .I2(n1235), 
            .I3(GND_net), .O(n1304));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i874_3_lut (.I0(n1204), .I1(n1268[29]), .I2(n1235), 
            .I3(GND_net), .O(n1303));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i877_3_lut (.I0(n1207), .I1(n1268[26]), .I2(n1235), 
            .I3(GND_net), .O(n1306));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i876_3_lut (.I0(n1206), .I1(n1268[27]), .I2(n1235), 
            .I3(GND_net), .O(n1305));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[31]), 
            .I3(n40445), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i880_3_lut (.I0(bit_ctr[23]), .I1(n1268[23]), .I2(n1235), 
            .I3(GND_net), .O(n1309));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i879_3_lut (.I0(n1209), .I1(n1268[24]), .I2(n1235), 
            .I3(GND_net), .O(n1308));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i810_3_lut (.I0(n1108), .I1(n1169[26]), .I2(n1136), 
            .I3(GND_net), .O(n1207));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i809_3_lut (.I0(n1107), .I1(n1169[27]), .I2(n1136), 
            .I3(GND_net), .O(n1206));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i808_3_lut (.I0(n1106), .I1(n1169[28]), .I2(n1136), 
            .I3(GND_net), .O(n1205));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i811_3_lut (.I0(n1109), .I1(n1169[25]), .I2(n1136), 
            .I3(GND_net), .O(n1208));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22709_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n36229));
    defparam i22709_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n36229), .I2(n1106), .I3(n1107), 
            .O(n12));   // verilog/neopixel.v(22[26:36])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1108), .I1(n12), .I2(n1104), .I3(n8_adj_4935), 
            .O(n1136));   // verilog/neopixel.v(22[26:36])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1828_3_lut (.I0(n2606), .I1(n2654[13]), .I2(n2621), 
            .I3(GND_net), .O(n2705));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1823_3_lut (.I0(n2601), .I1(n2654[18]), .I2(n2621), 
            .I3(GND_net), .O(n2700));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1823_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1826_3_lut (.I0(n2604), .I1(n2654[15]), .I2(n2621), 
            .I3(GND_net), .O(n2703));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i807_3_lut (.I0(n1105), .I1(n1169[29]), .I2(n1136), 
            .I3(GND_net), .O(n1204));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1822_3_lut (.I0(n2600), .I1(n2654[19]), .I2(n2621), 
            .I3(GND_net), .O(n2699));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1830_3_lut (.I0(n2608), .I1(n2654[11]), .I2(n2621), 
            .I3(GND_net), .O(n2707));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1829_3_lut (.I0(n2607), .I1(n2654[12]), .I2(n2621), 
            .I3(GND_net), .O(n2706));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1824_3_lut (.I0(n2602), .I1(n2654[17]), .I2(n2621), 
            .I3(GND_net), .O(n2701));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1824_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1819_3_lut (.I0(n2597), .I1(n2654[22]), .I2(n2621), 
            .I3(GND_net), .O(n2696));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i812_3_lut (.I0(bit_ctr[24]), .I1(n1169[24]), .I2(n1136), 
            .I3(GND_net), .O(n1209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), .I3(GND_net), 
            .O(n10));
    defparam i2_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i6_4_lut_adj_1540 (.I0(n1208), .I1(n1205), .I2(n1206), .I3(n1207), 
            .O(n14));
    defparam i6_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n1204), .I1(n14), .I2(n10), .I3(n1202), .O(n1235));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1821_3_lut (.I0(n2599), .I1(n2654[20]), .I2(n2621), 
            .I3(GND_net), .O(n2698));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i806_3_lut (.I0(n1104), .I1(n1169[30]), .I2(n1136), 
            .I3(GND_net), .O(n1203));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1813_3_lut (.I0(n2591), .I1(n2654[28]), .I2(n2621), 
            .I3(GND_net), .O(n2690));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i873_3_lut (.I0(n1203), .I1(n1268[30]), .I2(n1235), 
            .I3(GND_net), .O(n1302));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i878_3_lut (.I0(n1208), .I1(n1268[25]), .I2(n1235), 
            .I3(GND_net), .O(n1307));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(n1307), .I1(n1302), .I2(n1301), .I3(GND_net), 
            .O(n14_adj_4936));   // verilog/neopixel.v(22[26:36])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_2_lut (.I0(n1305), .I1(n1306), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4937));   // verilog/neopixel.v(22[26:36])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1541 (.I0(bit_ctr[22]), .I1(n14_adj_4936), .I2(n1308), 
            .I3(n1309), .O(n16));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1541.LUT_INIT = 16'hfefc;
    SB_LUT4 mod_5_i1815_3_lut (.I0(n2593), .I1(n2654[26]), .I2(n2621), 
            .I3(GND_net), .O(n2692));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut (.I0(n1303), .I1(n16), .I2(n12_adj_4937), .I3(n1304), 
            .O(n1334));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1814_3_lut (.I0(n2592), .I1(n2654[27]), .I2(n2621), 
            .I3(GND_net), .O(n2691));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1812_3_lut (.I0(n2590), .I1(n2654[29]), .I2(n2621), 
            .I3(GND_net), .O(n2689));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1818_3_lut (.I0(n2596), .I1(n2654[23]), .I2(n2621), 
            .I3(GND_net), .O(n2695));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1816_3_lut (.I0(n2594), .I1(n2654[25]), .I2(n2621), 
            .I3(GND_net), .O(n2693));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1816_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1820_3_lut (.I0(n2598), .I1(n2654[21]), .I2(n2621), 
            .I3(GND_net), .O(n2697));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1820_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1817_3_lut (.I0(n2595), .I1(n2654[24]), .I2(n2621), 
            .I3(GND_net), .O(n2694));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1832_3_lut (.I0(bit_ctr[9]), .I1(n2654[9]), .I2(n2621), 
            .I3(GND_net), .O(n2709));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1827_3_lut (.I0(n2605), .I1(n2654[14]), .I2(n2621), 
            .I3(GND_net), .O(n2704));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[30]), 
            .I3(n40444), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_3_lut (.I0(n2704), .I1(bit_ctr[8]), .I2(n2709), .I3(GND_net), 
            .O(n30));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i14_4_lut_adj_1542 (.I0(n2694), .I1(n2697), .I2(n2693), .I3(n2695), 
            .O(n37));
    defparam i14_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_2058__i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n6801), 
            .D(n133[20]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 i13_4_lut (.I0(n2689), .I1(n2691), .I2(n2692), .I3(n2690), 
            .O(n36));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_2058__i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n6801), 
            .D(n133[19]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_CARRY bit_ctr_2058_add_4_32 (.CI(n40444), .I0(GND_net), .I1(bit_ctr[30]), 
            .CO(n40445));
    SB_LUT4 i19_4_lut_adj_1543 (.I0(n37), .I1(n2698), .I2(n30), .I3(n2696), 
            .O(n42_adj_4938));
    defparam i19_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1544 (.I0(n2701), .I1(n2706), .I2(n2707), .I3(n2699), 
            .O(n40_adj_4939));
    defparam i17_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1545 (.I0(n2702), .I1(n36), .I2(n2688), .I3(n2687), 
            .O(n41_adj_4940));
    defparam i18_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_2058_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[29]), 
            .I3(n40443), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_adj_1546 (.I0(n2703), .I1(n2700), .I2(n2705), .I3(n2708), 
            .O(n39_adj_4941));
    defparam i16_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_CARRY bit_ctr_2058_add_4_31 (.CI(n40443), .I0(GND_net), .I1(bit_ctr[29]), 
            .CO(n40444));
    SB_CARRY mod_5_add_669_5 (.CI(n39231), .I0(n29447), .I1(VCC_net), 
            .CO(n39232));
    SB_LUT4 bit_ctr_2058_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[28]), 
            .I3(n40442), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_4_lut_adj_1547 (.I0(n39_adj_4941), .I1(n41_adj_4940), .I2(n40_adj_4939), 
            .I3(n42_adj_4938), .O(n2720));
    defparam i22_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1756_3_lut (.I0(n2502), .I1(n2555[18]), .I2(n2522), 
            .I3(GND_net), .O(n2601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1752_3_lut (.I0(n2498), .I1(n2555[22]), .I2(n2522), 
            .I3(GND_net), .O(n2597));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1753_3_lut (.I0(n2499), .I1(n2555[21]), .I2(n2522), 
            .I3(GND_net), .O(n2598));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1757_3_lut (.I0(n2503), .I1(n2555[17]), .I2(n2522), 
            .I3(GND_net), .O(n2602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1755_3_lut (.I0(n2501), .I1(n2555[19]), .I2(n2522), 
            .I3(GND_net), .O(n2600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1761_3_lut (.I0(n2507), .I1(n2555[13]), .I2(n2522), 
            .I3(GND_net), .O(n2606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1761_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1754_3_lut (.I0(n2500), .I1(n2555[20]), .I2(n2522), 
            .I3(GND_net), .O(n2599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1762_3_lut (.I0(n2508), .I1(n2555[12]), .I2(n2522), 
            .I3(GND_net), .O(n2607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1759_3_lut (.I0(n2505), .I1(n2555[15]), .I2(n2522), 
            .I3(GND_net), .O(n2604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1758_3_lut (.I0(n2504), .I1(n2555[16]), .I2(n2522), 
            .I3(GND_net), .O(n2603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1751_3_lut (.I0(n2497), .I1(n2555[23]), .I2(n2522), 
            .I3(GND_net), .O(n2596));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY bit_ctr_2058_add_4_30 (.CI(n40442), .I0(GND_net), .I1(bit_ctr[28]), 
            .CO(n40443));
    SB_LUT4 mod_5_i1760_3_lut (.I0(n2506), .I1(n2555[14]), .I2(n2522), 
            .I3(GND_net), .O(n2605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1746_3_lut (.I0(n2492), .I1(n2555[28]), .I2(n2522), 
            .I3(GND_net), .O(n2591));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1745_3_lut (.I0(n2491), .I1(n2555[29]), .I2(n2522), 
            .I3(GND_net), .O(n2590));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1744_3_lut (.I0(n2490), .I1(n2555[30]), .I2(n2522), 
            .I3(GND_net), .O(n2589));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1750_3_lut (.I0(n2496), .I1(n2555[24]), .I2(n2522), 
            .I3(GND_net), .O(n2595));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1748_3_lut (.I0(n2494), .I1(n2555[26]), .I2(n2522), 
            .I3(GND_net), .O(n2593));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1749_3_lut (.I0(n2495), .I1(n2555[25]), .I2(n2522), 
            .I3(GND_net), .O(n2594));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1747_3_lut (.I0(n2493), .I1(n2555[27]), .I2(n2522), 
            .I3(GND_net), .O(n2592));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1764_3_lut (.I0(bit_ctr[10]), .I1(n2555[10]), .I2(n2522), 
            .I3(GND_net), .O(n2609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1763_3_lut (.I0(n2509), .I1(n2555[11]), .I2(n2522), 
            .I3(GND_net), .O(n2608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(bit_ctr[9]), .I1(n2608), .I2(n2609), .I3(GND_net), 
            .O(n28));   // verilog/neopixel.v(22[26:36])
    defparam i6_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1548 (.I0(n2592), .I1(n2594), .I2(n2593), .I3(n2595), 
            .O(n35));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2589), .I1(n2590), .I2(n2588), .I3(n2591), 
            .O(n34));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1549 (.I0(n35), .I1(n2605), .I2(n28), .I3(n2596), 
            .O(n40_adj_4943));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1550 (.I0(n2603), .I1(n2604), .I2(n2607), .I3(n2599), 
            .O(n38_adj_4944));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2606), .I1(n34), .I2(n2600), .I3(GND_net), 
            .O(n39_adj_4945));   // verilog/neopixel.v(22[26:36])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1551 (.I0(n2602), .I1(n2598), .I2(n2597), .I3(n2601), 
            .O(n37_adj_4946));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1552 (.I0(n37_adj_4946), .I1(n39_adj_4945), .I2(n38_adj_4944), 
            .I3(n40_adj_4943), .O(n2621));   // verilog/neopixel.v(22[26:36])
    defparam i21_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2058_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[27]), 
            .I3(n40441), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1688_3_lut (.I0(n2402), .I1(n2456[19]), .I2(n2423), 
            .I3(GND_net), .O(n2501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1686_3_lut (.I0(n2400), .I1(n2456[21]), .I2(n2423), 
            .I3(GND_net), .O(n2499));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1692_3_lut (.I0(n2406), .I1(n2456[15]), .I2(n2423), 
            .I3(GND_net), .O(n2505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1694_3_lut (.I0(n2408), .I1(n2456[13]), .I2(n2423), 
            .I3(GND_net), .O(n2507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1693_3_lut (.I0(n2407), .I1(n2456[14]), .I2(n2423), 
            .I3(GND_net), .O(n2506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1681_3_lut (.I0(n2395), .I1(n2456[26]), .I2(n2423), 
            .I3(GND_net), .O(n2494));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1679_3_lut (.I0(n2393), .I1(n2456[28]), .I2(n2423), 
            .I3(GND_net), .O(n2492));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1680_3_lut (.I0(n2394), .I1(n2456[27]), .I2(n2423), 
            .I3(GND_net), .O(n2493));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1678_3_lut (.I0(n2392), .I1(n2456[29]), .I2(n2423), 
            .I3(GND_net), .O(n2491));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1685_3_lut (.I0(n2399), .I1(n2456[22]), .I2(n2423), 
            .I3(GND_net), .O(n2498));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1683_3_lut (.I0(n2397), .I1(n2456[24]), .I2(n2423), 
            .I3(GND_net), .O(n2496));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1684_3_lut (.I0(n2398), .I1(n2456[23]), .I2(n2423), 
            .I3(GND_net), .O(n2497));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1682_3_lut (.I0(n2396), .I1(n2456[25]), .I2(n2423), 
            .I3(GND_net), .O(n2495));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1691_3_lut (.I0(n2405), .I1(n2456[16]), .I2(n2423), 
            .I3(GND_net), .O(n2504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1690_3_lut (.I0(n2404), .I1(n2456[17]), .I2(n2423), 
            .I3(GND_net), .O(n2503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1695_3_lut (.I0(n2409), .I1(n2456[12]), .I2(n2423), 
            .I3(GND_net), .O(n2508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1689_3_lut (.I0(n2403), .I1(n2456[18]), .I2(n2423), 
            .I3(GND_net), .O(n2502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1689_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY bit_ctr_2058_add_4_29 (.CI(n40441), .I0(GND_net), .I1(bit_ctr[27]), 
            .CO(n40442));
    SB_LUT4 mod_5_i1696_3_lut (.I0(bit_ctr[11]), .I1(n2456[11]), .I2(n2423), 
            .I3(GND_net), .O(n2509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1687_3_lut (.I0(n2401), .I1(n2456[20]), .I2(n2423), 
            .I3(GND_net), .O(n2500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1677_3_lut (.I0(n2391), .I1(n2456[30]), .I2(n2423), 
            .I3(GND_net), .O(n2490));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n2490), .I1(n2489), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_3_lut_adj_1553 (.I0(bit_ctr[10]), .I1(n2500), .I2(n2509), 
            .I3(GND_net), .O(n28_adj_4948));
    defparam i7_3_lut_adj_1553.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1554 (.I0(n2502), .I1(n2508), .I2(n2503), .I3(n2504), 
            .O(n36_adj_4949));
    defparam i15_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1555 (.I0(n2495), .I1(n2497), .I2(n2496), .I3(n2498), 
            .O(n34_adj_4950));
    defparam i13_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1556 (.I0(n2491), .I1(n2493), .I2(n2492), .I3(n2494), 
            .O(n33_adj_4951));
    defparam i12_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1557 (.I0(n2506), .I1(n2507), .I2(n2505), .I3(n22), 
            .O(n37_adj_4952));
    defparam i16_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1558 (.I0(n2499), .I1(n36_adj_4949), .I2(n28_adj_4948), 
            .I3(n2501), .O(n39_adj_4953));
    defparam i18_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1559 (.I0(n39_adj_4953), .I1(n37_adj_4952), .I2(n33_adj_4951), 
            .I3(n34_adj_4950), .O(n2522));
    defparam i20_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_2058__i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n6801), 
            .D(n133[18]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2058_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[26]), 
            .I3(n40440), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n29401), .I2(VCC_net), 
            .I3(n39230), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_28 (.CI(n40440), .I0(GND_net), .I1(bit_ctr[26]), 
            .CO(n40441));
    SB_CARRY mod_5_add_669_4 (.CI(n39230), .I0(n29401), .I1(VCC_net), 
            .CO(n39231));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n26374), .I2(GND_net), 
            .I3(n39229), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_2058_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[25]), 
            .I3(n40439), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_669_3 (.CI(n39229), .I0(n26374), .I1(GND_net), 
            .CO(n39230));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1618_3_lut (.I0(n2300), .I1(n2357[22]), .I2(n2324), 
            .I3(GND_net), .O(n2399));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1617_3_lut (.I0(n2299), .I1(n2357[23]), .I2(n2324), 
            .I3(GND_net), .O(n2398));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1617_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n6801), 
            .D(n133[17]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFFESR bit_ctr_2058__i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n6801), 
            .D(n133[16]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_CARRY bit_ctr_2058_add_4_27 (.CI(n40439), .I0(GND_net), .I1(bit_ctr[25]), 
            .CO(n40440));
    SB_LUT4 mod_5_i1626_3_lut (.I0(n2308), .I1(n2357[14]), .I2(n2324), 
            .I3(GND_net), .O(n2407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1625_3_lut (.I0(n2307), .I1(n2357[15]), .I2(n2324), 
            .I3(GND_net), .O(n2406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1622_3_lut (.I0(n2304), .I1(n2357[18]), .I2(n2324), 
            .I3(GND_net), .O(n2403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1620_3_lut (.I0(n2302), .I1(n2357[20]), .I2(n2324), 
            .I3(GND_net), .O(n2401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1612_3_lut (.I0(n2294), .I1(n2357[28]), .I2(n2324), 
            .I3(GND_net), .O(n2393));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1611_3_lut (.I0(n2293), .I1(n2357[29]), .I2(n2324), 
            .I3(GND_net), .O(n2392));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1610_3_lut (.I0(n2292), .I1(n2357[30]), .I2(n2324), 
            .I3(GND_net), .O(n2391));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1627_3_lut (.I0(n2309), .I1(n2357[13]), .I2(n2324), 
            .I3(GND_net), .O(n2408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1614_3_lut (.I0(n2296), .I1(n2357[26]), .I2(n2324), 
            .I3(GND_net), .O(n2395));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1615_3_lut (.I0(n2297), .I1(n2357[25]), .I2(n2324), 
            .I3(GND_net), .O(n2396));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1613_3_lut (.I0(n2295), .I1(n2357[27]), .I2(n2324), 
            .I3(GND_net), .O(n2394));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1628_3_lut (.I0(bit_ctr[12]), .I1(n2357[12]), .I2(n2324), 
            .I3(GND_net), .O(n2409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1616_3_lut (.I0(n2298), .I1(n2357[24]), .I2(n2324), 
            .I3(GND_net), .O(n2397));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1624_3_lut (.I0(n2306), .I1(n2357[16]), .I2(n2324), 
            .I3(GND_net), .O(n2405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[24]), 
            .I3(n40438), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_26 (.CI(n40438), .I0(GND_net), .I1(bit_ctr[24]), 
            .CO(n40439));
    SB_LUT4 bit_ctr_2058_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[23]), 
            .I3(n40437), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_25 (.CI(n40437), .I0(GND_net), .I1(bit_ctr[23]), 
            .CO(n40438));
    SB_LUT4 bit_ctr_2058_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[22]), 
            .I3(n40436), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_24 (.CI(n40436), .I0(GND_net), .I1(bit_ctr[22]), 
            .CO(n40437));
    SB_LUT4 bit_ctr_2058_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[21]), 
            .I3(n40435), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_23 (.CI(n40435), .I0(GND_net), .I1(bit_ctr[21]), 
            .CO(n40436));
    SB_DFFESR bit_ctr_2058__i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n6801), 
            .D(n133[15]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1619_3_lut (.I0(n2301), .I1(n2357[21]), .I2(n2324), 
            .I3(GND_net), .O(n2400));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1623_3_lut (.I0(n2305), .I1(n2357[17]), .I2(n2324), 
            .I3(GND_net), .O(n2404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[20]), 
            .I3(n40434), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1621_3_lut (.I0(n2303), .I1(n2357[19]), .I2(n2324), 
            .I3(GND_net), .O(n2402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1621_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY bit_ctr_2058_add_4_22 (.CI(n40434), .I0(GND_net), .I1(bit_ctr[20]), 
            .CO(n40435));
    SB_LUT4 i14_4_lut_adj_1560 (.I0(n2402), .I1(n2404), .I2(n2400), .I3(n2405), 
            .O(n34_adj_4956));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1334), .I1(n1301), .I2(VCC_net), 
            .I3(n39999), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_10_lut (.I0(GND_net), .I1(n1302), .I2(VCC_net), 
            .I3(n39998), .O(n1367[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_3_lut_adj_1561 (.I0(n2397), .I1(bit_ctr[11]), .I2(n2409), 
            .I3(GND_net), .O(n25));   // verilog/neopixel.v(22[26:36])
    defparam i5_3_lut_adj_1561.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1562 (.I0(n2394), .I1(n2396), .I2(n2395), .I3(n2408), 
            .O(n32_adj_4957));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_2058_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[19]), 
            .I3(n40433), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_10 (.CI(n39998), .I0(n1302), .I1(VCC_net), 
            .CO(n39999));
    SB_LUT4 i11_4_lut (.I0(n2391), .I1(n2392), .I2(n2390), .I3(n2393), 
            .O(n31));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY bit_ctr_2058_add_4_21 (.CI(n40433), .I0(GND_net), .I1(bit_ctr[19]), 
            .CO(n40434));
    SB_LUT4 i15_4_lut_adj_1563 (.I0(n2401), .I1(n2403), .I2(n2406), .I3(n2407), 
            .O(n35_adj_4958));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1564 (.I0(n25), .I1(n34_adj_4956), .I2(n2398), 
            .I3(n2399), .O(n37_adj_4959));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_9_lut (.I0(GND_net), .I1(n1303), .I2(VCC_net), 
            .I3(n39997), .O(n1367[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_9 (.CI(n39997), .I0(n1303), .I1(VCC_net), .CO(n39998));
    SB_LUT4 i19_4_lut_adj_1565 (.I0(n37_adj_4959), .I1(n35_adj_4958), .I2(n31), 
            .I3(n32_adj_4957), .O(n2423));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_8_lut (.I0(GND_net), .I1(n1304), .I2(VCC_net), 
            .I3(n39996), .O(n1367[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n29724));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1549_3_lut (.I0(n2199), .I1(n2258[24]), .I2(n2225), 
            .I3(GND_net), .O(n2298));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1550_3_lut (.I0(n2200), .I1(n2258[23]), .I2(n2225), 
            .I3(GND_net), .O(n2299));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1548_3_lut (.I0(n2198), .I1(n2258[25]), .I2(n2225), 
            .I3(GND_net), .O(n2297));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1552_3_lut (.I0(n2202), .I1(n2258[21]), .I2(n2225), 
            .I3(GND_net), .O(n2301));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1552_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n29723));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_937_8 (.CI(n39996), .I0(n1304), .I1(VCC_net), .CO(n39997));
    SB_LUT4 mod_5_i1555_3_lut (.I0(n2205), .I1(n2258[18]), .I2(n2225), 
            .I3(GND_net), .O(n2304));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_937_7_lut (.I0(GND_net), .I1(n1305), .I2(VCC_net), 
            .I3(n39995), .O(n1367[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1559_3_lut (.I0(n2209), .I1(n2258[14]), .I2(n2225), 
            .I3(GND_net), .O(n2308));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1554_3_lut (.I0(n2204), .I1(n2258[19]), .I2(n2225), 
            .I3(GND_net), .O(n2303));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1557_3_lut (.I0(n2207), .I1(n2258[16]), .I2(n2225), 
            .I3(GND_net), .O(n2306));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1553_3_lut (.I0(n2203), .I1(n2258[20]), .I2(n2225), 
            .I3(GND_net), .O(n2302));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1551_3_lut (.I0(n2201), .I1(n2258[22]), .I2(n2225), 
            .I3(GND_net), .O(n2300));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1556_3_lut (.I0(n2206), .I1(n2258[17]), .I2(n2225), 
            .I3(GND_net), .O(n2305));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1543_3_lut (.I0(n2193), .I1(n2258[30]), .I2(n2225), 
            .I3(GND_net), .O(n2292));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1558_3_lut (.I0(n2208), .I1(n2258[15]), .I2(n2225), 
            .I3(GND_net), .O(n2307));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1560_3_lut (.I0(bit_ctr[13]), .I1(n2258[13]), .I2(n2225), 
            .I3(GND_net), .O(n2309));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[18]), 
            .I3(n40432), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1547_3_lut (.I0(n2197), .I1(n2258[26]), .I2(n2225), 
            .I3(GND_net), .O(n2296));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1545_3_lut (.I0(n2195), .I1(n2258[28]), .I2(n2225), 
            .I3(GND_net), .O(n2294));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1546_3_lut (.I0(n2196), .I1(n2258[27]), .I2(n2225), 
            .I3(GND_net), .O(n2295));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1544_3_lut (.I0(n2194), .I1(n2258[29]), .I2(n2225), 
            .I3(GND_net), .O(n2293));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1566 (.I0(n2293), .I1(n2295), .I2(n2294), .I3(n2296), 
            .O(n30_adj_4961));
    defparam i11_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i22651_2_lut (.I0(bit_ctr[12]), .I1(n2309), .I2(GND_net), 
            .I3(GND_net), .O(n36169));
    defparam i22651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15_4_lut_adj_1567 (.I0(n2307), .I1(n30_adj_4961), .I2(n2292), 
            .I3(n2291), .O(n34_adj_4962));
    defparam i15_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_937_7 (.CI(n39995), .I0(n1305), .I1(VCC_net), .CO(n39996));
    SB_LUT4 i13_4_lut_adj_1568 (.I0(n2305), .I1(n2300), .I2(n2302), .I3(n2306), 
            .O(n32_adj_4963));
    defparam i13_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_CARRY bit_ctr_2058_add_4_20 (.CI(n40432), .I0(GND_net), .I1(bit_ctr[18]), 
            .CO(n40433));
    SB_LUT4 i14_4_lut_adj_1569 (.I0(n2303), .I1(n2308), .I2(n2304), .I3(n2301), 
            .O(n33_adj_4964));
    defparam i14_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1570 (.I0(n2297), .I1(n2299), .I2(n2298), .I3(n36169), 
            .O(n31_adj_4965));
    defparam i12_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n29722));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_2058__i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n6801), 
            .D(n133[14]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n29721));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i18_4_lut_adj_1571 (.I0(n31_adj_4965), .I1(n33_adj_4964), .I2(n32_adj_4963), 
            .I3(n34_adj_4962), .O(n2324));
    defparam i18_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n29720));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n29719));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n29718));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n29717));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n29716));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n29715));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n29714));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n29713));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n29712));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_6_lut (.I0(GND_net), .I1(n1306), .I2(VCC_net), 
            .I3(n39994), .O(n1367[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n29711));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n29710));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n29709));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_937_6 (.CI(n39994), .I0(n1306), .I1(VCC_net), .CO(n39995));
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n29708));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n29707));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_5_lut (.I0(GND_net), .I1(n1307), .I2(VCC_net), 
            .I3(n39993), .O(n1367[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_5 (.CI(n39993), .I0(n1307), .I1(VCC_net), .CO(n39994));
    SB_LUT4 mod_5_i1482_3_lut (.I0(n2100), .I1(n2159[24]), .I2(n2126), 
            .I3(GND_net), .O(n2199));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1489_3_lut (.I0(n2107), .I1(n2159[17]), .I2(n2126), 
            .I3(GND_net), .O(n2206));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1486_3_lut (.I0(n2104), .I1(n2159[20]), .I2(n2126), 
            .I3(GND_net), .O(n2203));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1485_3_lut (.I0(n2103), .I1(n2159[21]), .I2(n2126), 
            .I3(GND_net), .O(n2202));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1481_3_lut (.I0(n2099), .I1(n2159[25]), .I2(n2126), 
            .I3(GND_net), .O(n2198));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1480_3_lut (.I0(n2098), .I1(n2159[26]), .I2(n2126), 
            .I3(GND_net), .O(n2197));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1480_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n6801), 
            .D(n133[13]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1484_3_lut (.I0(n2102), .I1(n2159[22]), .I2(n2126), 
            .I3(GND_net), .O(n2201));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1484_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR bit_ctr_2058__i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n6801), 
            .D(n133[12]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 bit_ctr_2058_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[17]), 
            .I3(n40431), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_19 (.CI(n40431), .I0(GND_net), .I1(bit_ctr[17]), 
            .CO(n40432));
    SB_LUT4 mod_5_i1479_3_lut (.I0(n2097), .I1(n2159[27]), .I2(n2126), 
            .I3(GND_net), .O(n2196));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1492_3_lut (.I0(bit_ctr[14]), .I1(n2159[14]), .I2(n2126), 
            .I3(GND_net), .O(n2209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1488_3_lut (.I0(n2106), .I1(n2159[18]), .I2(n2126), 
            .I3(GND_net), .O(n2205));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1487_3_lut (.I0(n2105), .I1(n2159[19]), .I2(n2126), 
            .I3(GND_net), .O(n2204));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1490_3_lut (.I0(n2108), .I1(n2159[16]), .I2(n2126), 
            .I3(GND_net), .O(n2207));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1483_3_lut (.I0(n2101), .I1(n2159[23]), .I2(n2126), 
            .I3(GND_net), .O(n2200));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1491_3_lut (.I0(n2109), .I1(n2159[15]), .I2(n2126), 
            .I3(GND_net), .O(n2208));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1478_3_lut (.I0(n2096), .I1(n2159[28]), .I2(n2126), 
            .I3(GND_net), .O(n2195));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1477_3_lut (.I0(n2095), .I1(n2159[29]), .I2(n2126), 
            .I3(GND_net), .O(n2194));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1476_3_lut (.I0(n2094), .I1(n2159[30]), .I2(n2126), 
            .I3(GND_net), .O(n2193));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut (.I0(n2193), .I1(n2194), .I2(n2192), .I3(n2195), 
            .O(n28_adj_4966));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n2208), .I1(n2200), .I2(GND_net), .I3(GND_net), 
            .O(n24));   // verilog/neopixel.v(22[26:36])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_3_lut (.I0(n2207), .I1(n28_adj_4966), .I2(n2204), .I3(GND_net), 
            .O(n32_adj_4967));   // verilog/neopixel.v(22[26:36])
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1572 (.I0(bit_ctr[13]), .I1(n24), .I2(n2205), 
            .I3(n2209), .O(n30_adj_4968));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1572.LUT_INIT = 16'hfefc;
    SB_LUT4 i13_4_lut_adj_1573 (.I0(n2202), .I1(n2203), .I2(n2206), .I3(n2199), 
            .O(n31_adj_4969));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1574 (.I0(n2196), .I1(n2201), .I2(n2197), .I3(n2198), 
            .O(n29));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1575 (.I0(n29), .I1(n31_adj_4969), .I2(n30_adj_4968), 
            .I3(n32_adj_4967), .O(n2225));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_4_lut (.I0(GND_net), .I1(n1308), .I2(VCC_net), 
            .I3(n39992), .O(n1367[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_2058_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[16]), 
            .I3(n40430), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_4 (.CI(n39992), .I0(n1308), .I1(VCC_net), .CO(n39993));
    SB_LUT4 i33300_3_lut (.I0(neopxl_color[0]), .I1(neopxl_color[1]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48737));
    defparam i33300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33301_3_lut (.I0(neopxl_color[2]), .I1(neopxl_color[3]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48738));
    defparam i33301_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n39229));
    SB_LUT4 i33442_3_lut (.I0(neopxl_color[6]), .I1(neopxl_color[7]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48879));
    defparam i33442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33441_3_lut (.I0(neopxl_color[4]), .I1(neopxl_color[5]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48878));
    defparam i33441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY bit_ctr_2058_add_4_18 (.CI(n40430), .I0(GND_net), .I1(bit_ctr[16]), 
            .CO(n40431));
    SB_LUT4 mod_5_add_937_3_lut (.I0(GND_net), .I1(n1309), .I2(GND_net), 
            .I3(n39991), .O(n1367[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_2058_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[15]), 
            .I3(n40429), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_3 (.CI(n39991), .I0(n1309), .I1(GND_net), .CO(n39992));
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_937_2_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(VCC_net), .O(n1367[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(GND_net), 
            .CO(n39991));
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY bit_ctr_2058_add_4_17 (.CI(n40429), .I0(GND_net), .I1(bit_ctr[15]), 
            .CO(n40430));
    SB_LUT4 bit_ctr_2058_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[14]), 
            .I3(n40428), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n29706));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n29705));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY bit_ctr_2058_add_4_16 (.CI(n40428), .I0(GND_net), .I1(bit_ctr[14]), 
            .CO(n40429));
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_2058_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[13]), 
            .I3(n40427), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_15 (.CI(n40427), .I0(GND_net), .I1(bit_ctr[13]), 
            .CO(n40428));
    SB_DFFESR bit_ctr_2058__i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n6801), 
            .D(n133[11]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_i1413_3_lut (.I0(n1999), .I1(n2060[26]), .I2(n2027), 
            .I3(GND_net), .O(n2098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1411_3_lut (.I0(n1997), .I1(n2060[28]), .I2(n2027), 
            .I3(GND_net), .O(n2096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1412_3_lut (.I0(n1998), .I1(n2060[27]), .I2(n2027), 
            .I3(GND_net), .O(n2097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1410_3_lut (.I0(n1996), .I1(n2060[29]), .I2(n2027), 
            .I3(GND_net), .O(n2095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1418_3_lut (.I0(n2004), .I1(n2060[21]), .I2(n2027), 
            .I3(GND_net), .O(n2103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1416_3_lut (.I0(n2002), .I1(n2060[23]), .I2(n2027), 
            .I3(GND_net), .O(n2101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1417_3_lut (.I0(n2003), .I1(n2060[22]), .I2(n2027), 
            .I3(GND_net), .O(n2102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1419_3_lut (.I0(n2005), .I1(n2060[20]), .I2(n2027), 
            .I3(GND_net), .O(n2104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1422_3_lut (.I0(n2008), .I1(n2060[17]), .I2(n2027), 
            .I3(GND_net), .O(n2107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1415_3_lut (.I0(n2001), .I1(n2060[24]), .I2(n2027), 
            .I3(GND_net), .O(n2100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1414_3_lut (.I0(n2000), .I1(n2060[25]), .I2(n2027), 
            .I3(GND_net), .O(n2099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1420_3_lut (.I0(n2006), .I1(n2060[19]), .I2(n2027), 
            .I3(GND_net), .O(n2105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1421_3_lut (.I0(n2007), .I1(n2060[18]), .I2(n2027), 
            .I3(GND_net), .O(n2106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1423_3_lut (.I0(n2009), .I1(n2060[16]), .I2(n2027), 
            .I3(GND_net), .O(n2108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_ctr_2058_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[12]), 
            .I3(n40426), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_14 (.CI(n40426), .I0(GND_net), .I1(bit_ctr[12]), 
            .CO(n40427));
    SB_LUT4 bit_ctr_2058_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[11]), 
            .I3(n40425), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1424_3_lut (.I0(bit_ctr[15]), .I1(n2060[15]), .I2(n2027), 
            .I3(GND_net), .O(n2109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1424_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY bit_ctr_2058_add_4_13 (.CI(n40425), .I0(GND_net), .I1(bit_ctr[11]), 
            .CO(n40426));
    SB_LUT4 bit_ctr_2058_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[10]), 
            .I3(n40424), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1409_3_lut (.I0(n1995), .I1(n2060[30]), .I2(n2027), 
            .I3(GND_net), .O(n2094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY bit_ctr_2058_add_4_12 (.CI(n40424), .I0(GND_net), .I1(bit_ctr[10]), 
            .CO(n40425));
    SB_LUT4 i1_2_lut_adj_1576 (.I0(n2094), .I1(n2093), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4972));
    defparam i1_2_lut_adj_1576.LUT_INIT = 16'heeee;
    SB_LUT4 i22647_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n36165));
    defparam i22647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 bit_ctr_2058_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[9]), 
            .I3(n40423), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut_adj_1577 (.I0(n2108), .I1(n2106), .I2(n2105), .I3(n18_adj_4972), 
            .O(n30_adj_4973));
    defparam i13_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_CARRY bit_ctr_2058_add_4_11 (.CI(n40423), .I0(GND_net), .I1(bit_ctr[9]), 
            .CO(n40424));
    SB_LUT4 i11_4_lut_adj_1578 (.I0(n2099), .I1(n36165), .I2(n2100), .I3(n2107), 
            .O(n28_adj_4974));
    defparam i11_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1579 (.I0(n2104), .I1(n2102), .I2(n2101), .I3(n2103), 
            .O(n29_adj_4975));
    defparam i12_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1580 (.I0(n2095), .I1(n2097), .I2(n2096), .I3(n2098), 
            .O(n27));
    defparam i10_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1581 (.I0(n27), .I1(n29_adj_4975), .I2(n28_adj_4974), 
            .I3(n30_adj_4973), .O(n2126));
    defparam i16_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_2058_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[8]), 
            .I3(n40422), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_10 (.CI(n40422), .I0(GND_net), .I1(bit_ctr[8]), 
            .CO(n40423));
    SB_LUT4 bit_ctr_2058_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[7]), 
            .I3(n40421), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1433), .I1(n1400), .I2(VCC_net), 
            .I3(n39728), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_ctr_2058_add_4_9 (.CI(n40421), .I0(GND_net), .I1(bit_ctr[7]), 
            .CO(n40422));
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(GND_net), .I1(n1401), .I2(VCC_net), 
            .I3(n39727), .O(n1466[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_11 (.CI(n39727), .I0(n1401), .I1(VCC_net), 
            .CO(n39728));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(GND_net), .I1(n1402), .I2(VCC_net), 
            .I3(n39726), .O(n1466[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_10 (.CI(n39726), .I0(n1402), .I1(VCC_net), 
            .CO(n39727));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(GND_net), .I1(n1403), .I2(VCC_net), 
            .I3(n39725), .O(n1466[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_2058_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[6]), 
            .I3(n40420), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_9 (.CI(n39725), .I0(n1403), .I1(VCC_net), 
            .CO(n39726));
    SB_CARRY bit_ctr_2058_add_4_8 (.CI(n40420), .I0(GND_net), .I1(bit_ctr[6]), 
            .CO(n40421));
    SB_LUT4 bit_ctr_2058_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[5]), 
            .I3(n40419), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_7 (.CI(n40419), .I0(GND_net), .I1(bit_ctr[5]), 
            .CO(n40420));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(GND_net), .I1(n1404), .I2(VCC_net), 
            .I3(n39724), .O(n1466[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_8 (.CI(n39724), .I0(n1404), .I1(VCC_net), 
            .CO(n39725));
    SB_LUT4 i22569_2_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(GND_net), .O(n36085));
    defparam i22569_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1582 (.I0(bit_ctr[8]), .I1(bit_ctr[18]), .I2(bit_ctr[24]), 
            .I3(bit_ctr[9]), .O(n48));
    defparam i20_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1583 (.I0(bit_ctr[26]), .I1(bit_ctr[28]), .I2(bit_ctr[6]), 
            .I3(bit_ctr[19]), .O(n46_adj_4977));
    defparam i18_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1584 (.I0(bit_ctr[13]), .I1(bit_ctr[20]), .I2(bit_ctr[23]), 
            .I3(bit_ctr[16]), .O(n47_adj_4978));
    defparam i19_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1585 (.I0(bit_ctr[15]), .I1(bit_ctr[14]), .I2(bit_ctr[21]), 
            .I3(bit_ctr[22]), .O(n45));
    defparam i17_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_2058_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[4]), 
            .I3(n40418), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_adj_1586 (.I0(bit_ctr[11]), .I1(bit_ctr[7]), .I2(bit_ctr[17]), 
            .I3(bit_ctr[29]), .O(n44_adj_4979));
    defparam i16_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1587 (.I0(bit_ctr[12]), .I1(bit_ctr[30]), .I2(n36085), 
            .I3(bit_ctr[25]), .O(n43_adj_4980));
    defparam i15_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47_adj_4978), .I2(n46_adj_4977), 
            .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY bit_ctr_2058_add_4_6 (.CI(n40418), .I0(GND_net), .I1(bit_ctr[4]), 
            .CO(n40419));
    SB_LUT4 bit_ctr_2058_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[3]), 
            .I3(n40417), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_7_lut (.I0(GND_net), .I1(n1405), .I2(VCC_net), 
            .I3(n39723), .O(n1466[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_7 (.CI(n39723), .I0(n1405), .I1(VCC_net), 
            .CO(n39724));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(GND_net), .I1(n1406), .I2(VCC_net), 
            .I3(n39722), .O(n1466[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_5 (.CI(n40417), .I0(GND_net), .I1(bit_ctr[3]), 
            .CO(n40418));
    SB_CARRY mod_5_add_1004_6 (.CI(n39722), .I0(n1406), .I1(VCC_net), 
            .CO(n39723));
    SB_LUT4 bit_ctr_2058_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[2]), 
            .I3(n40416), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_5_lut (.I0(GND_net), .I1(n1407), .I2(VCC_net), 
            .I3(n39721), .O(n1466[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_4 (.CI(n40416), .I0(GND_net), .I1(bit_ctr[2]), 
            .CO(n40417));
    SB_CARRY mod_5_add_1004_5 (.CI(n39721), .I0(n1407), .I1(VCC_net), 
            .CO(n39722));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(GND_net), .I1(n1408), .I2(VCC_net), 
            .I3(n39720), .O(n1466[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_2058_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[1]), 
            .I3(n40415), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_4 (.CI(n39720), .I0(n1408), .I1(VCC_net), 
            .CO(n39721));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(GND_net), .I1(n1409), .I2(GND_net), 
            .I3(n39719), .O(n1466[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_ctr_2058_add_4_3 (.CI(n40415), .I0(GND_net), .I1(bit_ctr[1]), 
            .CO(n40416));
    SB_CARRY mod_5_add_1004_3 (.CI(n39719), .I0(n1409), .I1(GND_net), 
            .CO(n39720));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(VCC_net), .O(n1466[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(GND_net), 
            .CO(n39719));
    SB_LUT4 bit_ctr_2058_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(bit_ctr[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_ctr_2058_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21_4_lut_adj_1588 (.I0(bit_ctr[27]), .I1(bit_ctr[31]), .I2(bit_ctr[10]), 
            .I3(bit_ctr[5]), .O(n49));
    defparam i21_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43_adj_4980), .I3(n44_adj_4979), 
            .O(\state_3__N_528[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY bit_ctr_2058_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_ctr[0]), 
            .CO(n40415));
    SB_LUT4 timer_2057_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n40414), .O(n133_adj_5090[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2057_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n40413), .O(n133_adj_5090[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_32 (.CI(n40413), .I0(GND_net), .I1(timer[30]), 
            .CO(n40414));
    SB_LUT4 timer_2057_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n40412), .O(n133_adj_5090[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_31 (.CI(n40412), .I0(GND_net), .I1(timer[29]), 
            .CO(n40413));
    SB_LUT4 timer_2057_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n40411), .O(n133_adj_5090[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_30 (.CI(n40411), .I0(GND_net), .I1(timer[28]), 
            .CO(n40412));
    SB_LUT4 timer_2057_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n40410), .O(n133_adj_5090[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_29 (.CI(n40410), .I0(GND_net), .I1(timer[27]), 
            .CO(n40411));
    SB_LUT4 timer_2057_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n40409), .O(n133_adj_5090[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_28 (.CI(n40409), .I0(GND_net), .I1(timer[26]), 
            .CO(n40410));
    SB_LUT4 i467_2_lut (.I0(LED_c), .I1(\state_3__N_528[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1923));   // verilog/neopixel.v(40[18] 45[12])
    defparam i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 timer_2057_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n40408), .O(n133_adj_5090[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1589 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n27992));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut_adj_1589.LUT_INIT = 16'hbbbb;
    SB_CARRY timer_2057_add_4_27 (.CI(n40408), .I0(GND_net), .I1(timer[25]), 
            .CO(n40409));
    SB_LUT4 timer_2057_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n40407), .O(n133_adj_5090[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_26 (.CI(n40407), .I0(GND_net), .I1(timer[24]), 
            .CO(n40408));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(CLK_c), .E(n29323), .D(state_3__N_528[0]), 
            .S(n29462));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_2057_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n40406), .O(n133_adj_5090[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(n49666), .I1(n6_adj_4990), .I2(n1923), .I3(\state[1] ), 
            .O(n29524));
    defparam i3_4_lut.LUT_INIT = 16'hc040;
    SB_LUT4 i26_4_lut_adj_1590 (.I0(n27992), .I1(n49686), .I2(\state[1] ), 
            .I3(n45055), .O(n6801));
    defparam i26_4_lut_adj_1590.LUT_INIT = 16'hc5c0;
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n29704));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1346_3_lut (.I0(n1900), .I1(n1961[26]), .I2(n1928), 
            .I3(GND_net), .O(n1999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1347_3_lut (.I0(n1901), .I1(n1961[25]), .I2(n1928), 
            .I3(GND_net), .O(n2000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1345_3_lut (.I0(n1899), .I1(n1961[27]), .I2(n1928), 
            .I3(GND_net), .O(n1998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1345_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2057_add_4_25 (.CI(n40406), .I0(GND_net), .I1(timer[23]), 
            .CO(n40407));
    SB_LUT4 mod_5_i1344_3_lut (.I0(n1898), .I1(n1961[28]), .I2(n1928), 
            .I3(GND_net), .O(n1997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1343_3_lut (.I0(n1897), .I1(n1961[29]), .I2(n1928), 
            .I3(GND_net), .O(n1996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1342_3_lut (.I0(n1896), .I1(n1961[30]), .I2(n1928), 
            .I3(GND_net), .O(n1995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1353_3_lut (.I0(n1907), .I1(n1961[19]), .I2(n1928), 
            .I3(GND_net), .O(n2006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1348_3_lut (.I0(n1902), .I1(n1961[24]), .I2(n1928), 
            .I3(GND_net), .O(n2001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1354_3_lut (.I0(n1908), .I1(n1961[18]), .I2(n1928), 
            .I3(GND_net), .O(n2007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1355_3_lut (.I0(n1909), .I1(n1961[17]), .I2(n1928), 
            .I3(GND_net), .O(n2008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1351_3_lut (.I0(n1905), .I1(n1961[21]), .I2(n1928), 
            .I3(GND_net), .O(n2004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1349_3_lut (.I0(n1903), .I1(n1961[23]), .I2(n1928), 
            .I3(GND_net), .O(n2002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2057_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n40405), .O(n133_adj_5090[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_24 (.CI(n40405), .I0(GND_net), .I1(timer[22]), 
            .CO(n40406));
    SB_LUT4 mod_5_i1350_3_lut (.I0(n1904), .I1(n1961[22]), .I2(n1928), 
            .I3(GND_net), .O(n2003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1352_3_lut (.I0(n1906), .I1(n1961[20]), .I2(n1928), 
            .I3(GND_net), .O(n2005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1356_3_lut (.I0(bit_ctr[16]), .I1(n1961[16]), .I2(n1928), 
            .I3(GND_net), .O(n2009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2057_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n40404), .O(n133_adj_5090[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_23 (.CI(n40404), .I0(GND_net), .I1(timer[21]), 
            .CO(n40405));
    SB_LUT4 i22645_2_lut (.I0(bit_ctr[15]), .I1(n2009), .I2(GND_net), 
            .I3(GND_net), .O(n36163));
    defparam i22645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1591 (.I0(n2005), .I1(n2003), .I2(n2002), .I3(n2004), 
            .O(n28_adj_4993));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_2057_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n40403), .O(n133_adj_5090[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1592 (.I0(n1998), .I1(n36163), .I2(n2000), .I3(n1999), 
            .O(n26_adj_4995));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1593 (.I0(n2008), .I1(n2007), .I2(n2001), .I3(n2006), 
            .O(n27_adj_4996));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1995), .I1(n1996), .I2(n1994), .I3(n1997), 
            .O(n25_adj_4997));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1594 (.I0(n25_adj_4997), .I1(n27_adj_4996), .I2(n26_adj_4995), 
            .I3(n28_adj_4993), .O(n2027));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_CARRY timer_2057_add_4_22 (.CI(n40403), .I0(GND_net), .I1(timer[20]), 
            .CO(n40404));
    SB_LUT4 timer_2057_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n40402), .O(n133_adj_5090[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_21 (.CI(n40402), .I0(GND_net), .I1(timer[19]), 
            .CO(n40403));
    SB_LUT4 timer_2057_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n40401), .O(n133_adj_5090[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_20 (.CI(n40401), .I0(GND_net), .I1(timer[18]), 
            .CO(n40402));
    SB_LUT4 timer_2057_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n40400), .O(n133_adj_5090[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_19 (.CI(n40400), .I0(GND_net), .I1(timer[17]), 
            .CO(n40401));
    SB_LUT4 timer_2057_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n40399), .O(n133_adj_5090[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_18 (.CI(n40399), .I0(GND_net), .I1(timer[16]), 
            .CO(n40400));
    SB_LUT4 timer_2057_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n40398), .O(n133_adj_5090[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_17 (.CI(n40398), .I0(GND_net), .I1(timer[15]), 
            .CO(n40399));
    SB_DFFESR bit_ctr_2058__i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n6801), 
            .D(n133[10]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2057_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n40397), .O(n133_adj_5090[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2057_add_4_16 (.CI(n40397), .I0(GND_net), .I1(timer[14]), 
            .CO(n40398));
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_2058__i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n6801), 
            .D(n133[9]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 timer_2057_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n40396), .O(n133_adj_5090[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2057_add_4_15 (.CI(n40396), .I0(GND_net), .I1(timer[13]), 
            .CO(n40397));
    SB_LUT4 timer_2057_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n40395), .O(n133_adj_5090[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_14 (.CI(n40395), .I0(GND_net), .I1(timer[12]), 
            .CO(n40396));
    SB_LUT4 i33423_3_lut (.I0(neopxl_color[8]), .I1(neopxl_color[9]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48860));
    defparam i33423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 timer_2057_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n40394), .O(n133_adj_5090[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33424_3_lut (.I0(neopxl_color[10]), .I1(neopxl_color[11]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48861));
    defparam i33424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33430_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48867));
    defparam i33430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33429_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48866));
    defparam i33429_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY timer_2057_add_4_13 (.CI(n40394), .I0(GND_net), .I1(timer[11]), 
            .CO(n40395));
    SB_LUT4 timer_2057_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n40393), .O(n133_adj_5090[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_12 (.CI(n40393), .I0(GND_net), .I1(timer[10]), 
            .CO(n40394));
    SB_LUT4 timer_2057_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n40392), .O(n133_adj_5090[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_11 (.CI(n40392), .I0(GND_net), .I1(timer[9]), 
            .CO(n40393));
    SB_LUT4 timer_2057_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n40391), .O(n133_adj_5090[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_10 (.CI(n40391), .I0(GND_net), .I1(timer[8]), 
            .CO(n40392));
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2057_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n40390), .O(n133_adj_5090[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_9 (.CI(n40390), .I0(GND_net), .I1(timer[7]), 
            .CO(n40391));
    SB_LUT4 timer_2057_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n40389), .O(n133_adj_5090[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_8 (.CI(n40389), .I0(GND_net), .I1(timer[6]), 
            .CO(n40390));
    SB_LUT4 timer_2057_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n40388), .O(n133_adj_5090[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_7 (.CI(n40388), .I0(GND_net), .I1(timer[5]), 
            .CO(n40389));
    SB_LUT4 timer_2057_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n40387), .O(n133_adj_5090[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_6 (.CI(n40387), .I0(GND_net), .I1(timer[4]), 
            .CO(n40388));
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2057_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n40386), .O(n133_adj_5090[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_5 (.CI(n40386), .I0(GND_net), .I1(timer[3]), 
            .CO(n40387));
    SB_LUT4 timer_2057_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n40385), .O(n133_adj_5090[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_4 (.CI(n40385), .I0(GND_net), .I1(timer[2]), 
            .CO(n40386));
    SB_LUT4 timer_2057_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n40384), .O(n133_adj_5090[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_2057_add_4_3 (.CI(n40384), .I0(GND_net), .I1(timer[1]), 
            .CO(n40385));
    SB_LUT4 timer_2057_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133_adj_5090[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2057_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2057_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n40384));
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1235), .I1(n1202), .I2(VCC_net), 
            .I3(n40376), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'h8228;
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n29703));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1283_3_lut (.I0(n1805), .I1(n1862[22]), .I2(n1829), 
            .I3(GND_net), .O(n1904));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1281_3_lut (.I0(n1803), .I1(n1862[24]), .I2(n1829), 
            .I3(GND_net), .O(n1902));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1285_3_lut (.I0(n1807), .I1(n1862[20]), .I2(n1829), 
            .I3(GND_net), .O(n1906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1288_3_lut (.I0(bit_ctr[17]), .I1(n1862[17]), .I2(n1829), 
            .I3(GND_net), .O(n1909));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1280_3_lut (.I0(n1802), .I1(n1862[25]), .I2(n1829), 
            .I3(GND_net), .O(n1901));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1279_3_lut (.I0(n1801), .I1(n1862[26]), .I2(n1829), 
            .I3(GND_net), .O(n1900));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1277_3_lut (.I0(n1799), .I1(n1862[28]), .I2(n1829), 
            .I3(GND_net), .O(n1898));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1278_3_lut (.I0(n1800), .I1(n1862[27]), .I2(n1829), 
            .I3(GND_net), .O(n1899));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1276_3_lut (.I0(n1798), .I1(n1862[29]), .I2(n1829), 
            .I3(GND_net), .O(n1897));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1275_3_lut (.I0(n1797), .I1(n1862[30]), .I2(n1829), 
            .I3(GND_net), .O(n1896));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1287_3_lut (.I0(n1809), .I1(n1862[18]), .I2(n1829), 
            .I3(GND_net), .O(n1908));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_870_9_lut (.I0(GND_net), .I1(n1203), .I2(VCC_net), 
            .I3(n40375), .O(n1268[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_9 (.CI(n40375), .I0(n1203), .I1(VCC_net), .CO(n40376));
    SB_LUT4 mod_5_add_870_8_lut (.I0(GND_net), .I1(n1204), .I2(VCC_net), 
            .I3(n40374), .O(n1268[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_8 (.CI(n40374), .I0(n1204), .I1(VCC_net), .CO(n40375));
    SB_LUT4 mod_5_i1282_3_lut (.I0(n1804), .I1(n1862[23]), .I2(n1829), 
            .I3(GND_net), .O(n1903));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_870_7_lut (.I0(GND_net), .I1(n1205), .I2(VCC_net), 
            .I3(n40373), .O(n1268[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n29702));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n29701));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n29700));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n29699));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n29698));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n29697));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n29696));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n29695));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n29694));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1286_3_lut (.I0(n1808), .I1(n1862[19]), .I2(n1829), 
            .I3(GND_net), .O(n1907));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1284_3_lut (.I0(n1806), .I1(n1862[21]), .I2(n1829), 
            .I3(GND_net), .O(n1905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1595 (.I0(n1905), .I1(n1907), .I2(n1903), .I3(n1908), 
            .O(n26_adj_5028));
    defparam i11_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(n1901), .I1(bit_ctr[16]), .I2(n1909), .I3(GND_net), 
            .O(n19_adj_5029));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1596 (.I0(n1896), .I1(n1895), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_5030));
    defparam i1_2_lut_adj_1596.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1597 (.I0(n1897), .I1(n1899), .I2(n1898), .I3(n1900), 
            .O(n24_adj_5031));
    defparam i9_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1598 (.I0(n19_adj_5029), .I1(n26_adj_5028), .I2(n1902), 
            .I3(n1904), .O(n28_adj_5032));
    defparam i13_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1599 (.I0(n1906), .I1(n28_adj_5032), .I2(n24_adj_5031), 
            .I3(n16_adj_5030), .O(n1928));
    defparam i14_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_870_7 (.CI(n40373), .I0(n1205), .I1(VCC_net), .CO(n40374));
    SB_LUT4 mod_5_add_870_6_lut (.I0(GND_net), .I1(n1206), .I2(VCC_net), 
            .I3(n40372), .O(n1268[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_6 (.CI(n40372), .I0(n1206), .I1(VCC_net), .CO(n40373));
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_870_5_lut (.I0(GND_net), .I1(n1207), .I2(VCC_net), 
            .I3(n40371), .O(n1268[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_5 (.CI(n40371), .I0(n1207), .I1(VCC_net), .CO(n40372));
    SB_LUT4 mod_5_add_870_4_lut (.I0(GND_net), .I1(n1208), .I2(VCC_net), 
            .I3(n40370), .O(n1268[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_4 (.CI(n40370), .I0(n1208), .I1(VCC_net), .CO(n40371));
    SB_LUT4 mod_5_add_870_3_lut (.I0(GND_net), .I1(n1209), .I2(GND_net), 
            .I3(n40369), .O(n1268[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_3 (.CI(n40369), .I0(n1209), .I1(GND_net), .CO(n40370));
    SB_LUT4 mod_5_add_870_2_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(VCC_net), .O(n1268[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(GND_net), 
            .CO(n40369));
    SB_DFF timer_2057__i0 (.Q(timer[0]), .C(CLK_c), .D(n133_adj_5090[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_736_8_lut (.I0(n50683), .I1(n50683), .I2(n1037), 
            .I3(n40920), .O(n8_adj_4935)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n50665), .I1(n50665), .I2(n1037), 
            .I3(n40919), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n40919), .I0(n50665), .I1(n1037), .CO(n40920));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n50661), .I1(n1006), .I2(n1037), 
            .I3(n40918), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n40918), .I0(n1006), .I1(n1037), .CO(n40919));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n50662), .I1(n1007), .I2(n1037), 
            .I3(n40917), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n40917), .I0(n1007), .I1(n1037), .CO(n40918));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n40916), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n40916), .I0(n1008), .I1(n1037), .CO(n40917));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n51353), 
            .I3(n40915), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n40915), .I0(n1009), .I1(n51353), .CO(n40916));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n51353), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n51353), 
            .CO(n40915));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1136), .I1(n8_adj_4935), .I2(VCC_net), 
            .I3(n40909), .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_803_8_lut (.I0(GND_net), .I1(n1104), .I2(VCC_net), 
            .I3(n40908), .O(n1169[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_8 (.CI(n40908), .I0(n1104), .I1(VCC_net), .CO(n40909));
    SB_LUT4 mod_5_add_803_7_lut (.I0(GND_net), .I1(n1105), .I2(VCC_net), 
            .I3(n40907), .O(n1169[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_7 (.CI(n40907), .I0(n1105), .I1(VCC_net), .CO(n40908));
    SB_LUT4 mod_5_add_803_6_lut (.I0(GND_net), .I1(n1106), .I2(VCC_net), 
            .I3(n40906), .O(n1169[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_6 (.CI(n40906), .I0(n1106), .I1(VCC_net), .CO(n40907));
    SB_LUT4 mod_5_add_803_5_lut (.I0(GND_net), .I1(n1107), .I2(VCC_net), 
            .I3(n40905), .O(n1169[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_5 (.CI(n40905), .I0(n1107), .I1(VCC_net), .CO(n40906));
    SB_LUT4 mod_5_add_803_4_lut (.I0(GND_net), .I1(n1108), .I2(VCC_net), 
            .I3(n40904), .O(n1169[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_4 (.CI(n40904), .I0(n1108), .I1(VCC_net), .CO(n40905));
    SB_LUT4 mod_5_add_803_3_lut (.I0(GND_net), .I1(n1109), .I2(GND_net), 
            .I3(n40903), .O(n1169[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_3 (.CI(n40903), .I0(n1109), .I1(GND_net), .CO(n40904));
    SB_LUT4 mod_5_add_803_2_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(VCC_net), .O(n1169[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(GND_net), 
            .CO(n40903));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n40902), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n40901), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_13 (.CI(n40901), .I0(n1599), .I1(n1631), .CO(n40902));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n40900), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n40900), .I0(n1600), .I1(n1631), .CO(n40901));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n40899), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n40899), .I0(n1601), .I1(n1631), .CO(n40900));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n40898), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1138_10 (.CI(n40898), .I0(n1602), .I1(n1631), .CO(n40899));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n40897), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n40897), .I0(n1603), .I1(n1631), .CO(n40898));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n40896), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n40896), .I0(n1604), .I1(n1631), .CO(n40897));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n40895), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n40895), .I0(n1605), .I1(n1631), .CO(n40896));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n40894), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n40894), .I0(n1606), .I1(n1631), .CO(n40895));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n40893), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n40893), .I0(n1607), .I1(n1631), .CO(n40894));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n40892), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n40892), .I0(n1608), .I1(n1631), .CO(n40893));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n51354), 
            .I3(n40891), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n40891), .I0(n1609), .I1(n51354), .CO(n40892));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n51354), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n51354), 
            .CO(n40891));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1730), .I1(n1697), .I2(VCC_net), 
            .I3(n40890), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(GND_net), .I1(n1698), .I2(VCC_net), 
            .I3(n40889), .O(n1763[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_14 (.CI(n40889), .I0(n1698), .I1(VCC_net), 
            .CO(n40890));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(GND_net), .I1(n1699), .I2(VCC_net), 
            .I3(n40888), .O(n1763[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_13 (.CI(n40888), .I0(n1699), .I1(VCC_net), 
            .CO(n40889));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(GND_net), .I1(n1700), .I2(VCC_net), 
            .I3(n40887), .O(n1763[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_12 (.CI(n40887), .I0(n1700), .I1(VCC_net), 
            .CO(n40888));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(GND_net), .I1(n1701), .I2(VCC_net), 
            .I3(n40886), .O(n1763[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_11 (.CI(n40886), .I0(n1701), .I1(VCC_net), 
            .CO(n40887));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(GND_net), .I1(n1702), .I2(VCC_net), 
            .I3(n40885), .O(n1763[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_10 (.CI(n40885), .I0(n1702), .I1(VCC_net), 
            .CO(n40886));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(GND_net), .I1(n1703), .I2(VCC_net), 
            .I3(n40884), .O(n1763[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_9 (.CI(n40884), .I0(n1703), .I1(VCC_net), 
            .CO(n40885));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(GND_net), .I1(n1704), .I2(VCC_net), 
            .I3(n40883), .O(n1763[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_8 (.CI(n40883), .I0(n1704), .I1(VCC_net), 
            .CO(n40884));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(GND_net), .I1(n1705), .I2(VCC_net), 
            .I3(n40882), .O(n1763[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_7 (.CI(n40882), .I0(n1705), .I1(VCC_net), 
            .CO(n40883));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(GND_net), .I1(n1706), .I2(VCC_net), 
            .I3(n40881), .O(n1763[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_6 (.CI(n40881), .I0(n1706), .I1(VCC_net), 
            .CO(n40882));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(GND_net), .I1(n1707), .I2(VCC_net), 
            .I3(n40880), .O(n1763[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_5 (.CI(n40880), .I0(n1707), .I1(VCC_net), 
            .CO(n40881));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(GND_net), .I1(n1708), .I2(VCC_net), 
            .I3(n40879), .O(n1763[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_4 (.CI(n40879), .I0(n1708), .I1(VCC_net), 
            .CO(n40880));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(GND_net), .I1(n1709), .I2(GND_net), 
            .I3(n40878), .O(n1763[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_3 (.CI(n40878), .I0(n1709), .I1(GND_net), 
            .CO(n40879));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(VCC_net), .O(n1763[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(GND_net), 
            .CO(n40878));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1829), .I1(n1796), .I2(VCC_net), 
            .I3(n40877), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(GND_net), .I1(n1797), .I2(VCC_net), 
            .I3(n40876), .O(n1862[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_15 (.CI(n40876), .I0(n1797), .I1(VCC_net), 
            .CO(n40877));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(GND_net), .I1(n1798), .I2(VCC_net), 
            .I3(n40875), .O(n1862[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_14 (.CI(n40875), .I0(n1798), .I1(VCC_net), 
            .CO(n40876));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(GND_net), .I1(n1799), .I2(VCC_net), 
            .I3(n40874), .O(n1862[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_13 (.CI(n40874), .I0(n1799), .I1(VCC_net), 
            .CO(n40875));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(GND_net), .I1(n1800), .I2(VCC_net), 
            .I3(n40873), .O(n1862[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_12 (.CI(n40873), .I0(n1800), .I1(VCC_net), 
            .CO(n40874));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(GND_net), .I1(n1801), .I2(VCC_net), 
            .I3(n40872), .O(n1862[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_11 (.CI(n40872), .I0(n1801), .I1(VCC_net), 
            .CO(n40873));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(GND_net), .I1(n1802), .I2(VCC_net), 
            .I3(n40871), .O(n1862[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_10 (.CI(n40871), .I0(n1802), .I1(VCC_net), 
            .CO(n40872));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(GND_net), .I1(n1803), .I2(VCC_net), 
            .I3(n40870), .O(n1862[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_9 (.CI(n40870), .I0(n1803), .I1(VCC_net), 
            .CO(n40871));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(GND_net), .I1(n1804), .I2(VCC_net), 
            .I3(n40869), .O(n1862[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_8 (.CI(n40869), .I0(n1804), .I1(VCC_net), 
            .CO(n40870));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(GND_net), .I1(n1805), .I2(VCC_net), 
            .I3(n40868), .O(n1862[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_7 (.CI(n40868), .I0(n1805), .I1(VCC_net), 
            .CO(n40869));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(GND_net), .I1(n1806), .I2(VCC_net), 
            .I3(n40867), .O(n1862[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_6 (.CI(n40867), .I0(n1806), .I1(VCC_net), 
            .CO(n40868));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(GND_net), .I1(n1807), .I2(VCC_net), 
            .I3(n40866), .O(n1862[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_5 (.CI(n40866), .I0(n1807), .I1(VCC_net), 
            .CO(n40867));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(GND_net), .I1(n1808), .I2(VCC_net), 
            .I3(n40865), .O(n1862[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_4 (.CI(n40865), .I0(n1808), .I1(VCC_net), 
            .CO(n40866));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(GND_net), .I1(n1809), .I2(GND_net), 
            .I3(n40864), .O(n1862[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_3 (.CI(n40864), .I0(n1809), .I1(GND_net), 
            .CO(n40865));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(VCC_net), .O(n1862[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(GND_net), 
            .CO(n40864));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1928), .I1(n1895), .I2(VCC_net), 
            .I3(n40863), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(GND_net), .I1(n1896), .I2(VCC_net), 
            .I3(n40862), .O(n1961[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_16 (.CI(n40862), .I0(n1896), .I1(VCC_net), 
            .CO(n40863));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(GND_net), .I1(n1897), .I2(VCC_net), 
            .I3(n40861), .O(n1961[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_15 (.CI(n40861), .I0(n1897), .I1(VCC_net), 
            .CO(n40862));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(GND_net), .I1(n1898), .I2(VCC_net), 
            .I3(n40860), .O(n1961[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_14 (.CI(n40860), .I0(n1898), .I1(VCC_net), 
            .CO(n40861));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(GND_net), .I1(n1899), .I2(VCC_net), 
            .I3(n40859), .O(n1961[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_13 (.CI(n40859), .I0(n1899), .I1(VCC_net), 
            .CO(n40860));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(GND_net), .I1(n1900), .I2(VCC_net), 
            .I3(n40858), .O(n1961[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_12 (.CI(n40858), .I0(n1900), .I1(VCC_net), 
            .CO(n40859));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(GND_net), .I1(n1901), .I2(VCC_net), 
            .I3(n40857), .O(n1961[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_11 (.CI(n40857), .I0(n1901), .I1(VCC_net), 
            .CO(n40858));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(GND_net), .I1(n1902), .I2(VCC_net), 
            .I3(n40856), .O(n1961[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_10 (.CI(n40856), .I0(n1902), .I1(VCC_net), 
            .CO(n40857));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(GND_net), .I1(n1903), .I2(VCC_net), 
            .I3(n40855), .O(n1961[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_9 (.CI(n40855), .I0(n1903), .I1(VCC_net), 
            .CO(n40856));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(GND_net), .I1(n1904), .I2(VCC_net), 
            .I3(n40854), .O(n1961[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_8 (.CI(n40854), .I0(n1904), .I1(VCC_net), 
            .CO(n40855));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(GND_net), .I1(n1905), .I2(VCC_net), 
            .I3(n40853), .O(n1961[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_7 (.CI(n40853), .I0(n1905), .I1(VCC_net), 
            .CO(n40854));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(GND_net), .I1(n1906), .I2(VCC_net), 
            .I3(n40852), .O(n1961[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_6 (.CI(n40852), .I0(n1906), .I1(VCC_net), 
            .CO(n40853));
    SB_DFFESR bit_ctr_2058__i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n6801), 
            .D(n133[8]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_add_1339_5_lut (.I0(GND_net), .I1(n1907), .I2(VCC_net), 
            .I3(n40851), .O(n1961[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_5 (.CI(n40851), .I0(n1907), .I1(VCC_net), 
            .CO(n40852));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(GND_net), .I1(n1908), .I2(VCC_net), 
            .I3(n40850), .O(n1961[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_4 (.CI(n40850), .I0(n1908), .I1(VCC_net), 
            .CO(n40851));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(GND_net), .I1(n1909), .I2(GND_net), 
            .I3(n40849), .O(n1961[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_3 (.CI(n40849), .I0(n1909), .I1(GND_net), 
            .CO(n40850));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(VCC_net), .O(n1961[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(GND_net), 
            .CO(n40849));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n2027), .I1(n1994), .I2(VCC_net), 
            .I3(n40848), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(GND_net), .I1(n1995), .I2(VCC_net), 
            .I3(n40847), .O(n2060[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_17 (.CI(n40847), .I0(n1995), .I1(VCC_net), 
            .CO(n40848));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(GND_net), .I1(n1996), .I2(VCC_net), 
            .I3(n40846), .O(n2060[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_16 (.CI(n40846), .I0(n1996), .I1(VCC_net), 
            .CO(n40847));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(GND_net), .I1(n1997), .I2(VCC_net), 
            .I3(n40845), .O(n2060[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_15 (.CI(n40845), .I0(n1997), .I1(VCC_net), 
            .CO(n40846));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(GND_net), .I1(n1998), .I2(VCC_net), 
            .I3(n40844), .O(n2060[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_14 (.CI(n40844), .I0(n1998), .I1(VCC_net), 
            .CO(n40845));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(GND_net), .I1(n1999), .I2(VCC_net), 
            .I3(n40843), .O(n2060[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_13 (.CI(n40843), .I0(n1999), .I1(VCC_net), 
            .CO(n40844));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(GND_net), .I1(n2000), .I2(VCC_net), 
            .I3(n40842), .O(n2060[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_12 (.CI(n40842), .I0(n2000), .I1(VCC_net), 
            .CO(n40843));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(GND_net), .I1(n2001), .I2(VCC_net), 
            .I3(n40841), .O(n2060[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_11 (.CI(n40841), .I0(n2001), .I1(VCC_net), 
            .CO(n40842));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(GND_net), .I1(n2002), .I2(VCC_net), 
            .I3(n40840), .O(n2060[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_10 (.CI(n40840), .I0(n2002), .I1(VCC_net), 
            .CO(n40841));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(GND_net), .I1(n2003), .I2(VCC_net), 
            .I3(n40839), .O(n2060[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_9 (.CI(n40839), .I0(n2003), .I1(VCC_net), 
            .CO(n40840));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(GND_net), .I1(n2004), .I2(VCC_net), 
            .I3(n40838), .O(n2060[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_33_lut (.I0(n48490), .I1(timer[31]), .I2(n1[31]), 
            .I3(n39279), .O(n27999)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n48488), .I1(timer[30]), .I2(n1[30]), 
            .I3(n39278), .O(n48490)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1406_8 (.CI(n40838), .I0(n2004), .I1(VCC_net), 
            .CO(n40839));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(GND_net), .I1(n2005), .I2(VCC_net), 
            .I3(n40837), .O(n2060[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_7 (.CI(n40837), .I0(n2005), .I1(VCC_net), 
            .CO(n40838));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(GND_net), .I1(n2006), .I2(VCC_net), 
            .I3(n40836), .O(n2060[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_6 (.CI(n40836), .I0(n2006), .I1(VCC_net), 
            .CO(n40837));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(GND_net), .I1(n2007), .I2(VCC_net), 
            .I3(n40835), .O(n2060[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_5 (.CI(n40835), .I0(n2007), .I1(VCC_net), 
            .CO(n40836));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(GND_net), .I1(n2008), .I2(VCC_net), 
            .I3(n40834), .O(n2060[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_4 (.CI(n40834), .I0(n2008), .I1(VCC_net), 
            .CO(n40835));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(GND_net), .I1(n2009), .I2(GND_net), 
            .I3(n40833), .O(n2060[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_3 (.CI(n40833), .I0(n2009), .I1(GND_net), 
            .CO(n40834));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(VCC_net), .O(n2060[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(GND_net), 
            .CO(n40833));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2126), .I1(n2093), .I2(VCC_net), 
            .I3(n40832), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(GND_net), .I1(n2094), .I2(VCC_net), 
            .I3(n40831), .O(n2159[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_18 (.CI(n40831), .I0(n2094), .I1(VCC_net), 
            .CO(n40832));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(GND_net), .I1(n2095), .I2(VCC_net), 
            .I3(n40830), .O(n2159[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_17 (.CI(n40830), .I0(n2095), .I1(VCC_net), 
            .CO(n40831));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(GND_net), .I1(n2096), .I2(VCC_net), 
            .I3(n40829), .O(n2159[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_16 (.CI(n40829), .I0(n2096), .I1(VCC_net), 
            .CO(n40830));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(GND_net), .I1(n2097), .I2(VCC_net), 
            .I3(n40828), .O(n2159[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_15 (.CI(n40828), .I0(n2097), .I1(VCC_net), 
            .CO(n40829));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(GND_net), .I1(n2098), .I2(VCC_net), 
            .I3(n40827), .O(n2159[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_14 (.CI(n40827), .I0(n2098), .I1(VCC_net), 
            .CO(n40828));
    SB_CARRY sub_14_add_2_32 (.CI(n39278), .I0(timer[30]), .I1(n1[30]), 
            .CO(n39279));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(GND_net), .I1(n2099), .I2(VCC_net), 
            .I3(n40826), .O(n2159[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_13 (.CI(n40826), .I0(n2099), .I1(VCC_net), 
            .CO(n40827));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(GND_net), .I1(n2100), .I2(VCC_net), 
            .I3(n40825), .O(n2159[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_12 (.CI(n40825), .I0(n2100), .I1(VCC_net), 
            .CO(n40826));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(GND_net), .I1(n2101), .I2(VCC_net), 
            .I3(n40824), .O(n2159[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_11 (.CI(n40824), .I0(n2101), .I1(VCC_net), 
            .CO(n40825));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(GND_net), .I1(n2102), .I2(VCC_net), 
            .I3(n40823), .O(n2159[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_10 (.CI(n40823), .I0(n2102), .I1(VCC_net), 
            .CO(n40824));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(GND_net), .I1(n2103), .I2(VCC_net), 
            .I3(n40822), .O(n2159[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_31_lut (.I0(n48486), .I1(timer[29]), .I2(n1[29]), 
            .I3(n39277), .O(n48488)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1473_9 (.CI(n40822), .I0(n2103), .I1(VCC_net), 
            .CO(n40823));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(GND_net), .I1(n2104), .I2(VCC_net), 
            .I3(n40821), .O(n2159[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_8 (.CI(n40821), .I0(n2104), .I1(VCC_net), 
            .CO(n40822));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(GND_net), .I1(n2105), .I2(VCC_net), 
            .I3(n40820), .O(n2159[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_7 (.CI(n40820), .I0(n2105), .I1(VCC_net), 
            .CO(n40821));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(GND_net), .I1(n2106), .I2(VCC_net), 
            .I3(n40819), .O(n2159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_6 (.CI(n40819), .I0(n2106), .I1(VCC_net), 
            .CO(n40820));
    SB_CARRY sub_14_add_2_31 (.CI(n39277), .I0(timer[29]), .I1(n1[29]), 
            .CO(n39278));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n48484), .I1(timer[28]), .I2(n1[28]), 
            .I3(n39276), .O(n48486)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1473_5_lut (.I0(GND_net), .I1(n2107), .I2(VCC_net), 
            .I3(n40818), .O(n2159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1215_3_lut (.I0(n1705), .I1(n1763[23]), .I2(n1730), 
            .I3(GND_net), .O(n1804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1211_3_lut (.I0(n1701), .I1(n1763[27]), .I2(n1730), 
            .I3(GND_net), .O(n1800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1210_3_lut (.I0(n1700), .I1(n1763[28]), .I2(n1730), 
            .I3(GND_net), .O(n1799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1209_3_lut (.I0(n1699), .I1(n1763[29]), .I2(n1730), 
            .I3(GND_net), .O(n1798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1209_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_30 (.CI(n39276), .I0(timer[28]), .I1(n1[28]), 
            .CO(n39277));
    SB_LUT4 sub_14_add_2_29_lut (.I0(n48482), .I1(timer[27]), .I2(n1[27]), 
            .I3(n39275), .O(n48484)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_i1208_3_lut (.I0(n1698), .I1(n1763[30]), .I2(n1730), 
            .I3(GND_net), .O(n1797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1208_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_29 (.CI(n39275), .I0(timer[27]), .I1(n1[27]), 
            .CO(n39276));
    SB_LUT4 mod_5_i1216_3_lut (.I0(n1706), .I1(n1763[22]), .I2(n1730), 
            .I3(GND_net), .O(n1805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1213_3_lut (.I0(n1703), .I1(n1763[25]), .I2(n1730), 
            .I3(GND_net), .O(n1802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1219_3_lut (.I0(n1709), .I1(n1763[19]), .I2(n1730), 
            .I3(GND_net), .O(n1808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1218_3_lut (.I0(n1708), .I1(n1763[20]), .I2(n1730), 
            .I3(GND_net), .O(n1807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1214_3_lut (.I0(n1704), .I1(n1763[24]), .I2(n1730), 
            .I3(GND_net), .O(n1803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1212_3_lut (.I0(n1702), .I1(n1763[26]), .I2(n1730), 
            .I3(GND_net), .O(n1801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1220_3_lut (.I0(bit_ctr[18]), .I1(n1763[18]), .I2(n1730), 
            .I3(GND_net), .O(n1809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1217_3_lut (.I0(n1707), .I1(n1763[21]), .I2(n1730), 
            .I3(GND_net), .O(n1806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_3_lut_adj_1600 (.I0(bit_ctr[17]), .I1(n1806), .I2(n1809), 
            .I3(GND_net), .O(n18_adj_5034));   // verilog/neopixel.v(22[26:36])
    defparam i4_3_lut_adj_1600.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1601 (.I0(n1801), .I1(n1803), .I2(n1807), .I3(n1808), 
            .O(n24_adj_5035));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1602 (.I0(n1797), .I1(n1798), .I2(n1796), .I3(n1799), 
            .O(n22_adj_5036));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1603 (.I0(n1800), .I1(n24_adj_5035), .I2(n18_adj_5034), 
            .I3(n1804), .O(n26_adj_5037));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1604 (.I0(n1802), .I1(n26_adj_5037), .I2(n22_adj_5036), 
            .I3(n1805), .O(n1829));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_28_lut (.I0(n48480), .I1(timer[26]), .I2(n1[26]), 
            .I3(n39274), .O(n48482)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1473_5 (.CI(n40818), .I0(n2107), .I1(VCC_net), 
            .CO(n40819));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(GND_net), .I1(n2108), .I2(VCC_net), 
            .I3(n40817), .O(n2159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_4 (.CI(n40817), .I0(n2108), .I1(VCC_net), 
            .CO(n40818));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(GND_net), .I1(n2109), .I2(GND_net), 
            .I3(n40816), .O(n2159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_3 (.CI(n40816), .I0(n2109), .I1(GND_net), 
            .CO(n40817));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(VCC_net), .O(n2159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(GND_net), 
            .CO(n40816));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2225), .I1(n2192), .I2(VCC_net), 
            .I3(n40815), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(GND_net), .I1(n2193), .I2(VCC_net), 
            .I3(n40814), .O(n2258[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_19 (.CI(n40814), .I0(n2193), .I1(VCC_net), 
            .CO(n40815));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(GND_net), .I1(n2194), .I2(VCC_net), 
            .I3(n40813), .O(n2258[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_18 (.CI(n40813), .I0(n2194), .I1(VCC_net), 
            .CO(n40814));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(GND_net), .I1(n2195), .I2(VCC_net), 
            .I3(n40812), .O(n2258[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_17 (.CI(n40812), .I0(n2195), .I1(VCC_net), 
            .CO(n40813));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(GND_net), .I1(n2196), .I2(VCC_net), 
            .I3(n40811), .O(n2258[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_16 (.CI(n40811), .I0(n2196), .I1(VCC_net), 
            .CO(n40812));
    SB_LUT4 i4_3_lut_adj_1605 (.I0(bit_ctr[18]), .I1(n1703), .I2(n1709), 
            .I3(GND_net), .O(n17_adj_5038));   // verilog/neopixel.v(22[26:36])
    defparam i4_3_lut_adj_1605.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1540_15_lut (.I0(GND_net), .I1(n2197), .I2(VCC_net), 
            .I3(n40810), .O(n2258[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut_adj_1606 (.I0(n1699), .I1(n1701), .I2(n1700), .I3(n1702), 
            .O(n21_adj_5039));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1607 (.I0(n1705), .I1(n1698), .I2(n1697), .I3(GND_net), 
            .O(n20));   // verilog/neopixel.v(22[26:36])
    defparam i7_3_lut_adj_1607.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_1540_15 (.CI(n40810), .I0(n2197), .I1(VCC_net), 
            .CO(n40811));
    SB_LUT4 i11_4_lut_adj_1608 (.I0(n21_adj_5039), .I1(n17_adj_5038), .I2(n1706), 
            .I3(n1707), .O(n24_adj_5040));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(GND_net), .I1(n2198), .I2(VCC_net), 
            .I3(n40809), .O(n2258[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_14 (.CI(n40809), .I0(n2198), .I1(VCC_net), 
            .CO(n40810));
    SB_LUT4 i12_4_lut_adj_1609 (.I0(n1708), .I1(n24_adj_5040), .I2(n20), 
            .I3(n1704), .O(n1730));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_13_lut (.I0(GND_net), .I1(n2199), .I2(VCC_net), 
            .I3(n40808), .O(n2258[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_13 (.CI(n40808), .I0(n2199), .I1(VCC_net), 
            .CO(n40809));
    SB_LUT4 i35916_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51354));
    defparam i35916_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_12_lut (.I0(GND_net), .I1(n2200), .I2(VCC_net), 
            .I3(n40807), .O(n2258[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_12 (.CI(n40807), .I0(n2200), .I1(VCC_net), 
            .CO(n40808));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(GND_net), .I1(n2201), .I2(VCC_net), 
            .I3(n40806), .O(n2258[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_28 (.CI(n39274), .I0(timer[26]), .I1(n1[26]), 
            .CO(n39275));
    SB_CARRY mod_5_add_1540_11 (.CI(n40806), .I0(n2201), .I1(VCC_net), 
            .CO(n40807));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(GND_net), .I1(n2202), .I2(VCC_net), 
            .I3(n40805), .O(n2258[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_10 (.CI(n40805), .I0(n2202), .I1(VCC_net), 
            .CO(n40806));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(GND_net), .I1(n2203), .I2(VCC_net), 
            .I3(n40804), .O(n2258[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_9 (.CI(n40804), .I0(n2203), .I1(VCC_net), 
            .CO(n40805));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(GND_net), .I1(n2204), .I2(VCC_net), 
            .I3(n40803), .O(n2258[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_8 (.CI(n40803), .I0(n2204), .I1(VCC_net), 
            .CO(n40804));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(GND_net), .I1(n2205), .I2(VCC_net), 
            .I3(n40802), .O(n2258[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_7 (.CI(n40802), .I0(n2205), .I1(VCC_net), 
            .CO(n40803));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(GND_net), .I1(n2206), .I2(VCC_net), 
            .I3(n40801), .O(n2258[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_6 (.CI(n40801), .I0(n2206), .I1(VCC_net), 
            .CO(n40802));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(GND_net), .I1(n2207), .I2(VCC_net), 
            .I3(n40800), .O(n2258[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_5 (.CI(n40800), .I0(n2207), .I1(VCC_net), 
            .CO(n40801));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(GND_net), .I1(n2208), .I2(VCC_net), 
            .I3(n40799), .O(n2258[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_4 (.CI(n40799), .I0(n2208), .I1(VCC_net), 
            .CO(n40800));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(GND_net), .I1(n2209), .I2(GND_net), 
            .I3(n40798), .O(n2258[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_3 (.CI(n40798), .I0(n2209), .I1(GND_net), 
            .CO(n40799));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(VCC_net), .O(n2258[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(GND_net), 
            .CO(n40798));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2324), .I1(n2291), .I2(VCC_net), 
            .I3(n40797), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(GND_net), .I1(n2292), .I2(VCC_net), 
            .I3(n40796), .O(n2357[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_27_lut (.I0(n48478), .I1(timer[25]), .I2(n1[25]), 
            .I3(n39273), .O(n48480)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1607_20 (.CI(n40796), .I0(n2292), .I1(VCC_net), 
            .CO(n40797));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(GND_net), .I1(n2293), .I2(VCC_net), 
            .I3(n40795), .O(n2357[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_19 (.CI(n40795), .I0(n2293), .I1(VCC_net), 
            .CO(n40796));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(GND_net), .I1(n2294), .I2(VCC_net), 
            .I3(n40794), .O(n2357[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_18 (.CI(n40794), .I0(n2294), .I1(VCC_net), 
            .CO(n40795));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(GND_net), .I1(n2295), .I2(VCC_net), 
            .I3(n40793), .O(n2357[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_27 (.CI(n39273), .I0(timer[25]), .I1(n1[25]), 
            .CO(n39274));
    SB_CARRY mod_5_add_1607_17 (.CI(n40793), .I0(n2295), .I1(VCC_net), 
            .CO(n40794));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(GND_net), .I1(n2296), .I2(VCC_net), 
            .I3(n40792), .O(n2357[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_16 (.CI(n40792), .I0(n2296), .I1(VCC_net), 
            .CO(n40793));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(GND_net), .I1(n2297), .I2(VCC_net), 
            .I3(n40791), .O(n2357[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_15 (.CI(n40791), .I0(n2297), .I1(VCC_net), 
            .CO(n40792));
    SB_LUT4 sub_14_add_2_26_lut (.I0(n48476), .I1(timer[24]), .I2(n1[24]), 
            .I3(n39272), .O(n48478)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1607_14_lut (.I0(GND_net), .I1(n2298), .I2(VCC_net), 
            .I3(n40790), .O(n2357[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_14 (.CI(n40790), .I0(n2298), .I1(VCC_net), 
            .CO(n40791));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(GND_net), .I1(n2299), .I2(VCC_net), 
            .I3(n40789), .O(n2357[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_13 (.CI(n40789), .I0(n2299), .I1(VCC_net), 
            .CO(n40790));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(GND_net), .I1(n2300), .I2(VCC_net), 
            .I3(n40788), .O(n2357[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_12 (.CI(n40788), .I0(n2300), .I1(VCC_net), 
            .CO(n40789));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(GND_net), .I1(n2301), .I2(VCC_net), 
            .I3(n40787), .O(n2357[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_11 (.CI(n40787), .I0(n2301), .I1(VCC_net), 
            .CO(n40788));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(GND_net), .I1(n2302), .I2(VCC_net), 
            .I3(n40786), .O(n2357[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n40786), .I0(n2302), .I1(VCC_net), 
            .CO(n40787));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(GND_net), .I1(n2303), .I2(VCC_net), 
            .I3(n40785), .O(n2357[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_9 (.CI(n40785), .I0(n2303), .I1(VCC_net), 
            .CO(n40786));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(GND_net), .I1(n2304), .I2(VCC_net), 
            .I3(n40784), .O(n2357[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_8 (.CI(n40784), .I0(n2304), .I1(VCC_net), 
            .CO(n40785));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(GND_net), .I1(n2305), .I2(VCC_net), 
            .I3(n40783), .O(n2357[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_7 (.CI(n40783), .I0(n2305), .I1(VCC_net), 
            .CO(n40784));
    SB_CARRY sub_14_add_2_26 (.CI(n39272), .I0(timer[24]), .I1(n1[24]), 
            .CO(n39273));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(GND_net), .I1(n2306), .I2(VCC_net), 
            .I3(n40782), .O(n2357[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_6 (.CI(n40782), .I0(n2306), .I1(VCC_net), 
            .CO(n40783));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(GND_net), .I1(n2307), .I2(VCC_net), 
            .I3(n40781), .O(n2357[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_5 (.CI(n40781), .I0(n2307), .I1(VCC_net), 
            .CO(n40782));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(GND_net), .I1(n2308), .I2(VCC_net), 
            .I3(n40780), .O(n2357[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_4 (.CI(n40780), .I0(n2308), .I1(VCC_net), 
            .CO(n40781));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(GND_net), .I1(n2309), .I2(GND_net), 
            .I3(n40779), .O(n2357[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_3 (.CI(n40779), .I0(n2309), .I1(GND_net), 
            .CO(n40780));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(VCC_net), .O(n2357[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(GND_net), 
            .CO(n40779));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2423), .I1(n2390), .I2(VCC_net), 
            .I3(n40778), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(GND_net), .I1(n2391), .I2(VCC_net), 
            .I3(n40777), .O(n2456[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_21 (.CI(n40777), .I0(n2391), .I1(VCC_net), 
            .CO(n40778));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(GND_net), .I1(n2392), .I2(VCC_net), 
            .I3(n40776), .O(n2456[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_20 (.CI(n40776), .I0(n2392), .I1(VCC_net), 
            .CO(n40777));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(GND_net), .I1(n2393), .I2(VCC_net), 
            .I3(n40775), .O(n2456[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_19 (.CI(n40775), .I0(n2393), .I1(VCC_net), 
            .CO(n40776));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(GND_net), .I1(n2394), .I2(VCC_net), 
            .I3(n40774), .O(n2456[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_18 (.CI(n40774), .I0(n2394), .I1(VCC_net), 
            .CO(n40775));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(GND_net), .I1(n2395), .I2(VCC_net), 
            .I3(n40773), .O(n2456[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_17 (.CI(n40773), .I0(n2395), .I1(VCC_net), 
            .CO(n40774));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(GND_net), .I1(n2396), .I2(VCC_net), 
            .I3(n40772), .O(n2456[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_16 (.CI(n40772), .I0(n2396), .I1(VCC_net), 
            .CO(n40773));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(GND_net), .I1(n2397), .I2(VCC_net), 
            .I3(n40771), .O(n2456[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_15 (.CI(n40771), .I0(n2397), .I1(VCC_net), 
            .CO(n40772));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(GND_net), .I1(n2398), .I2(VCC_net), 
            .I3(n40770), .O(n2456[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_14 (.CI(n40770), .I0(n2398), .I1(VCC_net), 
            .CO(n40771));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(GND_net), .I1(n2399), .I2(VCC_net), 
            .I3(n40769), .O(n2456[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_25_lut (.I0(n48474), .I1(timer[23]), .I2(n1[23]), 
            .I3(n39271), .O(n48476)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1674_13 (.CI(n40769), .I0(n2399), .I1(VCC_net), 
            .CO(n40770));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(GND_net), .I1(n2400), .I2(VCC_net), 
            .I3(n40768), .O(n2456[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_12 (.CI(n40768), .I0(n2400), .I1(VCC_net), 
            .CO(n40769));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(GND_net), .I1(n2401), .I2(VCC_net), 
            .I3(n40767), .O(n2456[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_11 (.CI(n40767), .I0(n2401), .I1(VCC_net), 
            .CO(n40768));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(GND_net), .I1(n2402), .I2(VCC_net), 
            .I3(n40766), .O(n2456[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_10 (.CI(n40766), .I0(n2402), .I1(VCC_net), 
            .CO(n40767));
    SB_CARRY sub_14_add_2_25 (.CI(n39271), .I0(timer[23]), .I1(n1[23]), 
            .CO(n39272));
    SB_LUT4 i15935_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n29323), 
            .I3(GND_net), .O(n29462));
    defparam i15935_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 mod_5_add_1674_9_lut (.I0(GND_net), .I1(n2403), .I2(VCC_net), 
            .I3(n40765), .O(n2456[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n40765), .I0(n2403), .I1(VCC_net), 
            .CO(n40766));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(GND_net), .I1(n2404), .I2(VCC_net), 
            .I3(n40764), .O(n2456[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_8 (.CI(n40764), .I0(n2404), .I1(VCC_net), 
            .CO(n40765));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(GND_net), .I1(n2405), .I2(VCC_net), 
            .I3(n40763), .O(n2456[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_7 (.CI(n40763), .I0(n2405), .I1(VCC_net), 
            .CO(n40764));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(GND_net), .I1(n2406), .I2(VCC_net), 
            .I3(n40762), .O(n2456[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_24_lut (.I0(n48472), .I1(timer[22]), .I2(n1[22]), 
            .I3(n39270), .O(n48474)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n39270), .I0(timer[22]), .I1(n1[22]), 
            .CO(n39271));
    SB_CARRY mod_5_add_1674_6 (.CI(n40762), .I0(n2406), .I1(VCC_net), 
            .CO(n40763));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(GND_net), .I1(n2407), .I2(VCC_net), 
            .I3(n40761), .O(n2456[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_5 (.CI(n40761), .I0(n2407), .I1(VCC_net), 
            .CO(n40762));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(GND_net), .I1(n2408), .I2(VCC_net), 
            .I3(n40760), .O(n2456[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_4 (.CI(n40760), .I0(n2408), .I1(VCC_net), 
            .CO(n40761));
    SB_LUT4 sub_14_add_2_23_lut (.I0(n48470), .I1(timer[21]), .I2(n1[21]), 
            .I3(n39269), .O(n48472)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1674_3_lut (.I0(GND_net), .I1(n2409), .I2(GND_net), 
            .I3(n40759), .O(n2456[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_3 (.CI(n40759), .I0(n2409), .I1(GND_net), 
            .CO(n40760));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(VCC_net), .O(n2456[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(GND_net), 
            .CO(n40759));
    SB_LUT4 mod_5_i1076_3_lut (.I0(n1502), .I1(n1565[28]), .I2(n1532), 
            .I3(GND_net), .O(n1601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2522), .I1(n2489), .I2(VCC_net), 
            .I3(n40758), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_i1075_3_lut (.I0(n1501), .I1(n1565[29]), .I2(n1532), 
            .I3(GND_net), .O(n1600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(GND_net), .I1(n2490), .I2(VCC_net), 
            .I3(n40757), .O(n2555[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1080_3_lut (.I0(n1506), .I1(n1565[24]), .I2(n1532), 
            .I3(GND_net), .O(n1605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1080_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1741_22 (.CI(n40757), .I0(n2490), .I1(VCC_net), 
            .CO(n40758));
    SB_LUT4 mod_5_i1074_3_lut (.I0(n1500), .I1(n1565[30]), .I2(n1532), 
            .I3(GND_net), .O(n1599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1074_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_14_add_2_23 (.CI(n39269), .I0(timer[21]), .I1(n1[21]), 
            .CO(n39270));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n48468), .I1(timer[20]), .I2(n1[20]), 
            .I3(n39268), .O(n48470)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1741_21_lut (.I0(GND_net), .I1(n2491), .I2(VCC_net), 
            .I3(n40756), .O(n2555[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_21 (.CI(n40756), .I0(n2491), .I1(VCC_net), 
            .CO(n40757));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(GND_net), .I1(n2492), .I2(VCC_net), 
            .I3(n40755), .O(n2555[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1083_3_lut (.I0(n1509), .I1(n1565[21]), .I2(n1532), 
            .I3(GND_net), .O(n1608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1081_3_lut (.I0(n1507), .I1(n1565[23]), .I2(n1532), 
            .I3(GND_net), .O(n1606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1082_3_lut (.I0(n1508), .I1(n1565[22]), .I2(n1532), 
            .I3(GND_net), .O(n1607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1082_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1741_20 (.CI(n40755), .I0(n2492), .I1(VCC_net), 
            .CO(n40756));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(GND_net), .I1(n2493), .I2(VCC_net), 
            .I3(n40754), .O(n2555[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_19 (.CI(n40754), .I0(n2493), .I1(VCC_net), 
            .CO(n40755));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(GND_net), .I1(n2494), .I2(VCC_net), 
            .I3(n40753), .O(n2555[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_18 (.CI(n40753), .I0(n2494), .I1(VCC_net), 
            .CO(n40754));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(GND_net), .I1(n2495), .I2(VCC_net), 
            .I3(n40752), .O(n2555[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1013_3_lut (.I0(n1407), .I1(n1466[24]), .I2(n1433), 
            .I3(GND_net), .O(n1506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1016_3_lut (.I0(bit_ctr[21]), .I1(n1466[21]), .I2(n1433), 
            .I3(GND_net), .O(n1509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1014_3_lut (.I0(n1408), .I1(n1466[23]), .I2(n1433), 
            .I3(GND_net), .O(n1507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1012_3_lut (.I0(n1406), .I1(n1466[25]), .I2(n1433), 
            .I3(GND_net), .O(n1505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1007_3_lut (.I0(n1401), .I1(n1466[30]), .I2(n1433), 
            .I3(GND_net), .O(n1500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1015_3_lut (.I0(n1409), .I1(n1466[22]), .I2(n1433), 
            .I3(GND_net), .O(n1508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1009_3_lut (.I0(n1403), .I1(n1466[28]), .I2(n1433), 
            .I3(GND_net), .O(n1502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1010_3_lut (.I0(n1404), .I1(n1466[27]), .I2(n1433), 
            .I3(GND_net), .O(n1503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut_adj_1610 (.I0(\state[1] ), .I1(\state[0] ), .I2(n6801), 
            .I3(GND_net), .O(n6_adj_4990));
    defparam i2_2_lut_3_lut_adj_1610.LUT_INIT = 16'h8080;
    SB_LUT4 mod_5_i1008_3_lut (.I0(n1402), .I1(n1466[29]), .I2(n1433), 
            .I3(GND_net), .O(n1501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1611 (.I0(n1501), .I1(n1503), .I2(n1502), .I3(n1504), 
            .O(n18_adj_5041));
    defparam i7_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1612 (.I0(n1508), .I1(n18_adj_5041), .I2(n1500), 
            .I3(n1499), .O(n20_adj_5042));
    defparam i9_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1613 (.I0(n1507), .I1(bit_ctr[20]), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_5043));
    defparam i4_3_lut_adj_1613.LUT_INIT = 16'heaea;
    SB_CARRY mod_5_add_1741_17 (.CI(n40752), .I0(n2495), .I1(VCC_net), 
            .CO(n40753));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(GND_net), .I1(n2496), .I2(VCC_net), 
            .I3(n40751), .O(n2555[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_16 (.CI(n40751), .I0(n2496), .I1(VCC_net), 
            .CO(n40752));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(GND_net), .I1(n2497), .I2(VCC_net), 
            .I3(n40750), .O(n2555[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_15 (.CI(n40750), .I0(n2497), .I1(VCC_net), 
            .CO(n40751));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(GND_net), .I1(n2498), .I2(VCC_net), 
            .I3(n40749), .O(n2555[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_14 (.CI(n40749), .I0(n2498), .I1(VCC_net), 
            .CO(n40750));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(GND_net), .I1(n2499), .I2(VCC_net), 
            .I3(n40748), .O(n2555[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_13 (.CI(n40748), .I0(n2499), .I1(VCC_net), 
            .CO(n40749));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(GND_net), .I1(n2500), .I2(VCC_net), 
            .I3(n40747), .O(n2555[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_12 (.CI(n40747), .I0(n2500), .I1(VCC_net), 
            .CO(n40748));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(GND_net), .I1(n2501), .I2(VCC_net), 
            .I3(n40746), .O(n2555[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_11 (.CI(n40746), .I0(n2501), .I1(VCC_net), 
            .CO(n40747));
    SB_LUT4 i10_4_lut_adj_1614 (.I0(n15_adj_5043), .I1(n20_adj_5042), .I2(n1505), 
            .I3(n1506), .O(n1532));
    defparam i10_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_22 (.CI(n39268), .I0(timer[20]), .I1(n1[20]), 
            .CO(n39269));
    SB_LUT4 mod_5_i1011_3_lut (.I0(n1405), .I1(n1466[26]), .I2(n1433), 
            .I3(GND_net), .O(n1504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1078_3_lut (.I0(n1504), .I1(n1565[26]), .I2(n1532), 
            .I3(GND_net), .O(n1603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_10_lut (.I0(GND_net), .I1(n2502), .I2(VCC_net), 
            .I3(n40745), .O(n2555[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1079_3_lut (.I0(n1505), .I1(n1565[25]), .I2(n1532), 
            .I3(GND_net), .O(n1604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_add_2_21_lut (.I0(n48466), .I1(timer[19]), .I2(n1[19]), 
            .I3(n39267), .O(n48468)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_i1084_3_lut (.I0(bit_ctr[20]), .I1(n1565[20]), .I2(n1532), 
            .I3(GND_net), .O(n1609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1077_3_lut (.I0(n1503), .I1(n1565[27]), .I2(n1532), 
            .I3(GND_net), .O(n1602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1077_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1741_10 (.CI(n40745), .I0(n2502), .I1(VCC_net), 
            .CO(n40746));
    SB_LUT4 i3_3_lut (.I0(n1602), .I1(bit_ctr[19]), .I2(n1609), .I3(GND_net), 
            .O(n15_adj_5044));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i7_4_lut_adj_1615 (.I0(n1607), .I1(n1606), .I2(n1608), .I3(n1598), 
            .O(n19_adj_5045));
    defparam i7_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut_adj_1616 (.I0(n1604), .I1(n1603), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5046));
    defparam i6_2_lut_adj_1616.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1617 (.I0(n19_adj_5045), .I1(n15_adj_5044), .I2(n1599), 
            .I3(n1605), .O(n22_adj_5047));
    defparam i10_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1618 (.I0(n1600), .I1(n22_adj_5047), .I2(n18_adj_5046), 
            .I3(n1601), .O(n1631));
    defparam i11_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_9_lut (.I0(GND_net), .I1(n2503), .I2(VCC_net), 
            .I3(n40744), .O(n2555[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_2058__i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n6801), 
            .D(n133[7]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_CARRY mod_5_add_1741_9 (.CI(n40744), .I0(n2503), .I1(VCC_net), 
            .CO(n40745));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(GND_net), .I1(n2504), .I2(VCC_net), 
            .I3(n40743), .O(n2555[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_8 (.CI(n40743), .I0(n2504), .I1(VCC_net), 
            .CO(n40744));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(GND_net), .I1(n2505), .I2(VCC_net), 
            .I3(n40742), .O(n2555[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_7 (.CI(n40742), .I0(n2505), .I1(VCC_net), 
            .CO(n40743));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(GND_net), .I1(n2506), .I2(VCC_net), 
            .I3(n40741), .O(n2555[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_6 (.CI(n40741), .I0(n2506), .I1(VCC_net), 
            .CO(n40742));
    SB_CARRY sub_14_add_2_21 (.CI(n39267), .I0(timer[19]), .I1(n1[19]), 
            .CO(n39268));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(GND_net), .I1(n2507), .I2(VCC_net), 
            .I3(n40740), .O(n2555[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_5 (.CI(n40740), .I0(n2507), .I1(VCC_net), 
            .CO(n40741));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(GND_net), .I1(n2508), .I2(VCC_net), 
            .I3(n40739), .O(n2555[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_20_lut (.I0(n48464), .I1(timer[18]), .I2(n1[18]), 
            .I3(n39266), .O(n48466)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1741_4 (.CI(n40739), .I0(n2508), .I1(VCC_net), 
            .CO(n40740));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(GND_net), .I1(n2509), .I2(GND_net), 
            .I3(n40738), .O(n2555[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_3 (.CI(n40738), .I0(n2509), .I1(GND_net), 
            .CO(n40739));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(VCC_net), .O(n2555[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(GND_net), 
            .CO(n40738));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2621), .I1(n2588), .I2(VCC_net), 
            .I3(n40737), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(GND_net), .I1(n2589), .I2(VCC_net), 
            .I3(n40736), .O(n2654[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n39266), .I0(timer[18]), .I1(n1[18]), 
            .CO(n39267));
    SB_CARRY mod_5_add_1808_23 (.CI(n40736), .I0(n2589), .I1(VCC_net), 
            .CO(n40737));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n48462), .I1(timer[17]), .I2(n1[17]), 
            .I3(n39265), .O(n48464)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1808_22_lut (.I0(GND_net), .I1(n2590), .I2(VCC_net), 
            .I3(n40735), .O(n2654[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_19 (.CI(n39265), .I0(timer[17]), .I1(n1[17]), 
            .CO(n39266));
    SB_CARRY mod_5_add_1808_22 (.CI(n40735), .I0(n2590), .I1(VCC_net), 
            .CO(n40736));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(GND_net), .I1(n2591), .I2(VCC_net), 
            .I3(n40734), .O(n2654[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_21 (.CI(n40734), .I0(n2591), .I1(VCC_net), 
            .CO(n40735));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(GND_net), .I1(n2592), .I2(VCC_net), 
            .I3(n40733), .O(n2654[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_20 (.CI(n40733), .I0(n2592), .I1(VCC_net), 
            .CO(n40734));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(GND_net), .I1(n2593), .I2(VCC_net), 
            .I3(n40732), .O(n2654[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_19 (.CI(n40732), .I0(n2593), .I1(VCC_net), 
            .CO(n40733));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(GND_net), .I1(n2594), .I2(VCC_net), 
            .I3(n40731), .O(n2654[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_18 (.CI(n40731), .I0(n2594), .I1(VCC_net), 
            .CO(n40732));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(GND_net), .I1(n2595), .I2(VCC_net), 
            .I3(n40730), .O(n2654[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_17 (.CI(n40730), .I0(n2595), .I1(VCC_net), 
            .CO(n40731));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(GND_net), .I1(n2596), .I2(VCC_net), 
            .I3(n40729), .O(n2654[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_16 (.CI(n40729), .I0(n2596), .I1(VCC_net), 
            .CO(n40730));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(GND_net), .I1(n2597), .I2(VCC_net), 
            .I3(n40728), .O(n2654[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_15 (.CI(n40728), .I0(n2597), .I1(VCC_net), 
            .CO(n40729));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(GND_net), .I1(n2598), .I2(VCC_net), 
            .I3(n40727), .O(n2654[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_18_lut (.I0(n48460), .I1(timer[16]), .I2(n1[16]), 
            .I3(n39264), .O(n48462)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_14 (.CI(n40727), .I0(n2598), .I1(VCC_net), 
            .CO(n40728));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(GND_net), .I1(n2599), .I2(VCC_net), 
            .I3(n40726), .O(n2654[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_13 (.CI(n40726), .I0(n2599), .I1(VCC_net), 
            .CO(n40727));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(GND_net), .I1(n2600), .I2(VCC_net), 
            .I3(n40725), .O(n2654[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_12 (.CI(n40725), .I0(n2600), .I1(VCC_net), 
            .CO(n40726));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(GND_net), .I1(n2601), .I2(VCC_net), 
            .I3(n40724), .O(n2654[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_11 (.CI(n40724), .I0(n2601), .I1(VCC_net), 
            .CO(n40725));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(GND_net), .I1(n2602), .I2(VCC_net), 
            .I3(n40723), .O(n2654[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_10 (.CI(n40723), .I0(n2602), .I1(VCC_net), 
            .CO(n40724));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(GND_net), .I1(n2603), .I2(VCC_net), 
            .I3(n40722), .O(n2654[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_9 (.CI(n40722), .I0(n2603), .I1(VCC_net), 
            .CO(n40723));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(GND_net), .I1(n2604), .I2(VCC_net), 
            .I3(n40721), .O(n2654[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_8 (.CI(n40721), .I0(n2604), .I1(VCC_net), 
            .CO(n40722));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(GND_net), .I1(n2605), .I2(VCC_net), 
            .I3(n40720), .O(n2654[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_7 (.CI(n40720), .I0(n2605), .I1(VCC_net), 
            .CO(n40721));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(GND_net), .I1(n2606), .I2(VCC_net), 
            .I3(n40719), .O(n2654[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_6 (.CI(n40719), .I0(n2606), .I1(VCC_net), 
            .CO(n40720));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(GND_net), .I1(n2607), .I2(VCC_net), 
            .I3(n40718), .O(n2654[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n39264), .I0(timer[16]), .I1(n1[16]), 
            .CO(n39265));
    SB_CARRY mod_5_add_1808_5 (.CI(n40718), .I0(n2607), .I1(VCC_net), 
            .CO(n40719));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(GND_net), .I1(n2608), .I2(VCC_net), 
            .I3(n40717), .O(n2654[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_4 (.CI(n40717), .I0(n2608), .I1(VCC_net), 
            .CO(n40718));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(GND_net), .I1(n2609), .I2(GND_net), 
            .I3(n40716), .O(n2654[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_3 (.CI(n40716), .I0(n2609), .I1(GND_net), 
            .CO(n40717));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(VCC_net), .O(n2654[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(GND_net), 
            .CO(n40716));
    SB_LUT4 sub_14_add_2_17_lut (.I0(n48458), .I1(timer[15]), .I2(n1[15]), 
            .I3(n39263), .O(n48460)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2720), .I1(n2687), .I2(VCC_net), 
            .I3(n40715), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(GND_net), .I1(n2688), .I2(VCC_net), 
            .I3(n40714), .O(n2753[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_24 (.CI(n40714), .I0(n2688), .I1(VCC_net), 
            .CO(n40715));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(GND_net), .I1(n2689), .I2(VCC_net), 
            .I3(n40713), .O(n2753[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_23 (.CI(n40713), .I0(n2689), .I1(VCC_net), 
            .CO(n40714));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(GND_net), .I1(n2690), .I2(VCC_net), 
            .I3(n40712), .O(n2753[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_22 (.CI(n40712), .I0(n2690), .I1(VCC_net), 
            .CO(n40713));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(GND_net), .I1(n2691), .I2(VCC_net), 
            .I3(n40711), .O(n2753[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_21 (.CI(n40711), .I0(n2691), .I1(VCC_net), 
            .CO(n40712));
    SB_CARRY sub_14_add_2_17 (.CI(n39263), .I0(timer[15]), .I1(n1[15]), 
            .CO(n39264));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(GND_net), .I1(n2692), .I2(VCC_net), 
            .I3(n40710), .O(n2753[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_20 (.CI(n40710), .I0(n2692), .I1(VCC_net), 
            .CO(n40711));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(GND_net), .I1(n2693), .I2(VCC_net), 
            .I3(n40709), .O(n2753[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_19 (.CI(n40709), .I0(n2693), .I1(VCC_net), 
            .CO(n40710));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(GND_net), .I1(n2694), .I2(VCC_net), 
            .I3(n40708), .O(n2753[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_18 (.CI(n40708), .I0(n2694), .I1(VCC_net), 
            .CO(n40709));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(GND_net), .I1(n2695), .I2(VCC_net), 
            .I3(n40707), .O(n2753[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_17 (.CI(n40707), .I0(n2695), .I1(VCC_net), 
            .CO(n40708));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(GND_net), .I1(n2696), .I2(VCC_net), 
            .I3(n40706), .O(n2753[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_16 (.CI(n40706), .I0(n2696), .I1(VCC_net), 
            .CO(n40707));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(GND_net), .I1(n2697), .I2(VCC_net), 
            .I3(n40705), .O(n2753[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_15 (.CI(n40705), .I0(n2697), .I1(VCC_net), 
            .CO(n40706));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(GND_net), .I1(n2698), .I2(VCC_net), 
            .I3(n40704), .O(n2753[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_14 (.CI(n40704), .I0(n2698), .I1(VCC_net), 
            .CO(n40705));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(GND_net), .I1(n2699), .I2(VCC_net), 
            .I3(n40703), .O(n2753[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_13 (.CI(n40703), .I0(n2699), .I1(VCC_net), 
            .CO(n40704));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(GND_net), .I1(n2700), .I2(VCC_net), 
            .I3(n40702), .O(n2753[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_12 (.CI(n40702), .I0(n2700), .I1(VCC_net), 
            .CO(n40703));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(GND_net), .I1(n2701), .I2(VCC_net), 
            .I3(n40701), .O(n2753[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_11 (.CI(n40701), .I0(n2701), .I1(VCC_net), 
            .CO(n40702));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(GND_net), .I1(n2702), .I2(VCC_net), 
            .I3(n40700), .O(n2753[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_10 (.CI(n40700), .I0(n2702), .I1(VCC_net), 
            .CO(n40701));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(GND_net), .I1(n2703), .I2(VCC_net), 
            .I3(n40699), .O(n2753[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_9 (.CI(n40699), .I0(n2703), .I1(VCC_net), 
            .CO(n40700));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(GND_net), .I1(n2704), .I2(VCC_net), 
            .I3(n40698), .O(n2753[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_8 (.CI(n40698), .I0(n2704), .I1(VCC_net), 
            .CO(n40699));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(GND_net), .I1(n2705), .I2(VCC_net), 
            .I3(n40697), .O(n2753[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_16_lut (.I0(n48456), .I1(timer[14]), .I2(n1[14]), 
            .I3(n39262), .O(n48458)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1875_7 (.CI(n40697), .I0(n2705), .I1(VCC_net), 
            .CO(n40698));
    SB_LUT4 i1_2_lut_adj_1619 (.I0(one_wire_N_679[2]), .I1(one_wire_N_679[3]), 
            .I2(GND_net), .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_1619.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1620 (.I0(one_wire_N_679[2]), .I1(n44921), .I2(GND_net), 
            .I3(GND_net), .O(n41104));
    defparam i2_2_lut_adj_1620.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1621 (.I0(one_wire_N_679[5]), .I1(one_wire_N_679[4]), 
            .I2(GND_net), .I3(GND_net), .O(n48440));   // verilog/neopixel.v(104[14:39])
    defparam i1_2_lut_adj_1621.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1622 (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[7]), 
            .I2(one_wire_N_679[6]), .I3(n48440), .O(n48446));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1623 (.I0(one_wire_N_679[10]), .I1(n27999), .I2(one_wire_N_679[9]), 
            .I3(n48446), .O(n27833));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i29741_4_lut (.I0(n27833), .I1(n41104), .I2(n4), .I3(\state[0] ), 
            .O(n45055));
    defparam i29741_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i22855_4_lut (.I0(one_wire_N_679[8]), .I1(n27999), .I2(one_wire_N_679[10]), 
            .I3(one_wire_N_679[9]), .O(n36377));
    defparam i22855_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i34388_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n49688));
    defparam i34388_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29695_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n45055), .I3(GND_net), .O(n45056));
    defparam i29695_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1624 (.I0(n45056), .I1(n49688), .I2(\state[1] ), 
            .I3(n36377), .O(n7));
    defparam i15_4_lut_adj_1624.LUT_INIT = 16'h3a0a;
    SB_LUT4 i35226_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(start_N_727));   // verilog/neopixel.v(36[4] 116[11])
    defparam i35226_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i29583_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n44939));
    defparam i29583_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i35175_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n44187));
    defparam i35175_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1625 (.I0(one_wire_N_679[2]), .I1(n44187), .I2(one_wire_N_679[3]), 
            .I3(n44921), .O(n103));
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'h45cd;
    SB_LUT4 i6_4_lut_adj_1626 (.I0(one_wire_N_679[7]), .I1(one_wire_N_679[9]), 
            .I2(n44939), .I3(n103), .O(n16_adj_5048));
    defparam i6_4_lut_adj_1626.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1627 (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[6]), 
            .I2(n16_adj_5048), .I3(one_wire_N_679[4]), .O(n6_adj_5049));
    defparam i1_4_lut_adj_1627.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_679[5]), .I1(one_wire_N_679[10]), .I2(n27999), 
            .I3(n6_adj_5049), .O(n51572));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1239_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_1239_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 mod_5_add_1875_6_lut (.I0(GND_net), .I1(n2706), .I2(VCC_net), 
            .I3(n40696), .O(n2753[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_6 (.CI(n40696), .I0(n2706), .I1(VCC_net), 
            .CO(n40697));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(GND_net), .I1(n2707), .I2(VCC_net), 
            .I3(n40695), .O(n2753[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_5 (.CI(n40695), .I0(n2707), .I1(VCC_net), 
            .CO(n40696));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(GND_net), .I1(n2708), .I2(VCC_net), 
            .I3(n40694), .O(n2753[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_4 (.CI(n40694), .I0(n2708), .I1(VCC_net), 
            .CO(n40695));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(GND_net), .I1(n2709), .I2(GND_net), 
            .I3(n40693), .O(n2753[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_3 (.CI(n40693), .I0(n2709), .I1(GND_net), 
            .CO(n40694));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n45124), .D(\neo_pixel_transmitter.done_N_742 ), 
            .R(n46958));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1875_2_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(VCC_net), .O(n2753[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(GND_net), 
            .CO(n40693));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2819), .I1(n2786), .I2(VCC_net), 
            .I3(n40692), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(GND_net), .I1(n2787), .I2(VCC_net), 
            .I3(n40691), .O(n2852[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_25 (.CI(n40691), .I0(n2787), .I1(VCC_net), 
            .CO(n40692));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(GND_net), .I1(n2788), .I2(VCC_net), 
            .I3(n40690), .O(n2852[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_24 (.CI(n40690), .I0(n2788), .I1(VCC_net), 
            .CO(n40691));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(GND_net), .I1(n2789), .I2(VCC_net), 
            .I3(n40689), .O(n2852[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_23 (.CI(n40689), .I0(n2789), .I1(VCC_net), 
            .CO(n40690));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(GND_net), .I1(n2790), .I2(VCC_net), 
            .I3(n40688), .O(n2852[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_22 (.CI(n40688), .I0(n2790), .I1(VCC_net), 
            .CO(n40689));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(GND_net), .I1(n2791), .I2(VCC_net), 
            .I3(n40687), .O(n2852[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_21 (.CI(n40687), .I0(n2791), .I1(VCC_net), 
            .CO(n40688));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(GND_net), .I1(n2792), .I2(VCC_net), 
            .I3(n40686), .O(n2852[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_20 (.CI(n40686), .I0(n2792), .I1(VCC_net), 
            .CO(n40687));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(GND_net), .I1(n2793), .I2(VCC_net), 
            .I3(n40685), .O(n2852[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_19 (.CI(n40685), .I0(n2793), .I1(VCC_net), 
            .CO(n40686));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(GND_net), .I1(n2794), .I2(VCC_net), 
            .I3(n40684), .O(n2852[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_18 (.CI(n40684), .I0(n2794), .I1(VCC_net), 
            .CO(n40685));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(GND_net), .I1(n2795), .I2(VCC_net), 
            .I3(n40683), .O(n2852[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_17 (.CI(n40683), .I0(n2795), .I1(VCC_net), 
            .CO(n40684));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(GND_net), .I1(n2796), .I2(VCC_net), 
            .I3(n40682), .O(n2852[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_16 (.CI(n40682), .I0(n2796), .I1(VCC_net), 
            .CO(n40683));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(GND_net), .I1(n2797), .I2(VCC_net), 
            .I3(n40681), .O(n2852[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_15 (.CI(n40681), .I0(n2797), .I1(VCC_net), 
            .CO(n40682));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(GND_net), .I1(n2798), .I2(VCC_net), 
            .I3(n40680), .O(n2852[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_14 (.CI(n40680), .I0(n2798), .I1(VCC_net), 
            .CO(n40681));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(GND_net), .I1(n2799), .I2(VCC_net), 
            .I3(n40679), .O(n2852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_13 (.CI(n40679), .I0(n2799), .I1(VCC_net), 
            .CO(n40680));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(GND_net), .I1(n2800), .I2(VCC_net), 
            .I3(n40678), .O(n2852[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_12 (.CI(n40678), .I0(n2800), .I1(VCC_net), 
            .CO(n40679));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(GND_net), .I1(n2801), .I2(VCC_net), 
            .I3(n40677), .O(n2852[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_11 (.CI(n40677), .I0(n2801), .I1(VCC_net), 
            .CO(n40678));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(GND_net), .I1(n2802), .I2(VCC_net), 
            .I3(n40676), .O(n2852[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_10 (.CI(n40676), .I0(n2802), .I1(VCC_net), 
            .CO(n40677));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(GND_net), .I1(n2803), .I2(VCC_net), 
            .I3(n40675), .O(n2852[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_9 (.CI(n40675), .I0(n2803), .I1(VCC_net), 
            .CO(n40676));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(GND_net), .I1(n2804), .I2(VCC_net), 
            .I3(n40674), .O(n2852[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_8 (.CI(n40674), .I0(n2804), .I1(VCC_net), 
            .CO(n40675));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(GND_net), .I1(n2805), .I2(VCC_net), 
            .I3(n40673), .O(n2852[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_7 (.CI(n40673), .I0(n2805), .I1(VCC_net), 
            .CO(n40674));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(GND_net), .I1(n2806), .I2(VCC_net), 
            .I3(n40672), .O(n2852[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_6 (.CI(n40672), .I0(n2806), .I1(VCC_net), 
            .CO(n40673));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(GND_net), .I1(n2807), .I2(VCC_net), 
            .I3(n40671), .O(n2852[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_5 (.CI(n40671), .I0(n2807), .I1(VCC_net), 
            .CO(n40672));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(GND_net), .I1(n2808), .I2(VCC_net), 
            .I3(n40670), .O(n2852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_4 (.CI(n40670), .I0(n2808), .I1(VCC_net), 
            .CO(n40671));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(GND_net), .I1(n2809), .I2(GND_net), 
            .I3(n40669), .O(n2852[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_3 (.CI(n40669), .I0(n2809), .I1(GND_net), 
            .CO(n40670));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(VCC_net), .O(n2852[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(GND_net), 
            .CO(n40669));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2918), .I1(n2885), .I2(VCC_net), 
            .I3(n40668), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(GND_net), .I1(n2886), .I2(VCC_net), 
            .I3(n40667), .O(n2951[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_26 (.CI(n40667), .I0(n2886), .I1(VCC_net), 
            .CO(n40668));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(GND_net), .I1(n2887), .I2(VCC_net), 
            .I3(n40666), .O(n2951[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_25 (.CI(n40666), .I0(n2887), .I1(VCC_net), 
            .CO(n40667));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(GND_net), .I1(n2888), .I2(VCC_net), 
            .I3(n40665), .O(n2951[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_24 (.CI(n40665), .I0(n2888), .I1(VCC_net), 
            .CO(n40666));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(GND_net), .I1(n2889), .I2(VCC_net), 
            .I3(n40664), .O(n2951[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_23 (.CI(n40664), .I0(n2889), .I1(VCC_net), 
            .CO(n40665));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(GND_net), .I1(n2890), .I2(VCC_net), 
            .I3(n40663), .O(n2951[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_22 (.CI(n40663), .I0(n2890), .I1(VCC_net), 
            .CO(n40664));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(GND_net), .I1(n2891), .I2(VCC_net), 
            .I3(n40662), .O(n2951[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_21 (.CI(n40662), .I0(n2891), .I1(VCC_net), 
            .CO(n40663));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(GND_net), .I1(n2892), .I2(VCC_net), 
            .I3(n40661), .O(n2951[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_20 (.CI(n40661), .I0(n2892), .I1(VCC_net), 
            .CO(n40662));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(GND_net), .I1(n2893), .I2(VCC_net), 
            .I3(n40660), .O(n2951[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_19 (.CI(n40660), .I0(n2893), .I1(VCC_net), 
            .CO(n40661));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(GND_net), .I1(n2894), .I2(VCC_net), 
            .I3(n40659), .O(n2951[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_18 (.CI(n40659), .I0(n2894), .I1(VCC_net), 
            .CO(n40660));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(GND_net), .I1(n2895), .I2(VCC_net), 
            .I3(n40658), .O(n2951[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_17 (.CI(n40658), .I0(n2895), .I1(VCC_net), 
            .CO(n40659));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(GND_net), .I1(n2896), .I2(VCC_net), 
            .I3(n40657), .O(n2951[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_16 (.CI(n40657), .I0(n2896), .I1(VCC_net), 
            .CO(n40658));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(GND_net), .I1(n2897), .I2(VCC_net), 
            .I3(n40656), .O(n2951[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_15 (.CI(n40656), .I0(n2897), .I1(VCC_net), 
            .CO(n40657));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(GND_net), .I1(n2898), .I2(VCC_net), 
            .I3(n40655), .O(n2951[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_14 (.CI(n40655), .I0(n2898), .I1(VCC_net), 
            .CO(n40656));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(GND_net), .I1(n2899), .I2(VCC_net), 
            .I3(n40654), .O(n2951[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_13 (.CI(n40654), .I0(n2899), .I1(VCC_net), 
            .CO(n40655));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(GND_net), .I1(n2900), .I2(VCC_net), 
            .I3(n40653), .O(n2951[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n40653), .I0(n2900), .I1(VCC_net), 
            .CO(n40654));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(GND_net), .I1(n2901), .I2(VCC_net), 
            .I3(n40652), .O(n2951[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_11 (.CI(n40652), .I0(n2901), .I1(VCC_net), 
            .CO(n40653));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(GND_net), .I1(n2902), .I2(VCC_net), 
            .I3(n40651), .O(n2951[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_10 (.CI(n40651), .I0(n2902), .I1(VCC_net), 
            .CO(n40652));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(GND_net), .I1(n2903), .I2(VCC_net), 
            .I3(n40650), .O(n2951[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_9 (.CI(n40650), .I0(n2903), .I1(VCC_net), 
            .CO(n40651));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(GND_net), .I1(n2904), .I2(VCC_net), 
            .I3(n40649), .O(n2951[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_8 (.CI(n40649), .I0(n2904), .I1(VCC_net), 
            .CO(n40650));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(GND_net), .I1(n2905), .I2(VCC_net), 
            .I3(n40648), .O(n2951[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_7 (.CI(n40648), .I0(n2905), .I1(VCC_net), 
            .CO(n40649));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(GND_net), .I1(n2906), .I2(VCC_net), 
            .I3(n40647), .O(n2951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_6 (.CI(n40647), .I0(n2906), .I1(VCC_net), 
            .CO(n40648));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(GND_net), .I1(n2907), .I2(VCC_net), 
            .I3(n40646), .O(n2951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_5 (.CI(n40646), .I0(n2907), .I1(VCC_net), 
            .CO(n40647));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(GND_net), .I1(n2908), .I2(VCC_net), 
            .I3(n40645), .O(n2951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n40645), .I0(n2908), .I1(VCC_net), 
            .CO(n40646));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(GND_net), .I1(n2909), .I2(GND_net), 
            .I3(n40644), .O(n2951[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_3 (.CI(n40644), .I0(n2909), .I1(GND_net), 
            .CO(n40645));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(VCC_net), .O(n2951[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(GND_net), 
            .CO(n40644));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n3017), .I1(n2984), .I2(VCC_net), 
            .I3(n40643), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(GND_net), .I1(n2985), .I2(VCC_net), 
            .I3(n40642), .O(n3050[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_27 (.CI(n40642), .I0(n2985), .I1(VCC_net), 
            .CO(n40643));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(GND_net), .I1(n2986), .I2(VCC_net), 
            .I3(n40641), .O(n3050[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_26 (.CI(n40641), .I0(n2986), .I1(VCC_net), 
            .CO(n40642));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(GND_net), .I1(n2987), .I2(VCC_net), 
            .I3(n40640), .O(n3050[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_25 (.CI(n40640), .I0(n2987), .I1(VCC_net), 
            .CO(n40641));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(GND_net), .I1(n2988), .I2(VCC_net), 
            .I3(n40639), .O(n3050[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_24 (.CI(n40639), .I0(n2988), .I1(VCC_net), 
            .CO(n40640));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(GND_net), .I1(n2989), .I2(VCC_net), 
            .I3(n40638), .O(n3050[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_23 (.CI(n40638), .I0(n2989), .I1(VCC_net), 
            .CO(n40639));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(GND_net), .I1(n2990), .I2(VCC_net), 
            .I3(n40637), .O(n3050[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_22 (.CI(n40637), .I0(n2990), .I1(VCC_net), 
            .CO(n40638));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(GND_net), .I1(n2991), .I2(VCC_net), 
            .I3(n40636), .O(n3050[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_21 (.CI(n40636), .I0(n2991), .I1(VCC_net), 
            .CO(n40637));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(GND_net), .I1(n2992), .I2(VCC_net), 
            .I3(n40635), .O(n3050[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_20 (.CI(n40635), .I0(n2992), .I1(VCC_net), 
            .CO(n40636));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(GND_net), .I1(n2993), .I2(VCC_net), 
            .I3(n40634), .O(n3050[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_19 (.CI(n40634), .I0(n2993), .I1(VCC_net), 
            .CO(n40635));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(GND_net), .I1(n2994), .I2(VCC_net), 
            .I3(n40633), .O(n3050[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_18 (.CI(n40633), .I0(n2994), .I1(VCC_net), 
            .CO(n40634));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(GND_net), .I1(n2995), .I2(VCC_net), 
            .I3(n40632), .O(n3050[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_17 (.CI(n40632), .I0(n2995), .I1(VCC_net), 
            .CO(n40633));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(GND_net), .I1(n2996), .I2(VCC_net), 
            .I3(n40631), .O(n3050[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_16 (.CI(n40631), .I0(n2996), .I1(VCC_net), 
            .CO(n40632));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(GND_net), .I1(n2997), .I2(VCC_net), 
            .I3(n40630), .O(n3050[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_15 (.CI(n40630), .I0(n2997), .I1(VCC_net), 
            .CO(n40631));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(GND_net), .I1(n2998), .I2(VCC_net), 
            .I3(n40629), .O(n3050[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_14 (.CI(n40629), .I0(n2998), .I1(VCC_net), 
            .CO(n40630));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(GND_net), .I1(n2999), .I2(VCC_net), 
            .I3(n40628), .O(n3050[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_13 (.CI(n40628), .I0(n2999), .I1(VCC_net), 
            .CO(n40629));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(GND_net), .I1(n3000), .I2(VCC_net), 
            .I3(n40627), .O(n3050[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_12 (.CI(n40627), .I0(n3000), .I1(VCC_net), 
            .CO(n40628));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(GND_net), .I1(n3001), .I2(VCC_net), 
            .I3(n40626), .O(n3050[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_11 (.CI(n40626), .I0(n3001), .I1(VCC_net), 
            .CO(n40627));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(GND_net), .I1(n3002), .I2(VCC_net), 
            .I3(n40625), .O(n3050[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_10 (.CI(n40625), .I0(n3002), .I1(VCC_net), 
            .CO(n40626));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(GND_net), .I1(n3003), .I2(VCC_net), 
            .I3(n40624), .O(n3050[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_9 (.CI(n40624), .I0(n3003), .I1(VCC_net), 
            .CO(n40625));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(GND_net), .I1(n3004), .I2(VCC_net), 
            .I3(n40623), .O(n3050[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_8 (.CI(n40623), .I0(n3004), .I1(VCC_net), 
            .CO(n40624));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(GND_net), .I1(n3005), .I2(VCC_net), 
            .I3(n40622), .O(n3050[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_7 (.CI(n40622), .I0(n3005), .I1(VCC_net), 
            .CO(n40623));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(GND_net), .I1(n3006), .I2(VCC_net), 
            .I3(n40621), .O(n3050[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_6 (.CI(n40621), .I0(n3006), .I1(VCC_net), 
            .CO(n40622));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(GND_net), .I1(n3007), .I2(VCC_net), 
            .I3(n40620), .O(n3050[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_5 (.CI(n40620), .I0(n3007), .I1(VCC_net), 
            .CO(n40621));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(GND_net), .I1(n3008), .I2(VCC_net), 
            .I3(n40619), .O(n3050[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_4 (.CI(n40619), .I0(n3008), .I1(VCC_net), 
            .CO(n40620));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(GND_net), .I1(n32241), .I2(GND_net), 
            .I3(n40618), .O(n3050[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_3 (.CI(n40618), .I0(n32241), .I1(GND_net), 
            .CO(n40619));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(VCC_net), .O(n3050[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(GND_net), 
            .CO(n40618));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n40617), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n40616), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n40616), .I0(n3084), .I1(n3116), .CO(n40617));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n40615), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n40615), .I0(n3085), .I1(n3116), .CO(n40616));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n40614), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n40614), .I0(n3086), .I1(n3116), .CO(n40615));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n40613), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n40613), .I0(n3087), .I1(n3116), .CO(n40614));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n40612), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n40612), .I0(n3088), .I1(n3116), .CO(n40613));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n40611), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n40611), .I0(n3089), .I1(n3116), .CO(n40612));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n40610), .O(n49_adj_5050)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n40610), .I0(n3090), .I1(n3116), .CO(n40611));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n40609), .O(n47_adj_5051)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n40609), .I0(n3091), .I1(n3116), .CO(n40610));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n40608), .O(n45_adj_5052)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n40608), .I0(n3092), .I1(n3116), .CO(n40609));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n40607), .O(n43_adj_5053)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n40607), .I0(n3093), .I1(n3116), .CO(n40608));
    SB_CARRY sub_14_add_2_16 (.CI(n39262), .I0(timer[14]), .I1(n1[14]), 
            .CO(n39263));
    SB_LUT4 sub_14_add_2_15_lut (.I0(n48454), .I1(timer[13]), .I2(n1[13]), 
            .I3(n39261), .O(n48456)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_DFFESR bit_ctr_2058__i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n6801), 
            .D(n133[6]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n40606), .O(n41_adj_5055)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n40606), .I0(n3094), .I1(n3116), .CO(n40607));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n40605), .O(n39_adj_5056)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n40605), .I0(n3095), .I1(n3116), .CO(n40606));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n40604), .O(n37_adj_5057)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n40604), .I0(n3096), .I1(n3116), .CO(n40605));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n40603), .O(n35_adj_5058)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n40603), .I0(n3097), .I1(n3116), .CO(n40604));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n40602), .O(n33_adj_5059)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n40602), .I0(n3098), .I1(n3116), .CO(n40603));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n40601), .O(n31_adj_5060)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n40601), .I0(n3099), .I1(n3116), .CO(n40602));
    SB_DFFESR bit_ctr_2058__i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n6801), 
            .D(n133[5]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n40600), .O(n29_adj_5061)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n40600), .I0(n3100), .I1(n3116), .CO(n40601));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n40599), .O(n27_adj_5062)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_2058__i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n6801), 
            .D(n133[4]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_CARRY mod_5_add_2143_11 (.CI(n40599), .I0(n3101), .I1(n3116), .CO(n40600));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n40598), .O(n25_adj_5063)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n40598), .I0(n3102), .I1(n3116), .CO(n40599));
    SB_DFFESR bit_ctr_2058__i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n6801), 
            .D(n133[3]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n40597), .O(n23_adj_5064)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_2058__i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n6801), 
            .D(n133[2]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_CARRY mod_5_add_2143_9 (.CI(n40597), .I0(n3103), .I1(n3116), .CO(n40598));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n40596), .O(n21_adj_5065)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n40596), .I0(n3104), .I1(n3116), .CO(n40597));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n40595), .O(n19_adj_5066)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n40595), .I0(n3105), .I1(n3116), .CO(n40596));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n40594), .O(n17_adj_5067)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n40594), .I0(n3106), .I1(n3116), .CO(n40595));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n40593), .O(n15_adj_5068)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n40593), .I0(n3107), .I1(n3116), .CO(n40594));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n40592), .O(n13_adj_5069)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n40592), .I0(n3108), .I1(n3116), .CO(n40593));
    SB_CARRY sub_14_add_2_15 (.CI(n39261), .I0(timer[13]), .I1(n1[13]), 
            .CO(n39262));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n51355), 
            .I3(n40591), .O(n11_adj_5070)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n40591), .I0(n3109), .I1(n51355), .CO(n40592));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n51355), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 bit_ctr_1__bdd_4_lut (.I0(bit_ctr[1]), .I1(n48887), .I2(n48888), 
            .I3(bit_ctr[2]), .O(n51417));
    defparam bit_ctr_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51417_bdd_4_lut (.I0(n51417), .I1(n48828), .I2(n48827), .I3(bit_ctr[2]), 
            .O(n51420));
    defparam n51417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF timer_2057__i1 (.Q(timer[1]), .C(CLK_c), .D(n133_adj_5090[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i2 (.Q(timer[2]), .C(CLK_c), .D(n133_adj_5090[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i3 (.Q(timer[3]), .C(CLK_c), .D(n133_adj_5090[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i4 (.Q(timer[4]), .C(CLK_c), .D(n133_adj_5090[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i5 (.Q(timer[5]), .C(CLK_c), .D(n133_adj_5090[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i6 (.Q(timer[6]), .C(CLK_c), .D(n133_adj_5090[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i7 (.Q(timer[7]), .C(CLK_c), .D(n133_adj_5090[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i8 (.Q(timer[8]), .C(CLK_c), .D(n133_adj_5090[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i9 (.Q(timer[9]), .C(CLK_c), .D(n133_adj_5090[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i10 (.Q(timer[10]), .C(CLK_c), .D(n133_adj_5090[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i11 (.Q(timer[11]), .C(CLK_c), .D(n133_adj_5090[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i12 (.Q(timer[12]), .C(CLK_c), .D(n133_adj_5090[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i13 (.Q(timer[13]), .C(CLK_c), .D(n133_adj_5090[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i14 (.Q(timer[14]), .C(CLK_c), .D(n133_adj_5090[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i15 (.Q(timer[15]), .C(CLK_c), .D(n133_adj_5090[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i16 (.Q(timer[16]), .C(CLK_c), .D(n133_adj_5090[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i17 (.Q(timer[17]), .C(CLK_c), .D(n133_adj_5090[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i18 (.Q(timer[18]), .C(CLK_c), .D(n133_adj_5090[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i19 (.Q(timer[19]), .C(CLK_c), .D(n133_adj_5090[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i20 (.Q(timer[20]), .C(CLK_c), .D(n133_adj_5090[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i21 (.Q(timer[21]), .C(CLK_c), .D(n133_adj_5090[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i22 (.Q(timer[22]), .C(CLK_c), .D(n133_adj_5090[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i23 (.Q(timer[23]), .C(CLK_c), .D(n133_adj_5090[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i24 (.Q(timer[24]), .C(CLK_c), .D(n133_adj_5090[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i25 (.Q(timer[25]), .C(CLK_c), .D(n133_adj_5090[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i26 (.Q(timer[26]), .C(CLK_c), .D(n133_adj_5090[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i27 (.Q(timer[27]), .C(CLK_c), .D(n133_adj_5090[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i28 (.Q(timer[28]), .C(CLK_c), .D(n133_adj_5090[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i29 (.Q(timer[29]), .C(CLK_c), .D(n133_adj_5090[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i30 (.Q(timer[30]), .C(CLK_c), .D(n133_adj_5090[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2057__i31 (.Q(timer[31]), .C(CLK_c), .D(n133_adj_5090[31]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n51355), 
            .CO(n40591));
    SB_DFFE state_i1 (.Q(\state[1] ), .C(CLK_c), .E(VCC_net), .D(n29633));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n29623));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_679[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n39260), .O(n48454)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_14 (.CI(n39260), .I0(timer[12]), .I1(n1[12]), 
            .CO(n39261));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n39259), .O(one_wire_N_679[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n39259), .I0(timer[11]), .I1(n1[11]), 
            .CO(n39260));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n39258), .O(one_wire_N_679[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n39258), .I0(timer[10]), .I1(n1[10]), 
            .CO(n39259));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n39257), .O(one_wire_N_679[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n39257), .I0(timer[9]), .I1(n1[9]), 
            .CO(n39258));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n39256), .O(one_wire_N_679[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n39256), .I0(timer[8]), .I1(n1[8]), 
            .CO(n39257));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n39255), .O(one_wire_N_679[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n39255), .I0(timer[7]), .I1(n1[7]), .CO(n39256));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n39254), .O(one_wire_N_679[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n39254), .I0(timer[6]), .I1(n1[6]), .CO(n39255));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n39253), .O(one_wire_N_679[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n39253), .I0(timer[5]), .I1(n1[5]), .CO(n39254));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n39252), .O(one_wire_N_679[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n39252), .I0(timer[4]), .I1(n1[4]), .CO(n39253));
    SB_LUT4 bit_ctr_1__bdd_4_lut_35970 (.I0(bit_ctr[1]), .I1(n48866), .I2(n48867), 
            .I3(bit_ctr[2]), .O(n51411));
    defparam bit_ctr_1__bdd_4_lut_35970.LUT_INIT = 16'he4aa;
    SB_LUT4 n51411_bdd_4_lut (.I0(n51411), .I1(n48861), .I2(n48860), .I3(bit_ctr[2]), 
            .O(n51414));
    defparam n51411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n39251), .O(one_wire_N_679[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n39251), .I0(timer[3]), .I1(n1[3]), .CO(n39252));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n39250), .O(one_wire_N_679[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1532), .I1(n1499), .I2(VCC_net), 
            .I3(n39382), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(GND_net), .I1(n1500), .I2(VCC_net), 
            .I3(n39381), .O(n1565[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_12 (.CI(n39381), .I0(n1500), .I1(VCC_net), 
            .CO(n39382));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(GND_net), .I1(n1501), .I2(VCC_net), 
            .I3(n39380), .O(n1565[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_11 (.CI(n39380), .I0(n1501), .I1(VCC_net), 
            .CO(n39381));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(GND_net), .I1(n1502), .I2(VCC_net), 
            .I3(n39379), .O(n1565[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_10 (.CI(n39379), .I0(n1502), .I1(VCC_net), 
            .CO(n39380));
    SB_CARRY sub_14_add_2_4 (.CI(n39250), .I0(timer[2]), .I1(n1[2]), .CO(n39251));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(GND_net), .I1(n1503), .I2(VCC_net), 
            .I3(n39378), .O(n1565[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_679[3]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n39249), .O(n44921)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1071_9 (.CI(n39378), .I0(n1503), .I1(VCC_net), 
            .CO(n39379));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(GND_net), .I1(n1504), .I2(VCC_net), 
            .I3(n39377), .O(n1565[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_8 (.CI(n39377), .I0(n1504), .I1(VCC_net), 
            .CO(n39378));
    SB_CARRY sub_14_add_2_3 (.CI(n39249), .I0(timer[1]), .I1(n1[1]), .CO(n39250));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(GND_net), .I1(n1505), .I2(VCC_net), 
            .I3(n39376), .O(n1565[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_7 (.CI(n39376), .I0(n1505), .I1(VCC_net), 
            .CO(n39377));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(GND_net), .I1(n1506), .I2(VCC_net), 
            .I3(n39375), .O(n1565[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_6 (.CI(n39375), .I0(n1506), .I1(VCC_net), 
            .CO(n39376));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(GND_net), .I1(n1507), .I2(VCC_net), 
            .I3(n39374), .O(n1565[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_5 (.CI(n39374), .I0(n1507), .I1(VCC_net), 
            .CO(n39375));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(GND_net), .I1(n1508), .I2(VCC_net), 
            .I3(n39373), .O(n1565[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_4 (.CI(n39373), .I0(n1508), .I1(VCC_net), 
            .CO(n39374));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(GND_net), .I1(n1509), .I2(GND_net), 
            .I3(n39372), .O(n1565[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_3 (.CI(n39372), .I0(n1509), .I1(GND_net), 
            .CO(n39373));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(VCC_net), .O(n1565[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(GND_net), 
            .CO(n39372));
    SB_LUT4 i35915_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51353));
    defparam i35915_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35224_2_lut (.I0(n971[28]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50662));   // verilog/neopixel.v(22[26:36])
    defparam i35224_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i35223_2_lut (.I0(n971[29]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50661));   // verilog/neopixel.v(22[26:36])
    defparam i35223_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i35227_2_lut (.I0(n971[30]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50665));   // verilog/neopixel.v(22[26:36])
    defparam i35227_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n39249));
    SB_LUT4 mod_5_i675_3_lut (.I0(n26374), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i673_3_lut (.I0(n29447), .I1(n971[29]), .I2(n2), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i674_3_lut (.I0(n29401), .I1(n971[28]), .I2(n2), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35245_2_lut (.I0(n971[31]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50683));   // verilog/neopixel.v(22[26:36])
    defparam i35245_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n7_adj_5071));
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i5_4_lut_adj_1628 (.I0(n50683), .I1(n7_adj_5071), .I2(n1006), 
            .I3(n8), .O(n1037));
    defparam i5_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_2058__i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n6801), 
            .D(n133[1]), .R(n29524));   // verilog/neopixel.v(69[23:32])
    SB_LUT4 i33390_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48827));
    defparam i33390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33391_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48828));
    defparam i33391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33451_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48888));
    defparam i33451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33450_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48887));
    defparam i33450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35917_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51355));
    defparam i35917_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i2089_3_lut (.I0(n2995), .I1(n3050[20]), .I2(n3017), 
            .I3(GND_net), .O(n3094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2087_3_lut (.I0(n2993), .I1(n3050[22]), .I2(n3017), 
            .I3(GND_net), .O(n3092));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18724_3_lut (.I0(n32241), .I1(n3050[6]), .I2(n3017), .I3(GND_net), 
            .O(n3108));
    defparam i18724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2091_3_lut (.I0(n2997), .I1(n3050[18]), .I2(n3017), 
            .I3(GND_net), .O(n3096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2093_3_lut (.I0(n2999), .I1(n3050[16]), .I2(n3017), 
            .I3(GND_net), .O(n3098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2101_3_lut (.I0(n3007), .I1(n3050[8]), .I2(n3017), 
            .I3(GND_net), .O(n3106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2097_3_lut (.I0(n3003), .I1(n3050[12]), .I2(n3017), 
            .I3(GND_net), .O(n3102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2098_3_lut (.I0(n3004), .I1(n3050[11]), .I2(n3017), 
            .I3(GND_net), .O(n3103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2079_3_lut (.I0(n2985), .I1(n3050[30]), .I2(n3017), 
            .I3(GND_net), .O(n3084));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2080_3_lut (.I0(n2986), .I1(n3050[29]), .I2(n3017), 
            .I3(GND_net), .O(n3085));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2102_3_lut (.I0(n3008), .I1(n3050[7]), .I2(n3017), 
            .I3(GND_net), .O(n3107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18743_3_lut (.I0(bit_ctr[5]), .I1(n3050[5]), .I2(n3017), 
            .I3(GND_net), .O(n3109));
    defparam i18743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2094_3_lut (.I0(n3000), .I1(n3050[15]), .I2(n3017), 
            .I3(GND_net), .O(n3099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2096_3_lut (.I0(n3002), .I1(n3050[13]), .I2(n3017), 
            .I3(GND_net), .O(n3101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2085_3_lut (.I0(n2991), .I1(n3050[24]), .I2(n3017), 
            .I3(GND_net), .O(n3090));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2082_3_lut (.I0(n2988), .I1(n3050[27]), .I2(n3017), 
            .I3(GND_net), .O(n3087));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2084_3_lut (.I0(n2990), .I1(n3050[25]), .I2(n3017), 
            .I3(GND_net), .O(n3089));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2092_3_lut (.I0(n2998), .I1(n3050[17]), .I2(n3017), 
            .I3(GND_net), .O(n3097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2100_3_lut (.I0(n3006), .I1(n3050[9]), .I2(n3017), 
            .I3(GND_net), .O(n3105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2099_3_lut (.I0(n3005), .I1(n3050[10]), .I2(n3017), 
            .I3(GND_net), .O(n3104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2090_3_lut (.I0(n2996), .I1(n3050[19]), .I2(n3017), 
            .I3(GND_net), .O(n3095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2088_3_lut (.I0(n2994), .I1(n3050[21]), .I2(n3017), 
            .I3(GND_net), .O(n3093));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2083_3_lut (.I0(n2989), .I1(n3050[26]), .I2(n3017), 
            .I3(GND_net), .O(n3088));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2081_3_lut (.I0(n2987), .I1(n3050[28]), .I2(n3017), 
            .I3(GND_net), .O(n3086));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2086_3_lut (.I0(n2992), .I1(n3050[23]), .I2(n3017), 
            .I3(GND_net), .O(n3091));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2095_3_lut (.I0(n3001), .I1(n3050[14]), .I2(n3017), 
            .I3(GND_net), .O(n3100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_2_lut (.I0(n3100), .I1(n3091), .I2(GND_net), .I3(GND_net), 
            .O(n36_adj_5072));
    defparam i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut_adj_1629 (.I0(n3095), .I1(n3104), .I2(n3105), .I3(n3097), 
            .O(n46_adj_5073));
    defparam i19_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1630 (.I0(n3086), .I1(n3088), .I2(n3083), .I3(n3093), 
            .O(n42_adj_5074));
    defparam i15_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1631 (.I0(bit_ctr[4]), .I1(n3099), .I2(n3109), 
            .I3(GND_net), .O(n34_adj_5075));
    defparam i7_3_lut_adj_1631.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1632 (.I0(n3089), .I1(n3087), .I2(n3090), .I3(n3101), 
            .O(n43_adj_5076));
    defparam i16_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1633 (.I0(n3103), .I1(n46_adj_5073), .I2(n36_adj_5072), 
            .I3(n3102), .O(n50));
    defparam i23_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1634 (.I0(n3107), .I1(n42_adj_5074), .I2(n3085), 
            .I3(n3084), .O(n48_adj_5077));
    defparam i21_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1635 (.I0(n43_adj_5076), .I1(n3092), .I2(n34_adj_5075), 
            .I3(n3094), .O(n49_adj_5078));
    defparam i22_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1636 (.I0(n3106), .I1(n3098), .I2(n3096), .I3(n3108), 
            .O(n47_adj_5079));
    defparam i20_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1637 (.I0(n47_adj_5079), .I1(n49_adj_5078), .I2(n48_adj_5077), 
            .I3(n50), .O(n3116));
    defparam i26_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i18740_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n29408));   // verilog/neopixel.v(18[12:19])
    defparam i18740_3_lut_4_lut.LUT_INIT = 16'hdb6d;
    SB_LUT4 i18742_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n26382));   // verilog/neopixel.v(18[12:19])
    defparam i18742_3_lut_4_lut.LUT_INIT = 16'hb6db;
    SB_LUT4 mod_5_i606_3_lut_3_lut_4_lut_3_lut (.I0(bit_ctr[27]), .I1(n26382), 
            .I2(n29408), .I3(GND_net), .O(n29447));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_3_lut_4_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i34580_3_lut_4_lut_3_lut (.I0(bit_ctr[27]), .I1(n26382), .I2(n29408), 
            .I3(GND_net), .O(n29401));   // verilog/neopixel.v(22[26:36])
    defparam i34580_3_lut_4_lut_3_lut.LUT_INIT = 16'h1919;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(bit_ctr[27]), .I1(n26382), .I2(n29408), 
            .I3(GND_net), .O(n26374));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h8585;
    SB_LUT4 mod_5_i2018_3_lut (.I0(n2892), .I1(n2951[24]), .I2(n2918), 
            .I3(GND_net), .O(n2991));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_4_lut (.I0(bit_ctr[26]), .I1(n26374), .I2(n29447), 
            .I3(n29401), .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 mod_5_i2016_3_lut (.I0(n2890), .I1(n2951[26]), .I2(n2918), 
            .I3(GND_net), .O(n2989));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2017_3_lut (.I0(n2891), .I1(n2951[25]), .I2(n2918), 
            .I3(GND_net), .O(n2990));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2015_3_lut (.I0(n2889), .I1(n2951[27]), .I2(n2918), 
            .I3(GND_net), .O(n2988));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2035_3_lut (.I0(n2909), .I1(n2951[7]), .I2(n2918), 
            .I3(GND_net), .O(n3008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2030_3_lut (.I0(n2904), .I1(n2951[12]), .I2(n2918), 
            .I3(GND_net), .O(n3003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2023_3_lut (.I0(n2897), .I1(n2951[19]), .I2(n2918), 
            .I3(GND_net), .O(n2996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2031_3_lut (.I0(n2905), .I1(n2951[11]), .I2(n2918), 
            .I3(GND_net), .O(n3004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2026_3_lut (.I0(n2900), .I1(n2951[16]), .I2(n2918), 
            .I3(GND_net), .O(n2999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2027_3_lut (.I0(n2901), .I1(n2951[15]), .I2(n2918), 
            .I3(GND_net), .O(n3000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2032_3_lut (.I0(n2906), .I1(n2951[10]), .I2(n2918), 
            .I3(GND_net), .O(n3005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2022_3_lut (.I0(n2896), .I1(n2951[20]), .I2(n2918), 
            .I3(GND_net), .O(n2995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2021_3_lut (.I0(n2895), .I1(n2951[21]), .I2(n2918), 
            .I3(GND_net), .O(n2994));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2020_3_lut (.I0(n2894), .I1(n2951[22]), .I2(n2918), 
            .I3(GND_net), .O(n2993));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2033_3_lut (.I0(n2907), .I1(n2951[9]), .I2(n2918), 
            .I3(GND_net), .O(n3006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2019_3_lut (.I0(n2893), .I1(n2951[23]), .I2(n2918), 
            .I3(GND_net), .O(n2992));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2028_3_lut (.I0(n2902), .I1(n2951[14]), .I2(n2918), 
            .I3(GND_net), .O(n3001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2025_3_lut (.I0(n2899), .I1(n2951[17]), .I2(n2918), 
            .I3(GND_net), .O(n2998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2024_3_lut (.I0(n2898), .I1(n2951[18]), .I2(n2918), 
            .I3(GND_net), .O(n2997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2029_3_lut (.I0(n2903), .I1(n2951[13]), .I2(n2918), 
            .I3(GND_net), .O(n3002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2014_3_lut (.I0(n2888), .I1(n2951[28]), .I2(n2918), 
            .I3(GND_net), .O(n2987));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2013_3_lut (.I0(n2887), .I1(n2951[29]), .I2(n2918), 
            .I3(GND_net), .O(n2986));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2012_3_lut (.I0(n2886), .I1(n2951[30]), .I2(n2918), 
            .I3(GND_net), .O(n2985));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18723_3_lut (.I0(bit_ctr[6]), .I1(n2951[6]), .I2(n2918), 
            .I3(GND_net), .O(n32241));
    defparam i18723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2034_3_lut (.I0(n2908), .I1(n2951[8]), .I2(n2918), 
            .I3(GND_net), .O(n3007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[5]), .I1(n3007), .I2(n32241), .I3(GND_net), 
            .O(n35_adj_5080));   // verilog/neopixel.v(22[26:36])
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1638 (.I0(n3002), .I1(n2997), .I2(n2998), .I3(n3001), 
            .O(n43_adj_5081));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1639 (.I0(n2985), .I1(n2986), .I2(n2984), .I3(n2987), 
            .O(n40_adj_5082));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1640 (.I0(n2995), .I1(n3005), .I2(n3000), .I3(n2999), 
            .O(n45_adj_5083));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1641 (.I0(n2992), .I1(n3006), .I2(n2993), .I3(n2994), 
            .O(n42_adj_5084));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1642 (.I0(n43_adj_5081), .I1(n35_adj_5080), .I2(n3004), 
            .I3(n2996), .O(n48_adj_5085));   // verilog/neopixel.v(22[26:36])
    defparam i22_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1643 (.I0(n2988), .I1(n2990), .I2(n2989), .I3(n2991), 
            .O(n41_adj_5086));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1644 (.I0(n45_adj_5083), .I1(n3003), .I2(n40_adj_5082), 
            .I3(n3008), .O(n49_adj_5087));   // verilog/neopixel.v(22[26:36])
    defparam i23_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n49_adj_5087), .I1(n41_adj_5086), .I2(n48_adj_5085), 
            .I3(n42_adj_5084), .O(n3017));   // verilog/neopixel.v(22[26:36])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(n23_adj_5064), .I1(n33_adj_5059), .I2(n21_adj_5065), 
            .I3(n13_adj_5069), .O(n48048));
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n27_adj_5062), .I1(n11_adj_5070), .I2(n17_adj_5067), 
            .I3(n15_adj_5068), .O(n48050));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(n19_adj_5066), .I1(n37_adj_5057), .I2(n39_adj_5056), 
            .I3(n31_adj_5060), .O(n48052));
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1648 (.I0(n25_adj_5063), .I1(n35_adj_5058), .I2(n41_adj_5055), 
            .I3(n29_adj_5061), .O(n48054));
    defparam i1_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i22667_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n36185));
    defparam i22667_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1649 (.I0(n48054), .I1(n48052), .I2(n48050), 
            .I3(n48048), .O(n48062));
    defparam i1_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(n45_adj_5052), .I1(n48062), .I2(n43_adj_5053), 
            .I3(n36185), .O(n48066));
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n51), .I1(n49_adj_5050), .I2(n47_adj_5051), 
            .I3(n48066), .O(n48072));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1652 (.I0(n57), .I1(n55), .I2(n53), .I3(n48072), 
            .O(n48078));
    defparam i1_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(n61), .I1(n63), .I2(n59), .I3(n48078), 
            .O(n41260));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1654 (.I0(\state[1] ), .I1(n36377), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n45525));
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'hf5fd;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(n45525), .I1(n45055), .I2(\state[1] ), 
            .I3(n27992), .O(n29323));
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'ha0a8;
    SB_LUT4 i34571_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n41260), .I3(GND_net), 
            .O(color_bit_N_722[4]));
    defparam i34571_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i34712_3_lut (.I0(n51420), .I1(bit_ctr[3]), .I2(n41260), .I3(GND_net), 
            .O(n49685));
    defparam i34712_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i35117_4_lut (.I0(n51360), .I1(n51414), .I2(bit_ctr[3]), .I3(n41260), 
            .O(n50555));   // verilog/neopixel.v(22[26:36])
    defparam i35117_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i21620_4_lut (.I0(n50555), .I1(\state_3__N_528[1] ), .I2(n49685), 
            .I3(color_bit_N_722[4]), .O(state_3__N_528[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i21620_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i34435_2_lut_3_lut (.I0(LED_c), .I1(\state_3__N_528[1] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n49686));
    defparam i34435_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i34424_3_lut_4_lut (.I0(n27833), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n4), .O(n49666));
    defparam i34424_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 mod_5_i941_3_lut (.I0(n1303), .I1(n1367[29]), .I2(n1334), 
            .I3(GND_net), .O(n1402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i943_3_lut (.I0(n1305), .I1(n1367[27]), .I2(n1334), 
            .I3(GND_net), .O(n1404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i940_3_lut (.I0(n1302), .I1(n1367[30]), .I2(n1334), 
            .I3(GND_net), .O(n1401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i945_3_lut (.I0(n1307), .I1(n1367[25]), .I2(n1334), 
            .I3(GND_net), .O(n1406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i947_3_lut (.I0(n1309), .I1(n1367[23]), .I2(n1334), 
            .I3(GND_net), .O(n1408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i944_3_lut (.I0(n1306), .I1(n1367[26]), .I2(n1334), 
            .I3(GND_net), .O(n1405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i942_3_lut (.I0(n1304), .I1(n1367[28]), .I2(n1334), 
            .I3(GND_net), .O(n1403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i946_3_lut (.I0(n1308), .I1(n1367[24]), .I2(n1334), 
            .I3(GND_net), .O(n1407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i948_3_lut (.I0(bit_ctr[22]), .I1(n1367[22]), .I2(n1334), 
            .I3(GND_net), .O(n1409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22671_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n36189));
    defparam i22671_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1656 (.I0(n1406), .I1(n1401), .I2(n1400), .I3(n36189), 
            .O(n16_adj_5088));   // verilog/neopixel.v(22[26:36])
    defparam i6_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1657 (.I0(n1407), .I1(n1403), .I2(n1405), .I3(n1408), 
            .O(n17_adj_5089));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1658 (.I0(n17_adj_5089), .I1(n1404), .I2(n16_adj_5088), 
            .I3(n1402), .O(n1433));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 i34731_3_lut_4_lut (.I0(n27833), .I1(n50168), .I2(start), 
            .I3(\state[1] ), .O(n50169));
    defparam i34731_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34397_2_lut_3_lut (.I0(one_wire_N_679[2]), .I1(one_wire_N_679[3]), 
            .I2(start), .I3(GND_net), .O(n49673));
    defparam i34397_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n36377), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n46958));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 bit_ctr_1__bdd_4_lut_35965 (.I0(bit_ctr[1]), .I1(n48878), .I2(n48879), 
            .I3(bit_ctr[2]), .O(n51357));
    defparam bit_ctr_1__bdd_4_lut_35965.LUT_INIT = 16'he4aa;
    SB_LUT4 n51357_bdd_4_lut (.I0(n51357), .I1(n48738), .I2(n48737), .I3(bit_ctr[2]), 
            .O(n51360));
    defparam n51357_bdd_4_lut.LUT_INIT = 16'haad8;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (n1653, ENCODER0_B_N_keep, ENCODER0_A_N_keep, 
            \a_new[1] , b_prev, n29689, n1617, direction_N_3907, encoder0_position, 
            GND_net, VCC_net) /* synthesis lattice_noprune=1 */ ;
    input n1653;
    input ENCODER0_B_N_keep;
    input ENCODER0_A_N_keep;
    output \a_new[1] ;
    output b_prev;
    input n29689;
    output n1617;
    output direction_N_3907;
    output [31:0]encoder0_position;
    input GND_net;
    input VCC_net;
    
    
    wire a_prev_N_3913, debounce_cnt;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire n29691, a_prev, n29690;
    wire [31:0]n133;
    
    wire direction_N_3906, n40554, n40553, n40552, n40551, n40550, 
        n40549, n40548, n40547, n40546, n40545, n40544, n40543, 
        n40542, n40541, n40540, n40539, n40538, n40537, n40536, 
        n40535, n40534, n40533, n40532, n40531, n40530, n40529, 
        n40528, n40527, n40526, n40525, n40524, direction_N_3910;
    
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1653), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1653), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1653), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i35188_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i35188_4_lut.LUT_INIT = 16'h8421;
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1653), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1653), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1653), .D(n29691));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1653), .D(n29690));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1617), .C(n1653), .D(n29689));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2066__i0 (.Q(encoder0_position[0]), .C(n1653), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 i16164_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29691));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16164_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE position_2066__i1 (.Q(encoder0_position[1]), .C(n1653), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 i16163_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n29690));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16163_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFFE position_2066__i2 (.Q(encoder0_position[2]), .C(n1653), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i3 (.Q(encoder0_position[3]), .C(n1653), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i4 (.Q(encoder0_position[4]), .C(n1653), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i5 (.Q(encoder0_position[5]), .C(n1653), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i6 (.Q(encoder0_position[6]), .C(n1653), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i7 (.Q(encoder0_position[7]), .C(n1653), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i8 (.Q(encoder0_position[8]), .C(n1653), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i9 (.Q(encoder0_position[9]), .C(n1653), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i10 (.Q(encoder0_position[10]), .C(n1653), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i11 (.Q(encoder0_position[11]), .C(n1653), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i12 (.Q(encoder0_position[12]), .C(n1653), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i13 (.Q(encoder0_position[13]), .C(n1653), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i14 (.Q(encoder0_position[14]), .C(n1653), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i15 (.Q(encoder0_position[15]), .C(n1653), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i16 (.Q(encoder0_position[16]), .C(n1653), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i17 (.Q(encoder0_position[17]), .C(n1653), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i18 (.Q(encoder0_position[18]), .C(n1653), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i19 (.Q(encoder0_position[19]), .C(n1653), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i20 (.Q(encoder0_position[20]), .C(n1653), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i21 (.Q(encoder0_position[21]), .C(n1653), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i22 (.Q(encoder0_position[22]), .C(n1653), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i23 (.Q(encoder0_position[23]), .C(n1653), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i24 (.Q(encoder0_position[24]), .C(n1653), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i25 (.Q(encoder0_position[25]), .C(n1653), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i26 (.Q(encoder0_position[26]), .C(n1653), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i27 (.Q(encoder0_position[27]), .C(n1653), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i28 (.Q(encoder0_position[28]), .C(n1653), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i29 (.Q(encoder0_position[29]), .C(n1653), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i30 (.Q(encoder0_position[30]), .C(n1653), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2066__i31 (.Q(encoder0_position[31]), .C(n1653), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 position_2066_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[31]), .I3(n40554), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2066_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[30]), .I3(n40553), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_32 (.CI(n40553), .I0(direction_N_3906), 
            .I1(encoder0_position[30]), .CO(n40554));
    SB_LUT4 position_2066_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[29]), .I3(n40552), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_31 (.CI(n40552), .I0(direction_N_3906), 
            .I1(encoder0_position[29]), .CO(n40553));
    SB_LUT4 position_2066_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[28]), .I3(n40551), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_30 (.CI(n40551), .I0(direction_N_3906), 
            .I1(encoder0_position[28]), .CO(n40552));
    SB_LUT4 position_2066_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[27]), .I3(n40550), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_29 (.CI(n40550), .I0(direction_N_3906), 
            .I1(encoder0_position[27]), .CO(n40551));
    SB_LUT4 position_2066_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[26]), .I3(n40549), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_28 (.CI(n40549), .I0(direction_N_3906), 
            .I1(encoder0_position[26]), .CO(n40550));
    SB_LUT4 position_2066_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[25]), .I3(n40548), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_27 (.CI(n40548), .I0(direction_N_3906), 
            .I1(encoder0_position[25]), .CO(n40549));
    SB_LUT4 position_2066_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[24]), .I3(n40547), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_26 (.CI(n40547), .I0(direction_N_3906), 
            .I1(encoder0_position[24]), .CO(n40548));
    SB_LUT4 position_2066_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[23]), .I3(n40546), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_25 (.CI(n40546), .I0(direction_N_3906), 
            .I1(encoder0_position[23]), .CO(n40547));
    SB_LUT4 position_2066_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[22]), .I3(n40545), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_24 (.CI(n40545), .I0(direction_N_3906), 
            .I1(encoder0_position[22]), .CO(n40546));
    SB_LUT4 position_2066_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[21]), .I3(n40544), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_23 (.CI(n40544), .I0(direction_N_3906), 
            .I1(encoder0_position[21]), .CO(n40545));
    SB_LUT4 position_2066_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[20]), .I3(n40543), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_22 (.CI(n40543), .I0(direction_N_3906), 
            .I1(encoder0_position[20]), .CO(n40544));
    SB_LUT4 position_2066_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[19]), .I3(n40542), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_21 (.CI(n40542), .I0(direction_N_3906), 
            .I1(encoder0_position[19]), .CO(n40543));
    SB_LUT4 position_2066_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[18]), .I3(n40541), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_20 (.CI(n40541), .I0(direction_N_3906), 
            .I1(encoder0_position[18]), .CO(n40542));
    SB_LUT4 position_2066_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[17]), .I3(n40540), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_19 (.CI(n40540), .I0(direction_N_3906), 
            .I1(encoder0_position[17]), .CO(n40541));
    SB_LUT4 position_2066_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[16]), .I3(n40539), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_18 (.CI(n40539), .I0(direction_N_3906), 
            .I1(encoder0_position[16]), .CO(n40540));
    SB_LUT4 position_2066_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[15]), .I3(n40538), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_17 (.CI(n40538), .I0(direction_N_3906), 
            .I1(encoder0_position[15]), .CO(n40539));
    SB_LUT4 position_2066_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[14]), .I3(n40537), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_16 (.CI(n40537), .I0(direction_N_3906), 
            .I1(encoder0_position[14]), .CO(n40538));
    SB_LUT4 position_2066_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[13]), .I3(n40536), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_15 (.CI(n40536), .I0(direction_N_3906), 
            .I1(encoder0_position[13]), .CO(n40537));
    SB_LUT4 position_2066_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[12]), .I3(n40535), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_14 (.CI(n40535), .I0(direction_N_3906), 
            .I1(encoder0_position[12]), .CO(n40536));
    SB_LUT4 position_2066_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[11]), .I3(n40534), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_13 (.CI(n40534), .I0(direction_N_3906), 
            .I1(encoder0_position[11]), .CO(n40535));
    SB_LUT4 position_2066_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[10]), .I3(n40533), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_12 (.CI(n40533), .I0(direction_N_3906), 
            .I1(encoder0_position[10]), .CO(n40534));
    SB_LUT4 position_2066_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[9]), .I3(n40532), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_11 (.CI(n40532), .I0(direction_N_3906), 
            .I1(encoder0_position[9]), .CO(n40533));
    SB_LUT4 position_2066_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[8]), .I3(n40531), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_10 (.CI(n40531), .I0(direction_N_3906), 
            .I1(encoder0_position[8]), .CO(n40532));
    SB_LUT4 position_2066_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[7]), .I3(n40530), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_9 (.CI(n40530), .I0(direction_N_3906), 
            .I1(encoder0_position[7]), .CO(n40531));
    SB_LUT4 position_2066_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[6]), .I3(n40529), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_8 (.CI(n40529), .I0(direction_N_3906), 
            .I1(encoder0_position[6]), .CO(n40530));
    SB_LUT4 position_2066_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[5]), .I3(n40528), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_7 (.CI(n40528), .I0(direction_N_3906), 
            .I1(encoder0_position[5]), .CO(n40529));
    SB_LUT4 position_2066_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[4]), .I3(n40527), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_6 (.CI(n40527), .I0(direction_N_3906), 
            .I1(encoder0_position[4]), .CO(n40528));
    SB_LUT4 position_2066_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[3]), .I3(n40526), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_5 (.CI(n40526), .I0(direction_N_3906), 
            .I1(encoder0_position[3]), .CO(n40527));
    SB_LUT4 position_2066_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[2]), .I3(n40525), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_4 (.CI(n40525), .I0(direction_N_3906), 
            .I1(encoder0_position[2]), .CO(n40526));
    SB_LUT4 position_2066_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[1]), .I3(n40524), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_3 (.CI(n40524), .I0(direction_N_3906), 
            .I1(encoder0_position[1]), .CO(n40525));
    SB_LUT4 position_2066_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2066_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2066_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n40524));
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(\a_new[1] ), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[10] , GND_net, IntegralLimit, \Kp[11] , \Kp[1] , 
            \Kp[0] , \Kp[12] , \Kp[13] , \Kp[14] , \Kp[2] , \Kp[3] , 
            \Kp[15] , \Ki[1] , \Ki[0] , \Kp[4] , \Kp[5] , \Kp[6] , 
            \Kp[7] , \Ki[2] , \Kp[8] , \Ki[3] , \Ki[4] , \Kp[9] , 
            \Ki[5] , \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , 
            \Ki[11] , \Ki[12] , \Ki[13] , PWMLimit, duty, clk32MHz, 
            \Ki[14] , \Ki[15] , VCC_net, setpoint, motor_state) /* synthesis syn_module_defined=1 */ ;
    input \Kp[10] ;
    input GND_net;
    input [23:0]IntegralLimit;
    input \Kp[11] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[15] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Ki[2] ;
    input \Kp[8] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Kp[9] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input [23:0]PWMLimit;
    output [23:0]duty;
    input clk32MHz;
    input \Ki[14] ;
    input \Ki[15] ;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    
    wire n752;
    wire [23:0]n1_adj_4928;
    
    wire n825, \PID_CONTROLLER.integral_23__N_3720 ;
    wire [23:0]n4096;
    
    wire n74, n5;
    wire [16:0]n16459;
    wire [15:0]n17036;
    
    wire n749, n40008, n898, n43, n39323;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n971, n1044, n147, n220, n1117, n17, n9, n11, n49788, 
        n49786, n51835;
    wire [0:0]n10322;
    wire [21:0]n10829;
    
    wire n40155, n50297, n50090, n51817, n50088, n50086, n51810, 
        n27, n15_adj_4510, n13, n11_adj_4511, n50046, n21, n19_adj_4512, 
        n17_adj_4513, n9_adj_4514, n49737, n16_adj_4515, n50026, n8, 
        n45, n24, n7_adj_4516, n5_adj_4517, n49747, n50062, n50058;
    wire [47:0]n106;
    
    wire n40154, n25_adj_4518, n23, n50465, n31, n29, n50383, 
        n37, n35, n33, n50566, n50092, n51804, n50080, n51798, 
        n12, n49760, n51822, n10, n30, n50391, n49769, n51802, 
        n50291, n51828, n50471, n51793, n50568, n51790, n16_adj_4519, 
        n49749, n24_adj_4520, n6_adj_4521, n50481, n50482, n49751, 
        n8_adj_4522, n51788, n50419, n50414;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3723 ;
    
    wire n3_adj_4523, n4_adj_4524, n50447, n50448, n12_adj_4525, n50036, 
        n10_adj_4526, n30_adj_4527, n50038, n50560, n50119, n50598, 
        n50599;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3672 ;
    
    wire n107, n39, n50587, n6_adj_4528, n50475, n50476, n50028, 
        n50423, n38, n50422, n41, n50030, n50543, n50125, n50545, 
        n4_adj_4529, n50479, n50480, n49762, n50558, n50416, n50604, 
        n50605, n50581, n49753, n50501, n40, \PID_CONTROLLER.integral_23__N_3722 , 
        n50503, n39324, n39322, n293, n366, n439, n512, n180, 
        n585, n253, n326, n658, n731, n399, n472, n545, n618, 
        n691, n764, n837, n910, n104, n40153, n35_adj_4535, n177, 
        n250, n40009, n676, n40007, n323, n603, n40006, n396, 
        n469, n542, n615, n688, n761, n834, n907, n980, n122, 
        n53, n195, n268, n341, n414, n487, n560, n101, n804, 
        n32, n877, n475, n402, n40152, n92, n23_adj_4539, n329, 
        n950, n165, n530, n40005, n1023, n174, n238, n256, n1096, 
        n183, n110, n41_adj_4542, n247, n320, n393, n311, n40151, 
        n384, n39321, n466;
    wire [23:0]duty_23__N_3772;
    
    wire n39_adj_4546, n41_adj_4547, n45_adj_4548, n37_adj_4549, n29_adj_4550, 
        n31_adj_4551, n43_adj_4552, n539, n612, n23_adj_4553, n25_adj_4554, 
        n685, n35_adj_4555, n11_adj_4556, n13_adj_4557, n15_adj_4558, 
        n27_adj_4559, n33_adj_4560, n9_adj_4561, n17_adj_4562, n19_adj_4563, 
        n21_adj_4564, n50013, n50006, n12_adj_4565, n10_adj_4566, 
        n30_adj_4567, n50024, n50255, n50251, n40150, n457, n40004;
    wire [23:0]duty_23__N_3648;
    
    wire n758, n50525, n50367, n50564, n40149, n16_adj_4568, n6_adj_4569, 
        n50443, n50444, n40003, n8_adj_4570, n40148, n24_adj_4571, 
        n49989, n39320, n49987, n50425, n50127, n4_adj_4572, n50441, 
        n50442, n40002, n50001, n49997, n50531, n50129, n50600, 
        n50601, n50585, n49991, n50547, n831, n50135, n904, n977, 
        n1050, n39319, n98, n39873;
    wire [10:0]n19011;
    
    wire n50549, n29_adj_4573, duty_23__N_3771;
    wire [23:0]n257;
    
    wire n41_adj_4574, n39_adj_4575, n45_adj_4576;
    wire [9:0]n19252;
    
    wire n39874, n40147, n43_adj_4577, n37_adj_4578, n39875, n40001, 
        n39318, n29_adj_4579, n31_adj_4580, n23_adj_4581, n25_adj_4582, 
        n40146, n35_adj_4583, n33_adj_4584, n11_adj_4585, n13_adj_4586, 
        n15_adj_4587, n27_adj_4589, n40000, n40145, n9_adj_4590, n17_adj_4591, 
        n19_adj_4592, n21_adj_4593, n49975, n49969, n12_adj_4594, 
        n39876, n10_adj_4595, n39877, n30_adj_4596, n39878, n49985, 
        n50209, n50205, n40144, n50519, n171, n50351, n244, n50562, 
        n16_adj_4597, n40143, n6_adj_4598, n50437, n50438, n8_adj_4599, 
        n24_adj_4600, n49954, n49952, n50427, n50137, n4_adj_4601, 
        n50435, n50436, n40142, n49964, n49962, n50533, n50139, 
        n50578, n50579, n50577, n49956, n50551, n50145, n50553, 
        n256_adj_4602;
    wire [23:0]duty_23__N_3747;
    
    wire n40141, n317, n390, n463, n536, n609, n682, n755, n40140, 
        n828, n901, n974, n107_adj_4604, n38_adj_4605, n1047, n1120, 
        n119, n50, n192, n180_adj_4607, n265_adj_4608, n253_adj_4609, 
        n338, n411, n484, n326_adj_4610, n557, n630, n95, n26_adj_4611, 
        n168, n241, n399_adj_4612, n314, n387, n460, n472_adj_4613, 
        n533, n606, n40139, n545_adj_4615, n679, n752_adj_4616, 
        n40138, n39317, n825_adj_4617, n898_adj_4618, n971_adj_4619, 
        n1044_adj_4620, n1117_adj_4621, n618_adj_4622, n92_adj_4623, 
        n23_adj_4624, n86, n17_adj_4626, n165_adj_4627, n238_adj_4628, 
        n311_adj_4629, n384_adj_4630, n457_adj_4631, n530_adj_4632, 
        n603_adj_4633, n39316, n676_adj_4634, n40137, n691_adj_4635, 
        n749_adj_4636, n159, n822, n232, n895, n968, n1041, n39315, 
        n1114, n764_adj_4637, n305, n116, n39314, n47, n40136, 
        n39228;
    wire [14:0]n17547;
    
    wire n39990, n39989, n189, n262_adj_4639, n335, n40135, n39313, 
        n39227, n40134, n408, n39988, n481, n837_adj_4640, n554, 
        n378, n39987, n627, n39226, n700, n89, n20_adj_4641, n162, 
        n235, n39225, n910_adj_4642, n308, n39312, n39986, n451, 
        n381, n524, n454, n39224, n527, n597, n600;
    wire [20:0]n13041;
    
    wire n40133, n39985, n39311, n40132, n39984, n822_adj_4644, 
        n673, n746, n39223, n39310;
    wire [23:0]n1_adj_4929;
    
    wire n819, n892, n670, n965, n39309, n40131, n39308, n679_adj_4651, 
        n39983, n606_adj_4652, n39982, n39307, n40130, n533_adj_4654, 
        n39981, n39306, n39305, n39304, n39303, n40129, n39222, 
        n460_adj_4660, n39980, n1038, n40128, n1111, n387_adj_4661, 
        n39979, n743, n86_adj_4662, n17_adj_4663, n40127, n895_adj_4665, 
        n314_adj_4666, n39978, n241_adj_4668, n39977, n1099, n40126, 
        n1026, n40125, n953, n40124, n880, n40123, n168_adj_4669, 
        n39976, n807, n40122, n734, n40121, n26_adj_4670, n95_adj_4671;
    wire [13:0]n17996;
    
    wire n1120_adj_4672, n39975, n1047_adj_4673, n39974, n974_adj_4674, 
        n39973, n661, n40120, n816, n901_adj_4675, n39972, n159_adj_4676, 
        n39221, n588, n40119, n828_adj_4677, n39971, n755_adj_4679, 
        n39970, n682_adj_4680, n39969, n515, n40118, n609_adj_4682, 
        n39968, n442, n40117, n536_adj_4683, n39967, n369, n40116, 
        n296, n40115, n463_adj_4684, n39966, n232_adj_4685, n305_adj_4686, 
        n390_adj_4688, n39965, n378_adj_4691, n223, n40114, n150_adj_4694, 
        n40113, n968_adj_4695, n317_adj_4698, n39964, n8_adj_4699, 
        n77, n4_adj_4700;
    wire [3:0]n19932;
    
    wire n6_adj_4701, n1041_adj_4703, n244_adj_4705, n39963, n1114_adj_4707;
    wire [19:0]n14291;
    
    wire n40112, n39302, n171_adj_4713, n39962, n29_adj_4715, n98_adj_4716, 
        n40111, n39220, n39301;
    wire [4:0]n19872;
    
    wire n89_adj_4719, n20_adj_4720, n451_adj_4721, n524_adj_4722, n889, 
        n597_adj_4723, n670_adj_4724, n39300;
    wire [12:0]n18387;
    
    wire n1050_adj_4725, n39961, n40110, n977_adj_4726, n39960;
    wire [0:0]n9791;
    wire [21:0]n10298;
    
    wire n39688;
    wire [47:0]n155;
    
    wire n39687, n39686, n162_adj_4727, n904_adj_4728, n39959, n39685, 
        n39299, n39684, n40109, n39219, n235_adj_4730, n39683, n39298, 
        n125, n56, n743_adj_4731, n198, n40108, n816_adj_4732, n889_adj_4733, 
        n39682, n962, n831_adj_4734, n39958, n962_adj_4735, n1035, 
        n1108, n39681, n39297, n40107, n1096_adj_4737, n39680, n271_adj_4738, 
        n308_adj_4739, n344, n1023_adj_4741, n39679, n950_adj_4742, 
        n39678, n113, n44, n186_adj_4743, n259_adj_4744, n332, n417, 
        n405, n478, n877_adj_4745, n39677, n551, n624, n1035_adj_4746, 
        n697, n204, n38911;
    wire [1:0]n19996;
    
    wire n804_adj_4748, n39676, n731_adj_4749, n39675, n658_adj_4750, 
        n39674, n131, n62, n585_adj_4752, n39673, n4_adj_4753;
    wire [2:0]n19972;
    
    wire n490, n12_adj_4754, n8_adj_4755, n11_adj_4756, n6_adj_4757, 
        n38820, n18_adj_4758, n13_adj_4759, n4_adj_4760, n45611, n39296, 
        n770, n83, n14_adj_4761, n758_adj_4762, n39957, n39295, 
        n512_adj_4763, n39672, n1102, n40106, n439_adj_4764, n39671, 
        n685_adj_4765, n39956, n1029, n40105, n612_adj_4766, n39955, 
        n122_adj_4767, n156, n53_adj_4768, n366_adj_4770, n39670, 
        n956, n40104, n229, n302, n539_adj_4771, n39954, n375, 
        n1108_adj_4772, n195_adj_4773, n268_adj_4774, n448, n293_adj_4775, 
        n39669, n883, n40103, n39294, n220_adj_4776, n39668, n381_adj_4777, 
        n521, n147_adj_4778, n39667, n5_adj_4779, n74_adj_4780;
    wire [20:0]n12554;
    
    wire n39666, n39665, n341_adj_4781, n810, n40102, n39293, n466_adj_4782, 
        n39953, n414_adj_4783, n39664, n487_adj_4784, n594, n667, 
        n740, n39663, n560_adj_4785, n454_adj_4786, n39662, n737, 
        n40101, n393_adj_4787, n39952, n119_adj_4788, n39292, n50_adj_4789, 
        n39291, n39661, n39660, n527_adj_4790, n1099_adj_4791, n39659, 
        n192_adj_4792, n1026_adj_4793, n39658, n953_adj_4794, n39657, 
        n265_adj_4795, n338_adj_4796, n39290, n320_adj_4797, n39951, 
        n880_adj_4798, n39656, n807_adj_4799, n39655, n664, n40100, 
        n734_adj_4800, n39654, n39218, n247_adj_4801, n39950, n661_adj_4802, 
        n39653, n411_adj_4803, n591, n40099, n174_adj_4804, n39949, 
        n518, n40098, n600_adj_4805, n588_adj_4806, n39652, n39289, 
        n484_adj_4808, n557_adj_4809, n445, n40097, n813, n886, 
        n959, n1032, n630_adj_4810, n116_adj_4811, n1105, n47_adj_4812, 
        n372, n40096, n299, n40095, n515_adj_4813, n39651, n32_adj_4814, 
        n101_adj_4815, n226, n40094, n442_adj_4816, n39650, n153_adj_4817, 
        n40093;
    wire [11:0]n18724;
    
    wire n980_adj_4818, n39948, n907_adj_4819, n39947, n80, n11_adj_4820, 
        n673_adj_4821, n548, n11_adj_4822, n80_adj_4823;
    wire [18:0]n15091;
    
    wire n40092, n83_adj_4825, n14_adj_4826, n369_adj_4827, n39649, 
        n296_adj_4828, n39648, n223_adj_4829, n39647, n189_adj_4830, 
        n39288, n834_adj_4832, n39946, n40091, n150_adj_4833, n39646, 
        n761_adj_4834, n39945, n688_adj_4835, n39944, n8_adj_4836, 
        n77_adj_4837, n746_adj_4838, n262_adj_4839, n615_adj_4840, n39943;
    wire [19:0]n13851;
    
    wire n39645, n40090, n40089, n542_adj_4841, n39942, n621, n39217, 
        n38836, n335_adj_4842, n819_adj_4843, n39644, n408_adj_4844, 
        n39216, n469_adj_4845, n39941, n153_adj_4846, n39643, n156_adj_4847, 
        n39287, n481_adj_4848, n40088, n39642, n229_adj_4849, n226_adj_4850, 
        n299_adj_4851, n39286, n39641, n302_adj_4852, n1105_adj_4853, 
        n40087, n694, n396_adj_4854, n39940, n39285, n39640, n1102_adj_4855, 
        n39639, n1032_adj_4856, n40086, n892_adj_4857, n1029_adj_4858, 
        n39638, n959_adj_4859, n40085, n375_adj_4860, n448_adj_4861, 
        n372_adj_4862, n521_adj_4863, n445_adj_4864, n594_adj_4865, 
        n554_adj_4866, n667_adj_4867, n767, n740_adj_4868, n38954;
    wire [1:0]n20004;
    
    wire n4_adj_4869, n956_adj_4870, n39637, n518_adj_4871, n627_adj_4872, 
        n323_adj_4873, n39939, n813_adj_4874, n700_adj_4875, n591_adj_4876, 
        n104_adj_4877, n840, n35_adj_4878;
    wire [2:0]n19987;
    
    wire n177_adj_4879, n250_adj_4880, n39938, n883_adj_4881, n39636, 
        n664_adj_4882, n886_adj_4883, n40084, n737_adj_4884, n810_adj_4885, 
        n39635, n39634, n39633, n39215, n39937, n39284, n39632, 
        n40083, n39631, n40082, n40081, n40080, n39630, n40079, 
        n39283, n39629, n40078, n40077, n40076, n39214, n39628, 
        n39627, n38979, n4_adj_4886, n40075, n40074, n39626, n39282;
    wire [17:0]n15812;
    
    wire n40073, n39213;
    wire [18:0]n14692;
    
    wire n39625, n40072, n39212, n39624, n39623, n40071, n39622, 
        n39621;
    wire [3:0]n19956;
    
    wire n39620, n39619, n39618, n39617, n39616, n39615, n39614, 
        n39613, n39612, n40070, n39611, n39211, n40069, n39610, 
        n39609, n39608, n39607;
    wire [8:0]n19451;
    
    wire n39606, n39605, n40068, n39604, n39603, n39602, n39601, 
        n39600, n39599, n39598, n39281, n4_adj_4887, n6_adj_4888;
    wire [17:0]n15452;
    
    wire n39589, n39588, n39587, n39586, n39585, n39584, n39210, 
        n39583, n40067, n39582, n39581, n39580, n39579, n39578;
    wire [4:0]n19907;
    
    wire n40066, n39577, n39576, n39013, n39280, n39209, n39575, 
        n39574, n39573, n39572, n40065, n39208;
    wire [16:0]n16136;
    
    wire n39571, n39570, n39569, n40064, n39568, n39567, n39566, 
        n40063, n39565, n39564, n39207, n39563, n39562, n39561, 
        n40062, n39560, n39559, n40061, n39558, n40060, n39557, 
        n39914, n39556, n39555;
    wire [7:0]n19612;
    
    wire n39554, n39553, n40059, n39206, n39552, n39913, n39551, 
        n39550, n39549, n39548, n39547, n40058;
    wire [15:0]n16748;
    
    wire n39546, n39545, n39912, n39544, n39543, n39542, n39541, 
        n40057, n39205, n39540, n39204, n40056, n39539, n39911, 
        n39538, n39537, n39536, n39535, n39534, n39533, n39532, 
        n39531, n39910;
    wire [14:0]n17292;
    
    wire n39530, n39529, n39528, n39527, n39526, n39525, n39524, 
        n39523, n39909, n39522, n39521, n39908, n39520, n39519, 
        n39518, n39907, n39203, n39517, n39516;
    wire [6:0]n19739;
    
    wire n39515, n39514, n39906, n39513, n39512, n39511, n39905, 
        n39510, n39904, n39509;
    wire [13:0]n17772;
    
    wire n39508, n39202, n39507, n39506, n39505, n39504, n39503, 
        n39201, n39502, n39501, n39500, n39499, n39498, n39497, 
        n39200, n39496, n39495, n39199;
    wire [12:0]n18192;
    
    wire n39494, n39493, n39198, n39492, n39491, n39197, n39490, 
        n39196, n39489, n39195, n39488, n39487, n39194, n39486, 
        n39193, n39485, n39484, n39483, n39482, n39192, n40032, 
        n39191;
    wire [5:0]n19836;
    
    wire n39481, n39480, n39479, n39478, n39477, n39476;
    wire [11:0]n18556;
    
    wire n39475, n39474, n39473, n39472, n39471, n39470, n39469, 
        n39468, n39467, n39466, n39465, n39464;
    wire [10:0]n18868;
    
    wire n39463, n39462, n39461, n39460, n39459, n39458, n39457, 
        n39456, n40031, n39455, n39454, n39453, n39190, n40030, 
        n45940, n490_adj_4889, n39452, n417_adj_4890, n39451, n1111_adj_4891, 
        n40029, n344_adj_4892, n39450, n39189, n271_adj_4893, n39449, 
        n198_adj_4894, n39448, n56_adj_4895, n125_adj_4896;
    wire [9:0]n19132;
    
    wire n840_adj_4897, n39440, n767_adj_4898, n39439, n694_adj_4899, 
        n39438, n621_adj_4900, n39437, n548_adj_4901, n39436, n475_adj_4902, 
        n39435, n402_adj_4903, n39434, n329_adj_4904, n39433, n256_adj_4905, 
        n39432, n183_adj_4906, n39431, n41_adj_4907, n110_adj_4908;
    wire [8:0]n19352;
    
    wire n770_adj_4909, n39417, n697_adj_4910, n39416, n624_adj_4911, 
        n39415, n551_adj_4912, n39414, n478_adj_4913, n39413, n405_adj_4914, 
        n39412, n1038_adj_4915, n40028, n332_adj_4916, n39411, n39188, 
        n259_adj_4917, n39410, n186_adj_4918, n39409, n965_adj_4919, 
        n40027, n44_adj_4920, n113_adj_4921, n39882;
    wire [7:0]n19532;
    
    wire n39408, n39407, n39881, n39406, n40026, n39880, n39187, 
        n39405, n39404, n40025, n39403, n39879, n39186, n39402, 
        n40024, n39401, n40023, n39185;
    wire [6:0]n19676;
    
    wire n39400, n39399, n39398, n40022, n39184, n39397, n39396, 
        n39395, n39394, n40021, n40020;
    wire [5:0]n19788;
    
    wire n39393, n39392, n39391, n39390, n40019, n39183, n39389, 
        n39388, n39387, n39386, n39385, n40018, n39384, n39383, 
        n40017, n40016, n39348, n39347, n39346, n39345, n40015, 
        n39344, n39343, n39342, n39341, n40014, n40013, n39340, 
        n39339, n40012, n39338, n39337, n39336, n40011, n39335, 
        n39334, n39333, n39332, n39331, n39330, n39329, n40010, 
        n39328, n39327, n39326, n39325, n12_adj_4922, n8_adj_4923, 
        n11_adj_4924, n6_adj_4925, n38861, n18_adj_4926, n13_adj_4927;
    
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21883_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21883_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6359_11_lut (.I0(GND_net), .I1(n17036[8]), .I2(n749), 
            .I3(n40008), .O(n16459[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4928[21]), .I3(n39323), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21882_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21882_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21881_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21881_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21880_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21880_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34351_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n49788));
    defparam i34351_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i34349_3_lut (.I0(n11), .I1(n9), .I2(n49788), .I3(GND_net), 
            .O(n49786));
    defparam i34349_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_224_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n51835));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_224_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n10829[21]), .I2(GND_net), 
            .I3(n40155), .O(n10322[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34859_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n51835), 
            .I2(IntegralLimit[7]), .I3(n49786), .O(n50297));
    defparam i34859_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34653_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n50297), .O(n50090));
    defparam i34653_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_206_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n51817));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_206_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34651_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n9), .O(n50088));
    defparam i34651_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34649_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n51817), 
            .I2(IntegralLimit[11]), .I3(n50088), .O(n50086));
    defparam i34649_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_199_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n51810));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_199_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34609_4_lut (.I0(n27), .I1(n15_adj_4510), .I2(n13), .I3(n11_adj_4511), 
            .O(n50046));
    defparam i34609_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34300_4_lut (.I0(n21), .I1(n19_adj_4512), .I2(n17_adj_4513), 
            .I3(n9_adj_4514), .O(n49737));
    defparam i34300_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4515));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34589_2_lut (.I0(n43), .I1(n19_adj_4512), .I2(GND_net), .I3(GND_net), 
            .O(n50026));
    defparam i34589_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4513), .I3(GND_net), 
            .O(n8));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4515), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34310_2_lut (.I0(n7_adj_4516), .I1(n5_adj_4517), .I2(GND_net), 
            .I3(GND_net), .O(n49747));
    defparam i34310_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i34625_4_lut (.I0(n13), .I1(n11_adj_4511), .I2(n9_adj_4514), 
            .I3(n49747), .O(n50062));
    defparam i34625_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34621_4_lut (.I0(n19_adj_4512), .I1(n17_adj_4513), .I2(n15_adj_4510), 
            .I3(n50062), .O(n50058));
    defparam i34621_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n10829[20]), .I2(GND_net), 
            .I3(n40154), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35027_4_lut (.I0(n25_adj_4518), .I1(n23), .I2(n21), .I3(n50058), 
            .O(n50465));
    defparam i35027_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34945_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n50465), 
            .O(n50383));
    defparam i34945_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35128_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n50383), 
            .O(n50566));
    defparam i35128_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34655_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n51835), 
            .I2(IntegralLimit[7]), .I3(n11), .O(n50092));
    defparam i34655_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_193_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n51804));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_193_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34643_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n51804), 
            .I2(IntegralLimit[14]), .I3(n50092), .O(n50080));
    defparam i34643_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_187_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n51798));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_187_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34323_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n49760));
    defparam i34323_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_211_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n51822));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_211_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34953_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n51817), 
            .I2(IntegralLimit[11]), .I3(n50090), .O(n50391));
    defparam i34953_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34332_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n51810), 
            .I2(IntegralLimit[13]), .I3(n50391), .O(n49769));
    defparam i34332_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_191_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n51802));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_191_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34853_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n51802), 
            .I2(IntegralLimit[15]), .I3(n49769), .O(n50291));
    defparam i34853_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_217_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n51828));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_217_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35033_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n51828), 
            .I2(IntegralLimit[17]), .I3(n50291), .O(n50471));
    defparam i35033_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_182_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n51793));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_182_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35130_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n51793), 
            .I2(IntegralLimit[19]), .I3(n50471), .O(n50568));
    defparam i35130_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_179_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n51790));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_179_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4519));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34312_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n49749));
    defparam i34312_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4519), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4520));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4521));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35043_3_lut (.I0(n6_adj_4521), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n50481));   // verilog/motorControl.v(31[10:34])
    defparam i35043_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35044_3_lut (.I0(n50481), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n50482));   // verilog/motorControl.v(31[10:34])
    defparam i35044_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34314_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n51810), 
            .I2(IntegralLimit[21]), .I3(n50086), .O(n49751));
    defparam i34314_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i34981_4_lut (.I0(n24_adj_4520), .I1(n8_adj_4522), .I2(n51788), 
            .I3(n49749), .O(n50419));   // verilog/motorControl.v(31[10:34])
    defparam i34981_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34976_3_lut (.I0(n50482), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n50414));   // verilog/motorControl.v(31[10:34])
    defparam i34976_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3723 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4523), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4524));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i35009_3_lut (.I0(n4_adj_4524), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n50447));   // verilog/motorControl.v(31[38:63])
    defparam i35009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35010_3_lut (.I0(n50447), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n50448));   // verilog/motorControl.v(31[38:63])
    defparam i35010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4525));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34599_2_lut (.I0(n33), .I1(n15_adj_4510), .I2(GND_net), .I3(GND_net), 
            .O(n50036));
    defparam i34599_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13), .I3(GND_net), 
            .O(n10_adj_4526));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4525), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_4527));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34601_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n50046), 
            .O(n50038));
    defparam i34601_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35122_4_lut (.I0(n30_adj_4527), .I1(n10_adj_4526), .I2(n35), 
            .I3(n50036), .O(n50560));   // verilog/motorControl.v(31[38:63])
    defparam i35122_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34682_3_lut (.I0(n50448), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n50119));   // verilog/motorControl.v(31[38:63])
    defparam i34682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35160_4_lut (.I0(n50119), .I1(n50560), .I2(n35), .I3(n50038), 
            .O(n50598));   // verilog/motorControl.v(31[38:63])
    defparam i35160_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35161_3_lut (.I0(n50598), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n50599));   // verilog/motorControl.v(31[38:63])
    defparam i35161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35149_3_lut (.I0(n50599), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n50587));   // verilog/motorControl.v(31[38:63])
    defparam i35149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4516), .I3(GND_net), 
            .O(n6_adj_4528));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35037_3_lut (.I0(n6_adj_4528), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21), .I3(GND_net), .O(n50475));   // verilog/motorControl.v(31[38:63])
    defparam i35037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35038_3_lut (.I0(n50475), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23), .I3(GND_net), .O(n50476));   // verilog/motorControl.v(31[38:63])
    defparam i35038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34591_4_lut (.I0(n43), .I1(n25_adj_4518), .I2(n23), .I3(n49737), 
            .O(n50028));
    defparam i34591_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34985_4_lut (.I0(n24), .I1(n8), .I2(n45), .I3(n50026), 
            .O(n50423));   // verilog/motorControl.v(31[38:63])
    defparam i34985_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34984_3_lut (.I0(n50476), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4518), .I3(GND_net), .O(n50422));   // verilog/motorControl.v(31[38:63])
    defparam i34984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34593_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n50566), 
            .O(n50030));
    defparam i34593_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35105_4_lut (.I0(n50422), .I1(n50423), .I2(n45), .I3(n50028), 
            .O(n50543));   // verilog/motorControl.v(31[38:63])
    defparam i35105_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34688_3_lut (.I0(n50587), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41), .I3(GND_net), .O(n50125));   // verilog/motorControl.v(31[38:63])
    defparam i34688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35107_4_lut (.I0(n50125), .I1(n50543), .I2(n45), .I3(n50030), 
            .O(n50545));   // verilog/motorControl.v(31[38:63])
    defparam i35107_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4529));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i35041_3_lut (.I0(n4_adj_4529), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n50479));   // verilog/motorControl.v(31[10:34])
    defparam i35041_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35042_3_lut (.I0(n50479), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n50480));   // verilog/motorControl.v(31[10:34])
    defparam i35042_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34325_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n51798), 
            .I2(IntegralLimit[16]), .I3(n50080), .O(n49762));
    defparam i34325_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i35120_4_lut (.I0(n30), .I1(n10), .I2(n51822), .I3(n49760), 
            .O(n50558));   // verilog/motorControl.v(31[10:34])
    defparam i35120_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34978_3_lut (.I0(n50480), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n50416));   // verilog/motorControl.v(31[10:34])
    defparam i34978_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35166_4_lut (.I0(n50416), .I1(n50558), .I2(n51822), .I3(n49762), 
            .O(n50604));   // verilog/motorControl.v(31[10:34])
    defparam i35166_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35167_3_lut (.I0(n50604), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n50605));   // verilog/motorControl.v(31[10:34])
    defparam i35167_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35143_3_lut (.I0(n50605), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n50581));   // verilog/motorControl.v(31[10:34])
    defparam i35143_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34316_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n51790), 
            .I2(IntegralLimit[21]), .I3(n50568), .O(n49753));
    defparam i34316_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_177_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n51788));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_177_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35063_4_lut (.I0(n50414), .I1(n50419), .I2(n51788), .I3(n49751), 
            .O(n50501));   // verilog/motorControl.v(31[10:34])
    defparam i35063_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35137_3_lut (.I0(n50581), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[10:34])
    defparam i35137_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35108_3_lut (.I0(n50545), .I1(\PID_CONTROLLER.integral_23__N_3723 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3722 ));   // verilog/motorControl.v(31[38:63])
    defparam i35108_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35065_4_lut (.I0(n40), .I1(n50501), .I2(n51788), .I3(n49753), 
            .O(n50503));   // verilog/motorControl.v(31[10:34])
    defparam i35065_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_850_4_lut  (.I0(n50503), .I1(\PID_CONTROLLER.integral_23__N_3722 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3720 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_850_4_lut .LUT_INIT = 16'h80c8;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n39323), .I0(GND_net), .I1(n1_adj_4928[21]), 
            .CO(n39324));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4928[20]), .I3(n39322), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21879_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21879_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_23 (.CI(n40154), .I0(n10829[20]), .I1(GND_net), 
            .CO(n40155));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n10829[19]), .I2(GND_net), 
            .I3(n40153), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4535));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6359_11 (.CI(n40008), .I0(n17036[8]), .I1(n749), .CO(n40009));
    SB_LUT4 add_6359_10_lut (.I0(GND_net), .I1(n17036[7]), .I2(n676), 
            .I3(n40007), .O(n16459[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6359_10 (.CI(n40007), .I0(n17036[7]), .I1(n676), .CO(n40008));
    SB_LUT4 add_6359_9_lut (.I0(GND_net), .I1(n17036[6]), .I2(n603), .I3(n40006), 
            .O(n16459[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_22 (.CI(n40153), .I0(n10829[19]), .I1(GND_net), 
            .CO(n40154));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n39322), .I0(GND_net), .I1(n1_adj_4928[20]), 
            .CO(n39323));
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n10829[18]), .I2(GND_net), 
            .I3(n40152), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4539));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6359_9 (.CI(n40006), .I0(n17036[6]), .I1(n603), .CO(n40007));
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6359_8_lut (.I0(GND_net), .I1(n17036[5]), .I2(n530), .I3(n40005), 
            .O(n16459[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n40152), .I0(n10829[18]), .I1(GND_net), 
            .CO(n40153));
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4542));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6359_8 (.CI(n40005), .I0(n17036[5]), .I1(n530), .CO(n40006));
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n10829[17]), .I2(GND_net), 
            .I3(n40151), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4928[19]), .I3(n39321), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3772[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4546));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3772[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4547));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3772[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4548));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3772[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4549));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3772[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4550));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3772[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4551));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4552));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3772[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4553));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i23_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_20 (.CI(n40151), .I0(n10829[17]), .I1(GND_net), 
            .CO(n40152));
    SB_LUT4 duty_23__I_851_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3772[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4554));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3772[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4555));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3772[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4556));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3772[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4557));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3772[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4558));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3772[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4559));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4560));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n39321), .I0(GND_net), .I1(n1_adj_4928[19]), 
            .CO(n39322));
    SB_LUT4 duty_23__I_851_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3772[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4561));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3772[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4562));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3772[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4563));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3772[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4564));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34576_4_lut (.I0(n21_adj_4564), .I1(n19_adj_4563), .I2(n17_adj_4562), 
            .I3(n9_adj_4561), .O(n50013));
    defparam i34576_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34569_4_lut (.I0(n27_adj_4559), .I1(n15_adj_4558), .I2(n13_adj_4557), 
            .I3(n11_adj_4556), .O(n50006));
    defparam i34569_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_851_i12_3_lut (.I0(duty_23__N_3772[7]), .I1(duty_23__N_3772[16]), 
            .I2(n33_adj_4560), .I3(GND_net), .O(n12_adj_4565));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i10_3_lut (.I0(duty_23__N_3772[5]), .I1(duty_23__N_3772[6]), 
            .I2(n13_adj_4557), .I3(GND_net), .O(n10_adj_4566));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i30_3_lut (.I0(n12_adj_4565), .I1(duty_23__N_3772[17]), 
            .I2(n35_adj_4555), .I3(GND_net), .O(n30_adj_4567));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34817_4_lut (.I0(n13_adj_4557), .I1(n11_adj_4556), .I2(n9_adj_4561), 
            .I3(n50024), .O(n50255));
    defparam i34817_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34813_4_lut (.I0(n19_adj_4563), .I1(n17_adj_4562), .I2(n15_adj_4558), 
            .I3(n50255), .O(n50251));
    defparam i34813_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n10829[16]), .I2(GND_net), 
            .I3(n40150), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n40150), .I0(n10829[16]), .I1(GND_net), 
            .CO(n40151));
    SB_LUT4 add_6359_7_lut (.I0(GND_net), .I1(n17036[4]), .I2(n457), .I3(n40004), 
            .O(n16459[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3648[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i35087_4_lut (.I0(n25_adj_4554), .I1(n23_adj_4553), .I2(n21_adj_4564), 
            .I3(n50251), .O(n50525));
    defparam i35087_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34929_4_lut (.I0(n31_adj_4551), .I1(n29_adj_4550), .I2(n27_adj_4559), 
            .I3(n50525), .O(n50367));
    defparam i34929_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35126_4_lut (.I0(n37_adj_4549), .I1(n35_adj_4555), .I2(n33_adj_4560), 
            .I3(n50367), .O(n50564));
    defparam i35126_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n10829[15]), .I2(GND_net), 
            .I3(n40149), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n40149), .I0(n10829[15]), .I1(GND_net), 
            .CO(n40150));
    SB_LUT4 duty_23__I_851_i16_3_lut (.I0(duty_23__N_3772[9]), .I1(duty_23__N_3772[21]), 
            .I2(n43_adj_4552), .I3(GND_net), .O(n16_adj_4568));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35005_3_lut (.I0(n6_adj_4569), .I1(duty_23__N_3772[10]), .I2(n21_adj_4564), 
            .I3(GND_net), .O(n50443));   // verilog/motorControl.v(36[10:25])
    defparam i35005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35006_3_lut (.I0(n50443), .I1(duty_23__N_3772[11]), .I2(n23_adj_4553), 
            .I3(GND_net), .O(n50444));   // verilog/motorControl.v(36[10:25])
    defparam i35006_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6359_7 (.CI(n40004), .I0(n17036[4]), .I1(n457), .CO(n40005));
    SB_LUT4 add_6359_6_lut (.I0(GND_net), .I1(n17036[3]), .I2(n384), .I3(n40003), 
            .O(n16459[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i8_3_lut (.I0(duty_23__N_3772[4]), .I1(duty_23__N_3772[8]), 
            .I2(n17_adj_4562), .I3(GND_net), .O(n8_adj_4570));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n10829[14]), .I2(GND_net), 
            .I3(n40148), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i24_3_lut (.I0(n16_adj_4568), .I1(duty_23__N_3772[22]), 
            .I2(n45_adj_4548), .I3(GND_net), .O(n24_adj_4571));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34552_4_lut (.I0(n43_adj_4552), .I1(n25_adj_4554), .I2(n23_adj_4553), 
            .I3(n50013), .O(n49989));
    defparam i34552_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4928[18]), .I3(n39320), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i34987_4_lut (.I0(n24_adj_4571), .I1(n8_adj_4570), .I2(n45_adj_4548), 
            .I3(n49987), .O(n50425));   // verilog/motorControl.v(36[10:25])
    defparam i34987_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34690_3_lut (.I0(n50444), .I1(duty_23__N_3772[12]), .I2(n25_adj_4554), 
            .I3(GND_net), .O(n50127));   // verilog/motorControl.v(36[10:25])
    defparam i34690_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6359_6 (.CI(n40003), .I0(n17036[3]), .I1(n384), .CO(n40004));
    SB_LUT4 duty_23__I_851_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(duty_23__N_3772[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4572));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i35003_3_lut (.I0(n4_adj_4572), .I1(duty_23__N_3772[13]), .I2(n27_adj_4559), 
            .I3(GND_net), .O(n50441));   // verilog/motorControl.v(36[10:25])
    defparam i35003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35004_3_lut (.I0(n50441), .I1(duty_23__N_3772[14]), .I2(n29_adj_4550), 
            .I3(GND_net), .O(n50442));   // verilog/motorControl.v(36[10:25])
    defparam i35004_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n39320), .I0(GND_net), .I1(n1_adj_4928[18]), 
            .CO(n39321));
    SB_LUT4 add_6359_5_lut (.I0(GND_net), .I1(n17036[2]), .I2(n311), .I3(n40002), 
            .O(n16459[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n40148), .I0(n10829[14]), .I1(GND_net), 
            .CO(n40149));
    SB_LUT4 i34564_4_lut (.I0(n33_adj_4560), .I1(n31_adj_4551), .I2(n29_adj_4550), 
            .I3(n50006), .O(n50001));
    defparam i34564_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35093_4_lut (.I0(n30_adj_4567), .I1(n10_adj_4566), .I2(n35_adj_4555), 
            .I3(n49997), .O(n50531));   // verilog/motorControl.v(36[10:25])
    defparam i35093_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34692_3_lut (.I0(n50442), .I1(duty_23__N_3772[15]), .I2(n31_adj_4551), 
            .I3(GND_net), .O(n50129));   // verilog/motorControl.v(36[10:25])
    defparam i34692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35162_4_lut (.I0(n50129), .I1(n50531), .I2(n35_adj_4555), 
            .I3(n50001), .O(n50600));   // verilog/motorControl.v(36[10:25])
    defparam i35162_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35163_3_lut (.I0(n50600), .I1(duty_23__N_3772[18]), .I2(n37_adj_4549), 
            .I3(GND_net), .O(n50601));   // verilog/motorControl.v(36[10:25])
    defparam i35163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35147_3_lut (.I0(n50601), .I1(duty_23__N_3772[19]), .I2(n39_adj_4546), 
            .I3(GND_net), .O(n50585));   // verilog/motorControl.v(36[10:25])
    defparam i35147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34554_4_lut (.I0(n43_adj_4552), .I1(n41_adj_4547), .I2(n39_adj_4546), 
            .I3(n50564), .O(n49991));
    defparam i34554_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_6359_5 (.CI(n40002), .I0(n17036[2]), .I1(n311), .CO(n40003));
    SB_LUT4 i35109_4_lut (.I0(n50127), .I1(n50425), .I2(n45_adj_4548), 
            .I3(n49989), .O(n50547));   // verilog/motorControl.v(36[10:25])
    defparam i35109_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34698_3_lut (.I0(n50585), .I1(duty_23__N_3772[20]), .I2(n41_adj_4547), 
            .I3(GND_net), .O(n50135));   // verilog/motorControl.v(36[10:25])
    defparam i34698_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4928[17]), .I3(n39319), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6521_2 (.CI(GND_net), .I0(n41_adj_4542), .I1(n110), .CO(n39873));
    SB_LUT4 add_6521_2_lut (.I0(GND_net), .I1(n41_adj_4542), .I2(n110), 
            .I3(GND_net), .O(n19011[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35111_4_lut (.I0(n50135), .I1(n50547), .I2(n45_adj_4548), 
            .I3(n49991), .O(n50549));   // verilog/motorControl.v(36[10:25])
    defparam i35111_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4573));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35112_3_lut (.I0(n50549), .I1(PWMLimit[23]), .I2(duty_23__N_3772[23]), 
            .I3(GND_net), .O(duty_23__N_3771));   // verilog/motorControl.v(36[10:25])
    defparam i35112_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n39319), .I0(GND_net), .I1(n1_adj_4928[17]), 
            .CO(n39320));
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4574));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4575));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4576));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6521_3 (.CI(n39873), .I0(n19252[0]), .I1(n183), .CO(n39874));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n10829[13]), .I2(n1096), 
            .I3(n40147), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4577));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4578));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6521_3_lut (.I0(GND_net), .I1(n19252[0]), .I2(n183), .I3(n39873), 
            .O(n19011[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_4 (.CI(n39874), .I0(n19252[1]), .I1(n256), .CO(n39875));
    SB_LUT4 add_6359_4_lut (.I0(GND_net), .I1(n17036[1]), .I2(n238), .I3(n40001), 
            .O(n16459[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4928[16]), .I3(n39318), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4579));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6359_4 (.CI(n40001), .I0(n17036[1]), .I1(n238), .CO(n40002));
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4580));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_16 (.CI(n40147), .I0(n10829[13]), .I1(n1096), 
            .CO(n40148));
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4581));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4582));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n10829[12]), .I2(n1023), 
            .I3(n40146), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_4_lut (.I0(GND_net), .I1(n19252[1]), .I2(n256), .I3(n39874), 
            .O(n19011[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n40146), .I0(n10829[12]), .I1(n1023), 
            .CO(n40147));
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4583));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4584));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4585));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4586));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4587));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4589));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_6359_3_lut (.I0(GND_net), .I1(n17036[0]), .I2(n165), .I3(n40000), 
            .O(n16459[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n10829[11]), .I2(n950), 
            .I3(n40145), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4590));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4591));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_6359_3 (.CI(n40000), .I0(n17036[0]), .I1(n165), .CO(n40001));
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4592));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4593));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34538_4_lut (.I0(n21_adj_4593), .I1(n19_adj_4592), .I2(n17_adj_4591), 
            .I3(n9_adj_4590), .O(n49975));
    defparam i34538_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34532_4_lut (.I0(n27_adj_4589), .I1(n15_adj_4587), .I2(n13_adj_4586), 
            .I3(n11_adj_4585), .O(n49969));
    defparam i34532_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4584), 
            .I3(GND_net), .O(n12_adj_4594));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6521_5 (.CI(n39875), .I0(n19252[2]), .I1(n329), .CO(n39876));
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4586), 
            .I3(GND_net), .O(n10_adj_4595));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6359_2_lut (.I0(GND_net), .I1(n23_adj_4539), .I2(n92), 
            .I3(GND_net), .O(n16459[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6521_5_lut (.I0(GND_net), .I1(n19252[2]), .I2(n329), .I3(n39875), 
            .O(n19011[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_6 (.CI(n39876), .I0(n19252[3]), .I1(n402), .CO(n39877));
    SB_CARRY add_6359_2 (.CI(GND_net), .I0(n23_adj_4539), .I1(n92), .CO(n40000));
    SB_CARRY mult_10_add_1225_14 (.CI(n40145), .I0(n10829[11]), .I1(n950), 
            .CO(n40146));
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4594), .I1(n257[17]), .I2(n35_adj_4583), 
            .I3(GND_net), .O(n30_adj_4596));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6521_7 (.CI(n39877), .I0(n19252[4]), .I1(n475), .CO(n39878));
    SB_LUT4 i34771_4_lut (.I0(n13_adj_4586), .I1(n11_adj_4585), .I2(n9_adj_4590), 
            .I3(n49985), .O(n50209));
    defparam i34771_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34767_4_lut (.I0(n19_adj_4592), .I1(n17_adj_4591), .I2(n15_adj_4587), 
            .I3(n50209), .O(n50205));
    defparam i34767_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n10829[10]), .I2(n877), 
            .I3(n40144), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35081_4_lut (.I0(n25_adj_4582), .I1(n23_adj_4581), .I2(n21_adj_4593), 
            .I3(n50205), .O(n50519));
    defparam i35081_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mult_10_add_1225_13 (.CI(n40144), .I0(n10829[10]), .I1(n877), 
            .CO(n40145));
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34913_4_lut (.I0(n31_adj_4580), .I1(n29_adj_4579), .I2(n27_adj_4589), 
            .I3(n50519), .O(n50351));
    defparam i34913_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35124_4_lut (.I0(n37_adj_4578), .I1(n35_adj_4583), .I2(n33_adj_4584), 
            .I3(n50351), .O(n50562));
    defparam i35124_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4577), 
            .I3(GND_net), .O(n16_adj_4597));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n10829[9]), .I2(n804), 
            .I3(n40143), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34999_3_lut (.I0(n6_adj_4598), .I1(n257[10]), .I2(n21_adj_4593), 
            .I3(GND_net), .O(n50437));   // verilog/motorControl.v(38[19:35])
    defparam i34999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35000_3_lut (.I0(n50437), .I1(n257[11]), .I2(n23_adj_4581), 
            .I3(GND_net), .O(n50438));   // verilog/motorControl.v(38[19:35])
    defparam i35000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4591), 
            .I3(GND_net), .O(n8_adj_4599));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4597), .I1(n257[22]), .I2(n45_adj_4576), 
            .I3(GND_net), .O(n24_adj_4600));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34517_4_lut (.I0(n43_adj_4577), .I1(n25_adj_4582), .I2(n23_adj_4581), 
            .I3(n49975), .O(n49954));
    defparam i34517_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mult_10_add_1225_12 (.CI(n40143), .I0(n10829[9]), .I1(n804), 
            .CO(n40144));
    SB_LUT4 i34989_4_lut (.I0(n24_adj_4600), .I1(n8_adj_4599), .I2(n45_adj_4576), 
            .I3(n49952), .O(n50427));   // verilog/motorControl.v(38[19:35])
    defparam i34989_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34700_3_lut (.I0(n50438), .I1(n257[12]), .I2(n25_adj_4582), 
            .I3(GND_net), .O(n50137));   // verilog/motorControl.v(38[19:35])
    defparam i34700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(n257[1]), 
            .I2(duty_23__N_3772[1]), .I3(n257[0]), .O(n4_adj_4601));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i34997_3_lut (.I0(n4_adj_4601), .I1(n257[13]), .I2(n27_adj_4589), 
            .I3(GND_net), .O(n50435));   // verilog/motorControl.v(38[19:35])
    defparam i34997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34998_3_lut (.I0(n50435), .I1(n257[14]), .I2(n29_adj_4579), 
            .I3(GND_net), .O(n50436));   // verilog/motorControl.v(38[19:35])
    defparam i34998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n10829[8]), .I2(n731), 
            .I3(n40142), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34527_4_lut (.I0(n33_adj_4584), .I1(n31_adj_4580), .I2(n29_adj_4579), 
            .I3(n49969), .O(n49964));
    defparam i34527_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35095_4_lut (.I0(n30_adj_4596), .I1(n10_adj_4595), .I2(n35_adj_4583), 
            .I3(n49962), .O(n50533));   // verilog/motorControl.v(38[19:35])
    defparam i35095_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34702_3_lut (.I0(n50436), .I1(n257[15]), .I2(n31_adj_4580), 
            .I3(GND_net), .O(n50139));   // verilog/motorControl.v(38[19:35])
    defparam i34702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35140_4_lut (.I0(n50139), .I1(n50533), .I2(n35_adj_4583), 
            .I3(n49964), .O(n50578));   // verilog/motorControl.v(38[19:35])
    defparam i35140_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35141_3_lut (.I0(n50578), .I1(n257[18]), .I2(n37_adj_4578), 
            .I3(GND_net), .O(n50579));   // verilog/motorControl.v(38[19:35])
    defparam i35141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35139_3_lut (.I0(n50579), .I1(n257[19]), .I2(n39_adj_4575), 
            .I3(GND_net), .O(n50577));   // verilog/motorControl.v(38[19:35])
    defparam i35139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34519_4_lut (.I0(n43_adj_4577), .I1(n41_adj_4574), .I2(n39_adj_4575), 
            .I3(n50562), .O(n49956));
    defparam i34519_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35113_4_lut (.I0(n50137), .I1(n50427), .I2(n45_adj_4576), 
            .I3(n49954), .O(n50551));   // verilog/motorControl.v(38[19:35])
    defparam i35113_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34708_3_lut (.I0(n50577), .I1(n257[20]), .I2(n41_adj_4574), 
            .I3(GND_net), .O(n50145));   // verilog/motorControl.v(38[19:35])
    defparam i34708_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35115_4_lut (.I0(n50145), .I1(n50551), .I2(n45_adj_4576), 
            .I3(n49956), .O(n50553));   // verilog/motorControl.v(38[19:35])
    defparam i35115_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35116_3_lut (.I0(n50553), .I1(duty_23__N_3772[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4602));   // verilog/motorControl.v(38[19:35])
    defparam i35116_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3772[0]), .I1(n257[0]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3747[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_11 (.CI(n40142), .I0(n10829[8]), .I1(n731), 
            .CO(n40143));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n10829[7]), .I2(n658), 
            .I3(n40141), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_10 (.CI(n40141), .I0(n10829[7]), .I1(n658), 
            .CO(n40142));
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6521_6_lut (.I0(GND_net), .I1(n19252[3]), .I2(n402), .I3(n39876), 
            .O(n19011[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n10829[6]), .I2(n585), 
            .I3(n40140), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4604));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4605));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_9 (.CI(n40140), .I0(n10829[6]), .I1(n585), 
            .CO(n40141));
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4607));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4608));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4609));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_4610));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4611));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_4612));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4613));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n10829[5]), .I2(n512), 
            .I3(n40139), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_1225_8 (.CI(n40139), .I0(n10829[5]), .I1(n512), 
            .CO(n40140));
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4616));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n10829[4]), .I2(n439), 
            .I3(n40138), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n39318), .I0(GND_net), .I1(n1_adj_4928[16]), 
            .CO(n39319));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4928[15]), .I3(n39317), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4617));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4619));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4620));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4622));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_7 (.CI(n40138), .I0(n10829[4]), .I1(n439), 
            .CO(n40139));
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4623));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n39317), .I0(GND_net), .I1(n1_adj_4928[15]), 
            .CO(n39318));
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4626));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4628));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4629));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4631));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4632));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4633));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4928[14]), .I3(n39316), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4634));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n10829[3]), .I2(n366), 
            .I3(n40137), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4635));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4636));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n39316), .I0(GND_net), .I1(n1_adj_4928[14]), 
            .CO(n39317));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4928[13]), .I3(n39315), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_10_add_1225_6 (.CI(n40137), .I0(n10829[3]), .I1(n366), 
            .CO(n40138));
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21721_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21721_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4637));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n39315), .I0(GND_net), .I1(n1_adj_4928[13]), 
            .CO(n39316));
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4928[12]), .I3(n39314), .O(n25_adj_4518)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n10829[2]), .I2(n293), 
            .I3(n40136), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n39314), .I0(GND_net), .I1(n1_adj_4928[12]), 
            .CO(n39315));
    SB_CARRY mult_10_add_1225_5 (.CI(n40136), .I0(n10829[2]), .I1(n293), 
            .CO(n40137));
    SB_LUT4 add_904_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n4096[23]), .I3(n39228), .O(\PID_CONTROLLER.integral_23__N_3672 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_17_lut (.I0(GND_net), .I1(n17547[14]), .I2(GND_net), 
            .I3(n39990), .O(n17036[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_16_lut (.I0(GND_net), .I1(n17547[13]), .I2(n1117), 
            .I3(n39989), .O(n17036[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4639));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n10829[1]), .I2(n220), 
            .I3(n40135), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4928[11]), .I3(n39313), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_10_add_1225_4 (.CI(n40135), .I0(n10829[1]), .I1(n220), 
            .CO(n40136));
    SB_CARRY add_6391_16 (.CI(n39989), .I0(n17547[13]), .I1(n1117), .CO(n39990));
    SB_LUT4 add_904_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n4096[22]), .I3(n39227), .O(\PID_CONTROLLER.integral_23__N_3672 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n10829[0]), .I2(n147), 
            .I3(n40134), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n39313), .I0(GND_net), .I1(n1_adj_4928[11]), 
            .CO(n39314));
    SB_LUT4 add_6391_15_lut (.I0(GND_net), .I1(n17547[12]), .I2(n1044), 
            .I3(n39988), .O(n17036[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_24 (.CI(n39227), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n4096[22]), .CO(n39228));
    SB_CARRY add_6391_15 (.CI(n39988), .I0(n17547[12]), .I1(n1044), .CO(n39989));
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4640));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21903_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21903_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6391_14_lut (.I0(GND_net), .I1(n17547[11]), .I2(n971), 
            .I3(n39987), .O(n17036[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_904_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n4096[21]), .I3(n39226), .O(\PID_CONTROLLER.integral_23__N_3672 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4641));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_904_23 (.CI(n39226), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n4096[21]), .CO(n39227));
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_904_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n4096[20]), .I3(n39225), .O(\PID_CONTROLLER.integral_23__N_3672 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4642));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_3 (.CI(n40134), .I0(n10829[0]), .I1(n147), 
            .CO(n40135));
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4928[10]), .I3(n39312), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6391_14 (.CI(n39987), .I0(n17547[11]), .I1(n971), .CO(n39988));
    SB_CARRY add_904_22 (.CI(n39225), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n4096[20]), .CO(n39226));
    SB_LUT4 add_6391_13_lut (.I0(GND_net), .I1(n17547[10]), .I2(n898), 
            .I3(n39986), .O(n17036[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n39312), .I0(GND_net), .I1(n1_adj_4928[10]), 
            .CO(n39313));
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n40134));
    SB_LUT4 add_904_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n4096[19]), .I3(n39224), .O(\PID_CONTROLLER.integral_23__N_3672 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6391_13 (.CI(n39986), .I0(n17547[10]), .I1(n898), .CO(n39987));
    SB_CARRY add_904_21 (.CI(n39224), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n4096[19]), .CO(n39225));
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4594_23_lut (.I0(GND_net), .I1(n13041[20]), .I2(GND_net), 
            .I3(n40133), .O(n10829[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_12_lut (.I0(GND_net), .I1(n17547[9]), .I2(n825), 
            .I3(n39985), .O(n17036[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4928[9]), .I3(n39311), .O(n19_adj_4512)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6391_12 (.CI(n39985), .I0(n17547[9]), .I1(n825), .CO(n39986));
    SB_LUT4 add_4594_22_lut (.I0(GND_net), .I1(n13041[19]), .I2(GND_net), 
            .I3(n40132), .O(n10829[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n39311), .I0(GND_net), .I1(n1_adj_4928[9]), 
            .CO(n39312));
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6391_11_lut (.I0(GND_net), .I1(n17547[8]), .I2(n752), 
            .I3(n39984), .O(n17036[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4644));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21902_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21902_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_904_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4096[18]), .I3(n39223), .O(\PID_CONTROLLER.integral_23__N_3672 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4928[8]), .I3(n39310), .O(n17_adj_4513)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n39310), .I0(GND_net), .I1(n1_adj_4928[8]), 
            .CO(n39311));
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4928[7]), .I3(n39309), .O(n15_adj_4510)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6391_11 (.CI(n39984), .I0(n17547[8]), .I1(n752), .CO(n39985));
    SB_CARRY add_4594_22 (.CI(n40132), .I0(n13041[19]), .I1(GND_net), 
            .CO(n40133));
    SB_LUT4 add_4594_21_lut (.I0(GND_net), .I1(n13041[18]), .I2(GND_net), 
            .I3(n40131), .O(n10829[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n39309), .I0(GND_net), .I1(n1_adj_4928[7]), 
            .CO(n39310));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4928[6]), .I3(n39308), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6391_10_lut (.I0(GND_net), .I1(n17547[7]), .I2(n679_adj_4651), 
            .I3(n39983), .O(n17036[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_10 (.CI(n39983), .I0(n17547[7]), .I1(n679_adj_4651), 
            .CO(n39984));
    SB_LUT4 add_6391_9_lut (.I0(GND_net), .I1(n17547[6]), .I2(n606_adj_4652), 
            .I3(n39982), .O(n17036[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_21 (.CI(n40131), .I0(n13041[18]), .I1(GND_net), 
            .CO(n40132));
    SB_CARRY add_6391_9 (.CI(n39982), .I0(n17547[6]), .I1(n606_adj_4652), 
            .CO(n39983));
    SB_CARRY unary_minus_5_add_3_8 (.CI(n39308), .I0(GND_net), .I1(n1_adj_4928[6]), 
            .CO(n39309));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4928[5]), .I3(n39307), .O(n11_adj_4511)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n39307), .I0(GND_net), .I1(n1_adj_4928[5]), 
            .CO(n39308));
    SB_CARRY add_904_20 (.CI(n39223), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n4096[18]), .CO(n39224));
    SB_LUT4 add_4594_20_lut (.I0(GND_net), .I1(n13041[17]), .I2(GND_net), 
            .I3(n40130), .O(n10829[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_8_lut (.I0(GND_net), .I1(n17547[5]), .I2(n533_adj_4654), 
            .I3(n39981), .O(n17036[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4928[4]), .I3(n39306), .O(n9_adj_4514)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n39306), .I0(GND_net), .I1(n1_adj_4928[4]), 
            .CO(n39307));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4928[3]), .I3(n39305), .O(n7_adj_4516)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n39305), .I0(GND_net), .I1(n1_adj_4928[3]), 
            .CO(n39306));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4928[2]), .I3(n39304), .O(n5_adj_4517)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n39304), .I0(GND_net), .I1(n1_adj_4928[2]), 
            .CO(n39305));
    SB_CARRY add_6391_8 (.CI(n39981), .I0(n17547[5]), .I1(n533_adj_4654), 
            .CO(n39982));
    SB_CARRY add_4594_20 (.CI(n40130), .I0(n13041[17]), .I1(GND_net), 
            .CO(n40131));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4928[1]), .I3(n39303), .O(n3_adj_4523)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4594_19_lut (.I0(GND_net), .I1(n13041[16]), .I2(GND_net), 
            .I3(n40129), .O(n10829[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n4096[17]), .I3(n39222), .O(\PID_CONTROLLER.integral_23__N_3672 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_19 (.CI(n40129), .I0(n13041[16]), .I1(GND_net), 
            .CO(n40130));
    SB_LUT4 add_6391_7_lut (.I0(GND_net), .I1(n17547[4]), .I2(n460_adj_4660), 
            .I3(n39980), .O(n17036[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n39303), .I0(GND_net), .I1(n1_adj_4928[1]), 
            .CO(n39304));
    SB_LUT4 add_4594_18_lut (.I0(GND_net), .I1(n13041[15]), .I2(GND_net), 
            .I3(n40128), .O(n10829[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_7 (.CI(n39980), .I0(n17547[4]), .I1(n460_adj_4660), 
            .CO(n39981));
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6391_6_lut (.I0(GND_net), .I1(n17547[3]), .I2(n387_adj_4661), 
            .I3(n39979), .O(n17036[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4662));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4663));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4594_18 (.CI(n40128), .I0(n13041[15]), .I1(GND_net), 
            .CO(n40129));
    SB_LUT4 add_4594_17_lut (.I0(GND_net), .I1(n13041[14]), .I2(GND_net), 
            .I3(n40127), .O(n10829[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21901_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21901_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6391_6 (.CI(n39979), .I0(n17547[3]), .I1(n387_adj_4661), 
            .CO(n39980));
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4665));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6391_5_lut (.I0(GND_net), .I1(n17547[2]), .I2(n314_adj_4666), 
            .I3(n39978), .O(n17036[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6391_5 (.CI(n39978), .I0(n17547[2]), .I1(n314_adj_4666), 
            .CO(n39979));
    SB_LUT4 add_6391_4_lut (.I0(GND_net), .I1(n17547[1]), .I2(n241_adj_4668), 
            .I3(n39977), .O(n17036[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_17 (.CI(n40127), .I0(n13041[14]), .I1(GND_net), 
            .CO(n40128));
    SB_LUT4 add_4594_16_lut (.I0(GND_net), .I1(n13041[13]), .I2(n1099), 
            .I3(n40126), .O(n10829[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_16 (.CI(n40126), .I0(n13041[13]), .I1(n1099), .CO(n40127));
    SB_LUT4 add_4594_15_lut (.I0(GND_net), .I1(n13041[12]), .I2(n1026), 
            .I3(n40125), .O(n10829[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_15 (.CI(n40125), .I0(n13041[12]), .I1(n1026), .CO(n40126));
    SB_CARRY add_6391_4 (.CI(n39977), .I0(n17547[1]), .I1(n241_adj_4668), 
            .CO(n39978));
    SB_LUT4 add_4594_14_lut (.I0(GND_net), .I1(n13041[11]), .I2(n953), 
            .I3(n40124), .O(n10829[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_14 (.CI(n40124), .I0(n13041[11]), .I1(n953), .CO(n40125));
    SB_LUT4 add_4594_13_lut (.I0(GND_net), .I1(n13041[10]), .I2(n880), 
            .I3(n40123), .O(n10829[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_13 (.CI(n40123), .I0(n13041[10]), .I1(n880), .CO(n40124));
    SB_LUT4 add_6391_3_lut (.I0(GND_net), .I1(n17547[0]), .I2(n168_adj_4669), 
            .I3(n39976), .O(n17036[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_12_lut (.I0(GND_net), .I1(n13041[9]), .I2(n807), 
            .I3(n40122), .O(n10829[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_3 (.CI(n39976), .I0(n17547[0]), .I1(n168_adj_4669), 
            .CO(n39977));
    SB_CARRY add_4594_12 (.CI(n40122), .I0(n13041[9]), .I1(n807), .CO(n40123));
    SB_LUT4 add_4594_11_lut (.I0(GND_net), .I1(n13041[8]), .I2(n734), 
            .I3(n40121), .O(n10829[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6391_2_lut (.I0(GND_net), .I1(n26_adj_4670), .I2(n95_adj_4671), 
            .I3(GND_net), .O(n17036[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6391_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6391_2 (.CI(GND_net), .I0(n26_adj_4670), .I1(n95_adj_4671), 
            .CO(n39976));
    SB_LUT4 add_6421_16_lut (.I0(GND_net), .I1(n17996[13]), .I2(n1120_adj_4672), 
            .I3(n39975), .O(n17547[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_15_lut (.I0(GND_net), .I1(n17996[12]), .I2(n1047_adj_4673), 
            .I3(n39974), .O(n17547[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_15 (.CI(n39974), .I0(n17996[12]), .I1(n1047_adj_4673), 
            .CO(n39975));
    SB_LUT4 add_6421_14_lut (.I0(GND_net), .I1(n17996[11]), .I2(n974_adj_4674), 
            .I3(n39973), .O(n17547[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_19 (.CI(n39222), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n4096[17]), .CO(n39223));
    SB_CARRY add_6421_14 (.CI(n39973), .I0(n17996[11]), .I1(n974_adj_4674), 
            .CO(n39974));
    SB_CARRY add_4594_11 (.CI(n40121), .I0(n13041[8]), .I1(n734), .CO(n40122));
    SB_LUT4 add_4594_10_lut (.I0(GND_net), .I1(n13041[7]), .I2(n661), 
            .I3(n40120), .O(n10829[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_10 (.CI(n40120), .I0(n13041[7]), .I1(n661), .CO(n40121));
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6421_13_lut (.I0(GND_net), .I1(n17996[10]), .I2(n901_adj_4675), 
            .I3(n39972), .O(n17547[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6421_13 (.CI(n39972), .I0(n17996[10]), .I1(n901_adj_4675), 
            .CO(n39973));
    SB_LUT4 add_904_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n4096[16]), .I3(n39221), .O(\PID_CONTROLLER.integral_23__N_3672 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_9_lut (.I0(GND_net), .I1(n13041[6]), .I2(n588), .I3(n40119), 
            .O(n10829[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_18 (.CI(n39221), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n4096[16]), .CO(n39222));
    SB_LUT4 add_6421_12_lut (.I0(GND_net), .I1(n17996[9]), .I2(n828_adj_4677), 
            .I3(n39971), .O(n17547[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_12 (.CI(n39971), .I0(n17996[9]), .I1(n828_adj_4677), 
            .CO(n39972));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4928[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3723 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_11_lut (.I0(GND_net), .I1(n17996[8]), .I2(n755_adj_4679), 
            .I3(n39970), .O(n17547[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_9 (.CI(n40119), .I0(n13041[6]), .I1(n588), .CO(n40120));
    SB_CARRY add_6421_11 (.CI(n39970), .I0(n17996[8]), .I1(n755_adj_4679), 
            .CO(n39971));
    SB_LUT4 add_6421_10_lut (.I0(GND_net), .I1(n17996[7]), .I2(n682_adj_4680), 
            .I3(n39969), .O(n17547[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_8_lut (.I0(GND_net), .I1(n13041[5]), .I2(n515), .I3(n40118), 
            .O(n10829[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6421_10 (.CI(n39969), .I0(n17996[7]), .I1(n682_adj_4680), 
            .CO(n39970));
    SB_CARRY add_4594_8 (.CI(n40118), .I0(n13041[5]), .I1(n515), .CO(n40119));
    SB_LUT4 add_6421_9_lut (.I0(GND_net), .I1(n17996[6]), .I2(n609_adj_4682), 
            .I3(n39968), .O(n17547[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_9 (.CI(n39968), .I0(n17996[6]), .I1(n609_adj_4682), 
            .CO(n39969));
    SB_LUT4 add_4594_7_lut (.I0(GND_net), .I1(n13041[4]), .I2(n442), .I3(n40117), 
            .O(n10829[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_8_lut (.I0(GND_net), .I1(n17996[5]), .I2(n536_adj_4683), 
            .I3(n39967), .O(n17547[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_7 (.CI(n40117), .I0(n13041[4]), .I1(n442), .CO(n40118));
    SB_LUT4 add_4594_6_lut (.I0(GND_net), .I1(n13041[3]), .I2(n369), .I3(n40116), 
            .O(n10829[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_8 (.CI(n39967), .I0(n17996[5]), .I1(n536_adj_4683), 
            .CO(n39968));
    SB_CARRY add_4594_6 (.CI(n40116), .I0(n13041[3]), .I1(n369), .CO(n40117));
    SB_LUT4 add_4594_5_lut (.I0(GND_net), .I1(n13041[2]), .I2(n296), .I3(n40115), 
            .O(n10829[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6421_7_lut (.I0(GND_net), .I1(n17996[4]), .I2(n463_adj_4684), 
            .I3(n39966), .O(n17547[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_7 (.CI(n39966), .I0(n17996[4]), .I1(n463_adj_4684), 
            .CO(n39967));
    SB_CARRY add_4594_5 (.CI(n40115), .I0(n13041[2]), .I1(n296), .CO(n40116));
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4686));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6421_6_lut (.I0(GND_net), .I1(n17996[3]), .I2(n390_adj_4688), 
            .I3(n39965), .O(n17547[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4594_4_lut (.I0(GND_net), .I1(n13041[1]), .I2(n223), .I3(n40114), 
            .O(n10829[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_4594_4 (.CI(n40114), .I0(n13041[1]), .I1(n223), .CO(n40115));
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6421_6 (.CI(n39965), .I0(n17996[3]), .I1(n390_adj_4688), 
            .CO(n39966));
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_4594_3_lut (.I0(GND_net), .I1(n13041[0]), .I2(n150_adj_4694), 
            .I3(n40113), .O(n10829[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4695));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4594_3 (.CI(n40113), .I0(n13041[0]), .I1(n150_adj_4694), 
            .CO(n40114));
    SB_LUT4 add_6421_5_lut (.I0(GND_net), .I1(n17996[2]), .I2(n317_adj_4698), 
            .I3(n39964), .O(n17547[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_2_lut (.I0(GND_net), .I1(n8_adj_4699), .I2(n77), 
            .I3(GND_net), .O(n10829[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25446_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n4_adj_4700), .I3(n19932[1]), .O(n6_adj_4701));   // verilog/motorControl.v(34[25:36])
    defparam i25446_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6421_5 (.CI(n39964), .I0(n17996[2]), .I1(n317_adj_4698), 
            .CO(n39965));
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4703));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3648[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3648[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3648[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3648[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3648[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3648[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3648[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3648[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3648[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3648[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3648[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3648[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3648[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3648[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3648[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3648[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i21900_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21900_2_lut.LUT_INIT = 16'h8888;
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3648[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4928[0]), 
            .CO(n39303));
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3648[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3648[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3648[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3648[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3648[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3648[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_6421_4_lut (.I0(GND_net), .I1(n17996[1]), .I2(n244_adj_4705), 
            .I3(n39963), .O(n17547[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_2 (.CI(GND_net), .I0(n8_adj_4699), .I1(n77), .CO(n40113));
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4707));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5841_22_lut (.I0(GND_net), .I1(n14291[19]), .I2(GND_net), 
            .I3(n40112), .O(n13041[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n39302), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6421_4 (.CI(n39963), .I0(n17996[1]), .I1(n244_adj_4705), 
            .CO(n39964));
    SB_LUT4 add_6421_3_lut (.I0(GND_net), .I1(n17996[0]), .I2(n171_adj_4713), 
            .I3(n39962), .O(n17547[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6421_3 (.CI(n39962), .I0(n17996[0]), .I1(n171_adj_4713), 
            .CO(n39963));
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6421_2_lut (.I0(GND_net), .I1(n29_adj_4715), .I2(n98_adj_4716), 
            .I3(GND_net), .O(n17547[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6421_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5841_21_lut (.I0(GND_net), .I1(n14291[18]), .I2(GND_net), 
            .I3(n40111), .O(n13041[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n4096[15]), .I3(n39220), .O(\PID_CONTROLLER.integral_23__N_3672 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n39301), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4929[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6421_2 (.CI(GND_net), .I0(n29_adj_4715), .I1(n98_adj_4716), 
            .CO(n39962));
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n19932[1]), .I3(n4_adj_4700), .O(n19872[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_CARRY add_904_17 (.CI(n39220), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n4096[15]), .CO(n39221));
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89_adj_4719));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4720));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4721));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4722));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4723));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_24 (.CI(n39301), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n39302));
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4724));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5841_21 (.CI(n40111), .I0(n14291[18]), .I1(GND_net), 
            .CO(n40112));
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n39300), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_15_lut (.I0(GND_net), .I1(n18387[12]), .I2(n1050_adj_4725), 
            .I3(n39961), .O(n17996[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_20_lut (.I0(GND_net), .I1(n14291[17]), .I2(GND_net), 
            .I3(n40110), .O(n13041[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_14_lut (.I0(GND_net), .I1(n18387[11]), .I2(n977_adj_4726), 
            .I3(n39960), .O(n17996[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I1(n10298[21]), .I2(GND_net), .I3(n39688), .O(n9791[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n10298[20]), .I2(GND_net), 
            .I3(n39687), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n39687), .I0(n10298[20]), .I1(GND_net), 
            .CO(n39688));
    SB_CARRY add_6449_14 (.CI(n39960), .I0(n18387[11]), .I1(n977_adj_4726), 
            .CO(n39961));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n10298[19]), .I2(GND_net), 
            .I3(n39686), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_23 (.CI(n39300), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n39301));
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162_adj_4727));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6449_13_lut (.I0(GND_net), .I1(n18387[10]), .I2(n904_adj_4728), 
            .I3(n39959), .O(n17996[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n39686), .I0(n10298[19]), .I1(GND_net), 
            .CO(n39687));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n10298[18]), .I2(GND_net), 
            .I3(n39685), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_13 (.CI(n39959), .I0(n18387[10]), .I1(n904_adj_4728), 
            .CO(n39960));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n39299), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_20 (.CI(n40110), .I0(n14291[17]), .I1(GND_net), 
            .CO(n40111));
    SB_CARRY mult_11_add_1225_21 (.CI(n39685), .I0(n10298[18]), .I1(GND_net), 
            .CO(n39686));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n10298[17]), .I2(GND_net), 
            .I3(n39684), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_19_lut (.I0(GND_net), .I1(n14291[16]), .I2(GND_net), 
            .I3(n40109), .O(n13041[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_19 (.CI(n40109), .I0(n14291[16]), .I1(GND_net), 
            .CO(n40110));
    SB_CARRY mult_11_add_1225_20 (.CI(n39684), .I0(n10298[17]), .I1(GND_net), 
            .CO(n39685));
    SB_CARRY sub_3_add_2_22 (.CI(n39299), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n39300));
    SB_LUT4 add_904_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n4096[14]), .I3(n39219), .O(\PID_CONTROLLER.integral_23__N_3672 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235_adj_4730));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n10298[16]), .I2(GND_net), 
            .I3(n39683), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n39298), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n39683), .I0(n10298[16]), .I1(GND_net), 
            .CO(n39684));
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5841_18_lut (.I0(GND_net), .I1(n14291[15]), .I2(GND_net), 
            .I3(n40108), .O(n13041[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4732));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4733));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n10298[15]), .I2(GND_net), 
            .I3(n39682), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_18 (.CI(n39682), .I0(n10298[15]), .I1(GND_net), 
            .CO(n39683));
    SB_LUT4 add_6449_12_lut (.I0(GND_net), .I1(n18387[9]), .I2(n831_adj_4734), 
            .I3(n39958), .O(n17996[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_12 (.CI(n39958), .I0(n18387[9]), .I1(n831_adj_4734), 
            .CO(n39959));
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4735));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21897_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21897_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_904_16 (.CI(n39219), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n4096[14]), .CO(n39220));
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n10298[14]), .I2(GND_net), 
            .I3(n39681), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_18 (.CI(n40108), .I0(n14291[15]), .I1(GND_net), 
            .CO(n40109));
    SB_CARRY sub_3_add_2_21 (.CI(n39298), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n39299));
    SB_CARRY mult_11_add_1225_17 (.CI(n39681), .I0(n10298[14]), .I1(GND_net), 
            .CO(n39682));
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n39297), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_17_lut (.I0(GND_net), .I1(n14291[14]), .I2(GND_net), 
            .I3(n40107), .O(n13041[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n39297), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n39298));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n10298[13]), .I2(n1096_adj_4737), 
            .I3(n39680), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4738));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308_adj_4739));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_16 (.CI(n39680), .I0(n10298[13]), .I1(n1096_adj_4737), 
            .CO(n39681));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n10298[12]), .I2(n1023_adj_4741), 
            .I3(n39679), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n39679), .I0(n10298[12]), .I1(n1023_adj_4741), 
            .CO(n39680));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n10298[11]), .I2(n950_adj_4742), 
            .I3(n39678), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_14 (.CI(n39678), .I0(n10298[11]), .I1(n950_adj_4742), 
            .CO(n39679));
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4744));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4701), .I1(\Ki[4] ), .I2(n19932[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), .O(n19872[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n10298[10]), .I2(n877_adj_4745), 
            .I3(n39677), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1519 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n19932[0]), .I3(n38911), .O(n19872[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1519.LUT_INIT = 16'h8778;
    SB_CARRY mult_11_add_1225_13 (.CI(n39677), .I0(n10298[10]), .I1(n877_adj_4745), 
            .CO(n39678));
    SB_LUT4 i25341_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n19996[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25341_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n10298[9]), .I2(n804_adj_4748), 
            .I3(n39676), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n39676), .I0(n10298[9]), .I1(n804_adj_4748), 
            .CO(n39677));
    SB_LUT4 i25438_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n38911), .I3(n19932[0]), .O(n4_adj_4700));   // verilog/motorControl.v(34[25:36])
    defparam i25438_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n10298[8]), .I2(n731_adj_4749), 
            .I3(n39675), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n39675), .I0(n10298[8]), .I1(n731_adj_4749), 
            .CO(n39676));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n10298[7]), .I2(n658_adj_4750), 
            .I3(n39674), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n39674), .I0(n10298[7]), .I1(n658_adj_4750), 
            .CO(n39675));
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n10298[6]), .I2(n585_adj_4752), 
            .I3(n39673), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25425_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n19872[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25425_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i2_4_lut_adj_1520 (.I0(n4_adj_4753), .I1(\Ki[3] ), .I2(n19972[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), .O(n19932[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1520.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1521 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [20]), .O(n12_adj_4754));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1521.LUT_INIT = 16'h9c50;
    SB_LUT4 i25454_4_lut (.I0(n19932[2]), .I1(\Ki[4] ), .I2(n6_adj_4701), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), .O(n8_adj_4755));   // verilog/motorControl.v(34[25:36])
    defparam i25454_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n11_adj_4756));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i25415_4_lut (.I0(n19972[1]), .I1(\Ki[3] ), .I2(n4_adj_4753), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), .O(n6_adj_4757));   // verilog/motorControl.v(34[25:36])
    defparam i25415_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i25343_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n38820));   // verilog/motorControl.v(34[25:36])
    defparam i25343_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4757), .I1(n11_adj_4756), .I2(n8_adj_4755), 
            .I3(n12_adj_4754), .O(n18_adj_4758));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [22]), .O(n13_adj_4759));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4759), .I1(n18_adj_4758), .I2(n38820), 
            .I3(n4_adj_4760), .O(n45611));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25427_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n38911));   // verilog/motorControl.v(34[25:36])
    defparam i25427_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n39296), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_9 (.CI(n39673), .I0(n10298[6]), .I1(n585_adj_4752), 
            .CO(n39674));
    SB_LUT4 add_6449_11_lut (.I0(GND_net), .I1(n18387[8]), .I2(n758_adj_4762), 
            .I3(n39957), .O(n17996[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n39296), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n39297));
    SB_CARRY add_5841_17 (.CI(n40107), .I0(n14291[14]), .I1(GND_net), 
            .CO(n40108));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n39295), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n10298[5]), .I2(n512_adj_4763), 
            .I3(n39672), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n39672), .I0(n10298[5]), .I1(n512_adj_4763), 
            .CO(n39673));
    SB_LUT4 add_5841_16_lut (.I0(GND_net), .I1(n14291[13]), .I2(n1102), 
            .I3(n40106), .O(n13041[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n10298[4]), .I2(n439_adj_4764), 
            .I3(n39671), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_16 (.CI(n40106), .I0(n14291[13]), .I1(n1102), .CO(n40107));
    SB_CARRY add_6449_11 (.CI(n39957), .I0(n18387[8]), .I1(n758_adj_4762), 
            .CO(n39958));
    SB_LUT4 add_6449_10_lut (.I0(GND_net), .I1(n18387[7]), .I2(n685_adj_4765), 
            .I3(n39956), .O(n17996[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_15_lut (.I0(GND_net), .I1(n14291[12]), .I2(n1029), 
            .I3(n40105), .O(n13041[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_15 (.CI(n40105), .I0(n14291[12]), .I1(n1029), .CO(n40106));
    SB_CARRY add_6449_10 (.CI(n39956), .I0(n18387[7]), .I1(n685_adj_4765), 
            .CO(n39957));
    SB_LUT4 add_6449_9_lut (.I0(GND_net), .I1(n18387[6]), .I2(n612_adj_4766), 
            .I3(n39955), .O(n17996[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n39295), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n39296));
    SB_CARRY mult_11_add_1225_7 (.CI(n39671), .I0(n10298[4]), .I1(n439_adj_4764), 
            .CO(n39672));
    SB_CARRY add_6449_9 (.CI(n39955), .I0(n18387[6]), .I1(n612_adj_4766), 
            .CO(n39956));
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4768));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n10298[3]), .I2(n366_adj_4770), 
            .I3(n39670), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_14_lut (.I0(GND_net), .I1(n14291[11]), .I2(n956), 
            .I3(n40104), .O(n13041[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6449_8_lut (.I0(GND_net), .I1(n18387[5]), .I2(n539_adj_4771), 
            .I3(n39954), .O(n17996[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4772));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21896_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21896_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4773));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4774));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_6 (.CI(n39670), .I0(n10298[3]), .I1(n366_adj_4770), 
            .CO(n39671));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n10298[2]), .I2(n293_adj_4775), 
            .I3(n39669), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_14 (.CI(n40104), .I0(n14291[11]), .I1(n956), .CO(n40105));
    SB_LUT4 add_5841_13_lut (.I0(GND_net), .I1(n14291[10]), .I2(n883), 
            .I3(n40103), .O(n13041[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_8 (.CI(n39954), .I0(n18387[5]), .I1(n539_adj_4771), 
            .CO(n39955));
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n39294), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n39669), .I0(n10298[2]), .I1(n293_adj_4775), 
            .CO(n39670));
    SB_CARRY add_5841_13 (.CI(n40103), .I0(n14291[10]), .I1(n883), .CO(n40104));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n10298[1]), .I2(n220_adj_4776), 
            .I3(n39668), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_17 (.CI(n39294), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n39295));
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381_adj_4777));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_4 (.CI(n39668), .I0(n10298[1]), .I1(n220_adj_4776), 
            .CO(n39669));
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n10298[0]), .I2(n147_adj_4778), 
            .I3(n39667), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n39667), .I0(n10298[0]), .I1(n147_adj_4778), 
            .CO(n39668));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4779), .I2(n74_adj_4780), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4779), .I1(n74_adj_4780), 
            .CO(n39667));
    SB_LUT4 add_4571_23_lut (.I0(GND_net), .I1(n12554[20]), .I2(GND_net), 
            .I3(n39666), .O(n10298[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4571_22_lut (.I0(GND_net), .I1(n12554[19]), .I2(GND_net), 
            .I3(n39665), .O(n10298[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4781));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4571_22 (.CI(n39665), .I0(n12554[19]), .I1(GND_net), 
            .CO(n39666));
    SB_LUT4 add_5841_12_lut (.I0(GND_net), .I1(n14291[9]), .I2(n810), 
            .I3(n40102), .O(n13041[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_12 (.CI(n40102), .I0(n14291[9]), .I1(n810), .CO(n40103));
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n39293), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_7_lut (.I0(GND_net), .I1(n18387[4]), .I2(n466_adj_4782), 
            .I3(n39953), .O(n17996[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4783));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4571_21_lut (.I0(GND_net), .I1(n12554[18]), .I2(GND_net), 
            .I3(n39664), .O(n10298[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4784));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4571_21 (.CI(n39664), .I0(n12554[18]), .I1(GND_net), 
            .CO(n39665));
    SB_LUT4 add_4571_20_lut (.I0(GND_net), .I1(n12554[17]), .I2(GND_net), 
            .I3(n39663), .O(n10298[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4785));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454_adj_4786));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_16 (.CI(n39293), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n39294));
    SB_CARRY add_4571_20 (.CI(n39663), .I0(n12554[17]), .I1(GND_net), 
            .CO(n39664));
    SB_LUT4 add_4571_19_lut (.I0(GND_net), .I1(n12554[16]), .I2(GND_net), 
            .I3(n39662), .O(n10298[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_19 (.CI(n39662), .I0(n12554[16]), .I1(GND_net), 
            .CO(n39663));
    SB_CARRY add_6449_7 (.CI(n39953), .I0(n18387[4]), .I1(n466_adj_4782), 
            .CO(n39954));
    SB_LUT4 add_5841_11_lut (.I0(GND_net), .I1(n14291[8]), .I2(n737), 
            .I3(n40101), .O(n13041[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_6_lut (.I0(GND_net), .I1(n18387[3]), .I2(n393_adj_4787), 
            .I3(n39952), .O(n17996[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4788));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n39292), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_11 (.CI(n40101), .I0(n14291[8]), .I1(n737), .CO(n40102));
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4789));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_15 (.CI(n39292), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n39293));
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n39291), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4571_18_lut (.I0(GND_net), .I1(n12554[15]), .I2(GND_net), 
            .I3(n39661), .O(n10298[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_18 (.CI(n39661), .I0(n12554[15]), .I1(GND_net), 
            .CO(n39662));
    SB_LUT4 add_4571_17_lut (.I0(GND_net), .I1(n12554[14]), .I2(GND_net), 
            .I3(n39660), .O(n10298[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527_adj_4790));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4571_17 (.CI(n39660), .I0(n12554[14]), .I1(GND_net), 
            .CO(n39661));
    SB_LUT4 add_4571_16_lut (.I0(GND_net), .I1(n12554[13]), .I2(n1099_adj_4791), 
            .I3(n39659), .O(n10298[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4792));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4571_16 (.CI(n39659), .I0(n12554[13]), .I1(n1099_adj_4791), 
            .CO(n39660));
    SB_LUT4 add_4571_15_lut (.I0(GND_net), .I1(n12554[12]), .I2(n1026_adj_4793), 
            .I3(n39658), .O(n10298[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_15 (.CI(n39658), .I0(n12554[12]), .I1(n1026_adj_4793), 
            .CO(n39659));
    SB_LUT4 add_4571_14_lut (.I0(GND_net), .I1(n12554[11]), .I2(n953_adj_4794), 
            .I3(n39657), .O(n10298[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_14 (.CI(n39657), .I0(n12554[11]), .I1(n953_adj_4794), 
            .CO(n39658));
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4795));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_14 (.CI(n39291), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n39292));
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4796));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6449_6 (.CI(n39952), .I0(n18387[3]), .I1(n393_adj_4787), 
            .CO(n39953));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n39290), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_5_lut (.I0(GND_net), .I1(n18387[2]), .I2(n320_adj_4797), 
            .I3(n39951), .O(n17996[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_13 (.CI(n39290), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n39291));
    SB_LUT4 add_4571_13_lut (.I0(GND_net), .I1(n12554[10]), .I2(n880_adj_4798), 
            .I3(n39656), .O(n10298[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6449_5 (.CI(n39951), .I0(n18387[2]), .I1(n320_adj_4797), 
            .CO(n39952));
    SB_CARRY add_4571_13 (.CI(n39656), .I0(n12554[10]), .I1(n880_adj_4798), 
            .CO(n39657));
    SB_LUT4 add_4571_12_lut (.I0(GND_net), .I1(n12554[9]), .I2(n807_adj_4799), 
            .I3(n39655), .O(n10298[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_12 (.CI(n39655), .I0(n12554[9]), .I1(n807_adj_4799), 
            .CO(n39656));
    SB_LUT4 add_5841_10_lut (.I0(GND_net), .I1(n14291[7]), .I2(n664), 
            .I3(n40100), .O(n13041[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_10 (.CI(n40100), .I0(n14291[7]), .I1(n664), .CO(n40101));
    SB_LUT4 add_4571_11_lut (.I0(GND_net), .I1(n12554[8]), .I2(n734_adj_4800), 
            .I3(n39654), .O(n10298[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_11 (.CI(n39654), .I0(n12554[8]), .I1(n734_adj_4800), 
            .CO(n39655));
    SB_LUT4 add_904_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n4096[13]), .I3(n39218), .O(\PID_CONTROLLER.integral_23__N_3672 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6449_4_lut (.I0(GND_net), .I1(n18387[1]), .I2(n247_adj_4801), 
            .I3(n39950), .O(n17996[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4571_10_lut (.I0(GND_net), .I1(n12554[7]), .I2(n661_adj_4802), 
            .I3(n39653), .O(n10298[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4803));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4571_10 (.CI(n39653), .I0(n12554[7]), .I1(n661_adj_4802), 
            .CO(n39654));
    SB_LUT4 add_5841_9_lut (.I0(GND_net), .I1(n14291[6]), .I2(n591), .I3(n40099), 
            .O(n13041[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_9 (.CI(n40099), .I0(n14291[6]), .I1(n591), .CO(n40100));
    SB_CARRY add_6449_4 (.CI(n39950), .I0(n18387[1]), .I1(n247_adj_4801), 
            .CO(n39951));
    SB_LUT4 add_6449_3_lut (.I0(GND_net), .I1(n18387[0]), .I2(n174_adj_4804), 
            .I3(n39949), .O(n17996[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_8_lut (.I0(GND_net), .I1(n14291[5]), .I2(n518), .I3(n40098), 
            .O(n13041[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_8 (.CI(n40098), .I0(n14291[5]), .I1(n518), .CO(n40099));
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600_adj_4805));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4571_9_lut (.I0(GND_net), .I1(n12554[6]), .I2(n588_adj_4806), 
            .I3(n39652), .O(n10298[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n39289), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4808));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4809));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5841_7_lut (.I0(GND_net), .I1(n14291[4]), .I2(n445), .I3(n40097), 
            .O(n13041[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_12 (.CI(n39289), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n39290));
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5841_7 (.CI(n40097), .I0(n14291[4]), .I1(n445), .CO(n40098));
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4811));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4812));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4571_9 (.CI(n39652), .I0(n12554[6]), .I1(n588_adj_4806), 
            .CO(n39653));
    SB_CARRY add_6449_3 (.CI(n39949), .I0(n18387[0]), .I1(n174_adj_4804), 
            .CO(n39950));
    SB_LUT4 add_5841_6_lut (.I0(GND_net), .I1(n14291[3]), .I2(n372), .I3(n40096), 
            .O(n13041[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21895_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21895_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5841_6 (.CI(n40096), .I0(n14291[3]), .I1(n372), .CO(n40097));
    SB_LUT4 add_5841_5_lut (.I0(GND_net), .I1(n14291[2]), .I2(n299), .I3(n40095), 
            .O(n13041[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4571_8_lut (.I0(GND_net), .I1(n12554[5]), .I2(n515_adj_4813), 
            .I3(n39651), .O(n10298[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_5 (.CI(n40095), .I0(n14291[2]), .I1(n299), .CO(n40096));
    SB_LUT4 add_6449_2_lut (.I0(GND_net), .I1(n32_adj_4814), .I2(n101_adj_4815), 
            .I3(GND_net), .O(n17996[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6449_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_8 (.CI(n39651), .I0(n12554[5]), .I1(n515_adj_4813), 
            .CO(n39652));
    SB_CARRY add_6449_2 (.CI(GND_net), .I0(n32_adj_4814), .I1(n101_adj_4815), 
            .CO(n39949));
    SB_LUT4 add_5841_4_lut (.I0(GND_net), .I1(n14291[1]), .I2(n226), .I3(n40094), 
            .O(n13041[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4571_7_lut (.I0(GND_net), .I1(n12554[4]), .I2(n442_adj_4816), 
            .I3(n39650), .O(n10298[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_4 (.CI(n40094), .I0(n14291[1]), .I1(n226), .CO(n40095));
    SB_LUT4 add_5841_3_lut (.I0(GND_net), .I1(n14291[0]), .I2(n153_adj_4817), 
            .I3(n40093), .O(n13041[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_3 (.CI(n40093), .I0(n14291[0]), .I1(n153_adj_4817), 
            .CO(n40094));
    SB_LUT4 add_6475_14_lut (.I0(GND_net), .I1(n18724[11]), .I2(n980_adj_4818), 
            .I3(n39948), .O(n18387[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_13_lut (.I0(GND_net), .I1(n18724[10]), .I2(n907_adj_4819), 
            .I3(n39947), .O(n18387[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_7 (.CI(n39650), .I0(n12554[4]), .I1(n442_adj_4816), 
            .CO(n39651));
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4820));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673_adj_4821));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6475_13 (.CI(n39947), .I0(n18724[10]), .I1(n907_adj_4819), 
            .CO(n39948));
    SB_LUT4 add_5841_2_lut (.I0(GND_net), .I1(n11_adj_4822), .I2(n80_adj_4823), 
            .I3(GND_net), .O(n13041[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_2 (.CI(GND_net), .I0(n11_adj_4822), .I1(n80_adj_4823), 
            .CO(n40093));
    SB_LUT4 i21894_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21894_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_21_lut (.I0(GND_net), .I1(n15091[18]), .I2(GND_net), 
            .I3(n40092), .O(n14291[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4825));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4826));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4571_6_lut (.I0(GND_net), .I1(n12554[3]), .I2(n369_adj_4827), 
            .I3(n39649), .O(n10298[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_6 (.CI(n39649), .I0(n12554[3]), .I1(n369_adj_4827), 
            .CO(n39650));
    SB_LUT4 add_4571_5_lut (.I0(GND_net), .I1(n12554[2]), .I2(n296_adj_4828), 
            .I3(n39648), .O(n10298[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_5 (.CI(n39648), .I0(n12554[2]), .I1(n296_adj_4828), 
            .CO(n39649));
    SB_LUT4 add_4571_4_lut (.I0(GND_net), .I1(n12554[1]), .I2(n223_adj_4829), 
            .I3(n39647), .O(n10298[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4830));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n39288), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_4 (.CI(n39647), .I0(n12554[1]), .I1(n223_adj_4829), 
            .CO(n39648));
    SB_LUT4 add_6475_12_lut (.I0(GND_net), .I1(n18724[9]), .I2(n834_adj_4832), 
            .I3(n39946), .O(n18387[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_20_lut (.I0(GND_net), .I1(n15091[17]), .I2(GND_net), 
            .I3(n40091), .O(n14291[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_20 (.CI(n40091), .I0(n15091[17]), .I1(GND_net), 
            .CO(n40092));
    SB_LUT4 add_4571_3_lut (.I0(GND_net), .I1(n12554[0]), .I2(n150_adj_4833), 
            .I3(n39646), .O(n10298[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_12 (.CI(n39946), .I0(n18724[9]), .I1(n834_adj_4832), 
            .CO(n39947));
    SB_LUT4 add_6475_11_lut (.I0(GND_net), .I1(n18724[8]), .I2(n761_adj_4834), 
            .I3(n39945), .O(n18387[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_11 (.CI(n39945), .I0(n18724[8]), .I1(n761_adj_4834), 
            .CO(n39946));
    SB_LUT4 add_6475_10_lut (.I0(GND_net), .I1(n18724[7]), .I2(n688_adj_4835), 
            .I3(n39944), .O(n18387[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_3 (.CI(n39646), .I0(n12554[0]), .I1(n150_adj_4833), 
            .CO(n39647));
    SB_CARRY add_6475_10 (.CI(n39944), .I0(n18724[7]), .I1(n688_adj_4835), 
            .CO(n39945));
    SB_LUT4 add_4571_2_lut (.I0(GND_net), .I1(n8_adj_4836), .I2(n77_adj_4837), 
            .I3(GND_net), .O(n10298[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4571_2 (.CI(GND_net), .I0(n8_adj_4836), .I1(n77_adj_4837), 
            .CO(n39646));
    SB_CARRY add_904_15 (.CI(n39218), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n4096[13]), .CO(n39219));
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4838));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4839));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6475_9_lut (.I0(GND_net), .I1(n18724[6]), .I2(n615_adj_4840), 
            .I3(n39943), .O(n18387[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_9 (.CI(n39943), .I0(n18724[6]), .I1(n615_adj_4840), 
            .CO(n39944));
    SB_LUT4 add_5816_22_lut (.I0(GND_net), .I1(n13851[19]), .I2(GND_net), 
            .I3(n39645), .O(n12554[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_19_lut (.I0(GND_net), .I1(n15091[16]), .I2(GND_net), 
            .I3(n40090), .O(n14291[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_19 (.CI(n40090), .I0(n15091[16]), .I1(GND_net), 
            .CO(n40091));
    SB_LUT4 add_6250_18_lut (.I0(GND_net), .I1(n15091[15]), .I2(GND_net), 
            .I3(n40089), .O(n14291[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_8_lut (.I0(GND_net), .I1(n18724[5]), .I2(n542_adj_4841), 
            .I3(n39942), .O(n18387[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_904_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n4096[12]), .I3(n39217), .O(\PID_CONTROLLER.integral_23__N_3672 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_8 (.CI(n39942), .I0(n18724[5]), .I1(n542_adj_4841), 
            .CO(n39943));
    SB_CARRY add_904_14 (.CI(n39217), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n4096[12]), .CO(n39218));
    SB_LUT4 i25369_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n38836), .I3(n19996[0]), .O(n4_adj_4760));   // verilog/motorControl.v(34[25:36])
    defparam i25369_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4842));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_11 (.CI(n39288), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n39289));
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4843));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5816_21_lut (.I0(GND_net), .I1(n13851[18]), .I2(GND_net), 
            .I3(n39644), .O(n12554[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_21 (.CI(n39644), .I0(n13851[18]), .I1(GND_net), 
            .CO(n39645));
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4844));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_904_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n4096[11]), .I3(n39216), .O(\PID_CONTROLLER.integral_23__N_3672 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_7_lut (.I0(GND_net), .I1(n18724[4]), .I2(n469_adj_4845), 
            .I3(n39941), .O(n18387[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4846));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6250_18 (.CI(n40089), .I0(n15091[15]), .I1(GND_net), 
            .CO(n40090));
    SB_LUT4 add_5816_20_lut (.I0(GND_net), .I1(n13851[17]), .I2(GND_net), 
            .I3(n39643), .O(n12554[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4847));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n39287), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4848));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5816_20 (.CI(n39643), .I0(n13851[17]), .I1(GND_net), 
            .CO(n39644));
    SB_LUT4 add_6250_17_lut (.I0(GND_net), .I1(n15091[14]), .I2(GND_net), 
            .I3(n40088), .O(n14291[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5816_19_lut (.I0(GND_net), .I1(n13851[16]), .I2(GND_net), 
            .I3(n39642), .O(n12554[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4849));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4850));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_10 (.CI(n39287), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n39288));
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4851));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21893_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21893_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5816_19 (.CI(n39642), .I0(n13851[16]), .I1(GND_net), 
            .CO(n39643));
    SB_CARRY add_6250_17 (.CI(n40088), .I0(n15091[14]), .I1(GND_net), 
            .CO(n40089));
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n39286), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_7 (.CI(n39941), .I0(n18724[4]), .I1(n469_adj_4845), 
            .CO(n39942));
    SB_LUT4 add_5816_18_lut (.I0(GND_net), .I1(n13851[15]), .I2(GND_net), 
            .I3(n39641), .O(n12554[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4852));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_16_lut (.I0(GND_net), .I1(n15091[13]), .I2(n1105_adj_4853), 
            .I3(n40087), .O(n14291[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_9 (.CI(n39286), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n39287));
    SB_CARRY add_5816_18 (.CI(n39641), .I0(n13851[15]), .I1(GND_net), 
            .CO(n39642));
    SB_LUT4 add_6475_6_lut (.I0(GND_net), .I1(n18724[3]), .I2(n396_adj_4854), 
            .I3(n39940), .O(n18387[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_6 (.CI(n39940), .I0(n18724[3]), .I1(n396_adj_4854), 
            .CO(n39941));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n39285), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5816_17_lut (.I0(GND_net), .I1(n13851[14]), .I2(GND_net), 
            .I3(n39640), .O(n12554[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_16 (.CI(n40087), .I0(n15091[13]), .I1(n1105_adj_4853), 
            .CO(n40088));
    SB_CARRY add_5816_17 (.CI(n39640), .I0(n13851[14]), .I1(GND_net), 
            .CO(n39641));
    SB_LUT4 add_5816_16_lut (.I0(GND_net), .I1(n13851[13]), .I2(n1102_adj_4855), 
            .I3(n39639), .O(n12554[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_15_lut (.I0(GND_net), .I1(n15091[12]), .I2(n1032_adj_4856), 
            .I3(n40086), .O(n14291[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4857));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5816_16 (.CI(n39639), .I0(n13851[13]), .I1(n1102_adj_4855), 
            .CO(n39640));
    SB_LUT4 add_5816_15_lut (.I0(GND_net), .I1(n13851[12]), .I2(n1029_adj_4858), 
            .I3(n39638), .O(n12554[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_15 (.CI(n40086), .I0(n15091[12]), .I1(n1032_adj_4856), 
            .CO(n40087));
    SB_LUT4 add_6250_14_lut (.I0(GND_net), .I1(n15091[11]), .I2(n959_adj_4859), 
            .I3(n40085), .O(n14291[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4860));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448_adj_4861));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4862));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521_adj_4863));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4864));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594_adj_4865));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4866));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667_adj_4867));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740_adj_4868));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5816_15 (.CI(n39638), .I0(n13851[12]), .I1(n1029_adj_4858), 
            .CO(n39639));
    SB_CARRY sub_3_add_2_8 (.CI(n39285), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n39286));
    SB_CARRY add_6250_14 (.CI(n40085), .I0(n15091[11]), .I1(n959_adj_4859), 
            .CO(n40086));
    SB_LUT4 i25477_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n38954), 
            .I3(n20004[0]), .O(n4_adj_4869));   // verilog/motorControl.v(34[16:22])
    defparam i25477_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_5816_14_lut (.I0(GND_net), .I1(n13851[11]), .I2(n956_adj_4870), 
            .I3(n39637), .O(n12554[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4871));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4872));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5816_14 (.CI(n39637), .I0(n13851[11]), .I1(n956_adj_4870), 
            .CO(n39638));
    SB_LUT4 add_6475_5_lut (.I0(GND_net), .I1(n18724[2]), .I2(n323_adj_4873), 
            .I3(n39939), .O(n18387[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1522 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n19996[0]), .I3(n38836), .O(n19972[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1522.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813_adj_4874));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4875));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4876));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4878));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1523 (.I0(\Kp[2] ), .I1(n1[20]), .I2(n20004[0]), 
            .I3(n38954), .O(n19987[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1523.LUT_INIT = 16'h8778;
    SB_LUT4 i25464_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n19987[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25464_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4879));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21892_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21892_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6475_5 (.CI(n39939), .I0(n18724[2]), .I1(n323_adj_4873), 
            .CO(n39940));
    SB_LUT4 add_6475_4_lut (.I0(GND_net), .I1(n18724[1]), .I2(n250_adj_4880), 
            .I3(n39938), .O(n18387[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1524 (.I0(n62), .I1(n131), .I2(n19972[0]), 
            .I3(n204), .O(n19932[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1524.LUT_INIT = 16'h8778;
    SB_LUT4 i25466_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n38954));   // verilog/motorControl.v(34[16:22])
    defparam i25466_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_6475_4 (.CI(n39938), .I0(n18724[1]), .I1(n250_adj_4880), 
            .CO(n39939));
    SB_LUT4 add_5816_13_lut (.I0(GND_net), .I1(n13851[10]), .I2(n883_adj_4881), 
            .I3(n39636), .O(n12554[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4882));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6250_13_lut (.I0(GND_net), .I1(n15091[10]), .I2(n886_adj_4883), 
            .I3(n40084), .O(n14291[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_13 (.CI(n39636), .I0(n13851[10]), .I1(n883_adj_4881), 
            .CO(n39637));
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4884));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5816_12_lut (.I0(GND_net), .I1(n13851[9]), .I2(n810_adj_4885), 
            .I3(n39635), .O(n12554[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_12 (.CI(n39635), .I0(n13851[9]), .I1(n810_adj_4885), 
            .CO(n39636));
    SB_LUT4 add_5816_11_lut (.I0(GND_net), .I1(n13851[8]), .I2(n737_adj_4884), 
            .I3(n39634), .O(n12554[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_11 (.CI(n39634), .I0(n13851[8]), .I1(n737_adj_4884), 
            .CO(n39635));
    SB_LUT4 add_5816_10_lut (.I0(GND_net), .I1(n13851[7]), .I2(n664_adj_4882), 
            .I3(n39633), .O(n12554[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_13 (.CI(n39216), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n4096[11]), .CO(n39217));
    SB_CARRY add_5816_10 (.CI(n39633), .I0(n13851[7]), .I1(n664_adj_4882), 
            .CO(n39634));
    SB_LUT4 add_904_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n4096[10]), .I3(n39215), .O(\PID_CONTROLLER.integral_23__N_3672 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_13 (.CI(n40084), .I0(n15091[10]), .I1(n886_adj_4883), 
            .CO(n40085));
    SB_LUT4 add_6475_3_lut (.I0(GND_net), .I1(n18724[0]), .I2(n177_adj_4879), 
            .I3(n39937), .O(n18387[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_3 (.CI(n39937), .I0(n18724[0]), .I1(n177_adj_4879), 
            .CO(n39938));
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n39284), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6475_2_lut (.I0(GND_net), .I1(n35_adj_4878), .I2(n104_adj_4877), 
            .I3(GND_net), .O(n18387[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6475_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5816_9_lut (.I0(GND_net), .I1(n13851[6]), .I2(n591_adj_4876), 
            .I3(n39632), .O(n12554[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_9 (.CI(n39632), .I0(n13851[6]), .I1(n591_adj_4876), 
            .CO(n39633));
    SB_LUT4 add_6250_12_lut (.I0(GND_net), .I1(n15091[9]), .I2(n813_adj_4874), 
            .I3(n40083), .O(n14291[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_12 (.CI(n40083), .I0(n15091[9]), .I1(n813_adj_4874), 
            .CO(n40084));
    SB_LUT4 add_5816_8_lut (.I0(GND_net), .I1(n13851[5]), .I2(n518_adj_4871), 
            .I3(n39631), .O(n12554[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_8 (.CI(n39631), .I0(n13851[5]), .I1(n518_adj_4871), 
            .CO(n39632));
    SB_LUT4 add_6250_11_lut (.I0(GND_net), .I1(n15091[8]), .I2(n740_adj_4868), 
            .I3(n40082), .O(n14291[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_11 (.CI(n40082), .I0(n15091[8]), .I1(n740_adj_4868), 
            .CO(n40083));
    SB_LUT4 add_6250_10_lut (.I0(GND_net), .I1(n15091[7]), .I2(n667_adj_4867), 
            .I3(n40081), .O(n14291[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6475_2 (.CI(GND_net), .I0(n35_adj_4878), .I1(n104_adj_4877), 
            .CO(n39937));
    SB_CARRY add_6250_10 (.CI(n40081), .I0(n15091[7]), .I1(n667_adj_4867), 
            .CO(n40082));
    SB_LUT4 add_6250_9_lut (.I0(GND_net), .I1(n15091[6]), .I2(n594_adj_4865), 
            .I3(n40080), .O(n14291[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_9 (.CI(n40080), .I0(n15091[6]), .I1(n594_adj_4865), 
            .CO(n40081));
    SB_LUT4 add_5816_7_lut (.I0(GND_net), .I1(n13851[4]), .I2(n445_adj_4864), 
            .I3(n39630), .O(n12554[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_12 (.CI(n39215), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n4096[10]), .CO(n39216));
    SB_LUT4 add_6250_8_lut (.I0(GND_net), .I1(n15091[5]), .I2(n521_adj_4863), 
            .I3(n40079), .O(n14291[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_7 (.CI(n39284), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n39285));
    SB_CARRY add_5816_7 (.CI(n39630), .I0(n13851[4]), .I1(n445_adj_4864), 
            .CO(n39631));
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n39283), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_8 (.CI(n40079), .I0(n15091[5]), .I1(n521_adj_4863), 
            .CO(n40080));
    SB_LUT4 add_5816_6_lut (.I0(GND_net), .I1(n13851[3]), .I2(n372_adj_4862), 
            .I3(n39629), .O(n12554[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_7_lut (.I0(GND_net), .I1(n15091[4]), .I2(n448_adj_4861), 
            .I3(n40078), .O(n14291[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_7 (.CI(n40078), .I0(n15091[4]), .I1(n448_adj_4861), 
            .CO(n40079));
    SB_CARRY add_5816_6 (.CI(n39629), .I0(n13851[3]), .I1(n372_adj_4862), 
            .CO(n39630));
    SB_LUT4 add_6250_6_lut (.I0(GND_net), .I1(n15091[3]), .I2(n375_adj_4860), 
            .I3(n40077), .O(n14291[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_6 (.CI(n40077), .I0(n15091[3]), .I1(n375_adj_4860), 
            .CO(n40078));
    SB_LUT4 add_6250_5_lut (.I0(GND_net), .I1(n15091[2]), .I2(n302_adj_4852), 
            .I3(n40076), .O(n14291[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n4096[9]), .I3(n39214), .O(\PID_CONTROLLER.integral_23__N_3672 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5816_5_lut (.I0(GND_net), .I1(n13851[2]), .I2(n299_adj_4851), 
            .I3(n39628), .O(n12554[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_5 (.CI(n39628), .I0(n13851[2]), .I1(n299_adj_4851), 
            .CO(n39629));
    SB_CARRY add_6250_5 (.CI(n40076), .I0(n15091[2]), .I1(n302_adj_4852), 
            .CO(n40077));
    SB_CARRY add_904_11 (.CI(n39214), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n4096[9]), .CO(n39215));
    SB_LUT4 add_5816_4_lut (.I0(GND_net), .I1(n13851[1]), .I2(n226_adj_4850), 
            .I3(n39627), .O(n12554[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_4 (.CI(n39627), .I0(n13851[1]), .I1(n226_adj_4850), 
            .CO(n39628));
    SB_LUT4 i25500_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n38979), 
            .I3(n19987[0]), .O(n4_adj_4886));   // verilog/motorControl.v(34[16:22])
    defparam i25500_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_6250_4_lut (.I0(GND_net), .I1(n15091[1]), .I2(n229_adj_4849), 
            .I3(n40075), .O(n14291[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_4 (.CI(n40075), .I0(n15091[1]), .I1(n229_adj_4849), 
            .CO(n40076));
    SB_LUT4 add_6250_3_lut (.I0(GND_net), .I1(n15091[0]), .I2(n156_adj_4847), 
            .I3(n40074), .O(n14291[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n39283), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n39284));
    SB_LUT4 add_5816_3_lut (.I0(GND_net), .I1(n13851[0]), .I2(n153_adj_4846), 
            .I3(n39626), .O(n12554[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6250_3 (.CI(n40074), .I0(n15091[0]), .I1(n156_adj_4847), 
            .CO(n40075));
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n39282), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6250_2_lut (.I0(GND_net), .I1(n14_adj_4826), .I2(n83_adj_4825), 
            .I3(GND_net), .O(n14291[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6250_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_3 (.CI(n39626), .I0(n13851[0]), .I1(n153_adj_4846), 
            .CO(n39627));
    SB_CARRY add_6250_2 (.CI(GND_net), .I0(n14_adj_4826), .I1(n83_adj_4825), 
            .CO(n40074));
    SB_LUT4 add_6289_20_lut (.I0(GND_net), .I1(n15812[17]), .I2(GND_net), 
            .I3(n40073), .O(n15091[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n4096[8]), .I3(n39213), .O(\PID_CONTROLLER.integral_23__N_3672 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_10 (.CI(n39213), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n4096[8]), .CO(n39214));
    SB_LUT4 add_5816_2_lut (.I0(GND_net), .I1(n11_adj_4820), .I2(n80), 
            .I3(GND_net), .O(n12554[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5816_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5816_2 (.CI(GND_net), .I0(n11_adj_4820), .I1(n80), .CO(n39626));
    SB_LUT4 add_6230_21_lut (.I0(GND_net), .I1(n14692[18]), .I2(GND_net), 
            .I3(n39625), .O(n13851[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_19_lut (.I0(GND_net), .I1(n15812[16]), .I2(GND_net), 
            .I3(n40072), .O(n15091[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_19 (.CI(n40072), .I0(n15812[16]), .I1(GND_net), 
            .CO(n40073));
    SB_CARRY sub_3_add_2_5 (.CI(n39282), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n39283));
    SB_LUT4 add_904_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n4096[7]), .I3(n39212), .O(\PID_CONTROLLER.integral_23__N_3672 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6230_20_lut (.I0(GND_net), .I1(n14692[17]), .I2(GND_net), 
            .I3(n39624), .O(n13851[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_20 (.CI(n39624), .I0(n14692[17]), .I1(GND_net), 
            .CO(n39625));
    SB_LUT4 add_6230_19_lut (.I0(GND_net), .I1(n14692[16]), .I2(GND_net), 
            .I3(n39623), .O(n13851[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_18_lut (.I0(GND_net), .I1(n15812[15]), .I2(GND_net), 
            .I3(n40071), .O(n15091[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_19 (.CI(n39623), .I0(n14692[16]), .I1(GND_net), 
            .CO(n39624));
    SB_LUT4 add_6230_18_lut (.I0(GND_net), .I1(n14692[15]), .I2(GND_net), 
            .I3(n39622), .O(n13851[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_18 (.CI(n39622), .I0(n14692[15]), .I1(GND_net), 
            .CO(n39623));
    SB_LUT4 add_6230_17_lut (.I0(GND_net), .I1(n14692[14]), .I2(GND_net), 
            .I3(n39621), .O(n13851[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_17 (.CI(n39621), .I0(n14692[14]), .I1(GND_net), 
            .CO(n39622));
    SB_LUT4 i2_3_lut_4_lut_adj_1525 (.I0(\Kp[2] ), .I1(n1[19]), .I2(n19987[0]), 
            .I3(n38979), .O(n19956[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1525.LUT_INIT = 16'h8778;
    SB_LUT4 add_6230_16_lut (.I0(GND_net), .I1(n14692[13]), .I2(n1105), 
            .I3(n39620), .O(n13851[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_16 (.CI(n39620), .I0(n14692[13]), .I1(n1105), .CO(n39621));
    SB_LUT4 add_6230_15_lut (.I0(GND_net), .I1(n14692[12]), .I2(n1032), 
            .I3(n39619), .O(n13851[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_15 (.CI(n39619), .I0(n14692[12]), .I1(n1032), .CO(n39620));
    SB_CARRY add_6289_18 (.CI(n40071), .I0(n15812[15]), .I1(GND_net), 
            .CO(n40072));
    SB_LUT4 add_6230_14_lut (.I0(GND_net), .I1(n14692[11]), .I2(n959), 
            .I3(n39618), .O(n13851[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25487_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n19956[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25487_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_6230_14 (.CI(n39618), .I0(n14692[11]), .I1(n959), .CO(n39619));
    SB_LUT4 add_6230_13_lut (.I0(GND_net), .I1(n14692[10]), .I2(n886), 
            .I3(n39617), .O(n13851[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_13 (.CI(n39617), .I0(n14692[10]), .I1(n886), .CO(n39618));
    SB_LUT4 add_6230_12_lut (.I0(GND_net), .I1(n14692[9]), .I2(n813), 
            .I3(n39616), .O(n13851[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25489_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n38979));   // verilog/motorControl.v(34[16:22])
    defparam i25489_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_6230_12 (.CI(n39616), .I0(n14692[9]), .I1(n813), .CO(n39617));
    SB_LUT4 add_6230_11_lut (.I0(GND_net), .I1(n14692[8]), .I2(n740), 
            .I3(n39615), .O(n13851[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_9 (.CI(n39212), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n4096[7]), .CO(n39213));
    SB_CARRY add_6230_11 (.CI(n39615), .I0(n14692[8]), .I1(n740), .CO(n39616));
    SB_LUT4 add_6230_10_lut (.I0(GND_net), .I1(n14692[7]), .I2(n667), 
            .I3(n39614), .O(n13851[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_10 (.CI(n39614), .I0(n14692[7]), .I1(n667), .CO(n39615));
    SB_LUT4 add_6230_9_lut (.I0(GND_net), .I1(n14692[6]), .I2(n594), .I3(n39613), 
            .O(n13851[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_9 (.CI(n39613), .I0(n14692[6]), .I1(n594), .CO(n39614));
    SB_LUT4 add_6230_8_lut (.I0(GND_net), .I1(n14692[5]), .I2(n521), .I3(n39612), 
            .O(n13851[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_17_lut (.I0(GND_net), .I1(n15812[14]), .I2(GND_net), 
            .I3(n40070), .O(n15091[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_17 (.CI(n40070), .I0(n15812[14]), .I1(GND_net), 
            .CO(n40071));
    SB_CARRY add_6230_8 (.CI(n39612), .I0(n14692[5]), .I1(n521), .CO(n39613));
    SB_LUT4 add_6230_7_lut (.I0(GND_net), .I1(n14692[4]), .I2(n448), .I3(n39611), 
            .O(n13851[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n4096[6]), .I3(n39211), .O(\PID_CONTROLLER.integral_23__N_3672 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_16_lut (.I0(GND_net), .I1(n15812[13]), .I2(n1108_adj_4772), 
            .I3(n40069), .O(n15091[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_7 (.CI(n39611), .I0(n14692[4]), .I1(n448), .CO(n39612));
    SB_LUT4 add_6230_6_lut (.I0(GND_net), .I1(n14692[3]), .I2(n375), .I3(n39610), 
            .O(n13851[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_6 (.CI(n39610), .I0(n14692[3]), .I1(n375), .CO(n39611));
    SB_LUT4 add_6230_5_lut (.I0(GND_net), .I1(n14692[2]), .I2(n302), .I3(n39609), 
            .O(n13851[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_5 (.CI(n39609), .I0(n14692[2]), .I1(n302), .CO(n39610));
    SB_LUT4 add_6230_4_lut (.I0(GND_net), .I1(n14692[1]), .I2(n229), .I3(n39608), 
            .O(n13851[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_8 (.CI(n39211), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n4096[6]), .CO(n39212));
    SB_CARRY add_6230_4 (.CI(n39608), .I0(n14692[1]), .I1(n229), .CO(n39609));
    SB_LUT4 add_6230_3_lut (.I0(GND_net), .I1(n14692[0]), .I2(n156), .I3(n39607), 
            .O(n13851[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_3 (.CI(n39607), .I0(n14692[0]), .I1(n156), .CO(n39608));
    SB_LUT4 add_6230_2_lut (.I0(GND_net), .I1(n14_adj_4761), .I2(n83), 
            .I3(GND_net), .O(n13851[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6230_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6230_2 (.CI(GND_net), .I0(n14_adj_4761), .I1(n83), .CO(n39607));
    SB_LUT4 add_6541_11_lut (.I0(GND_net), .I1(n19451[8]), .I2(n770), 
            .I3(n39606), .O(n19252[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_16 (.CI(n40069), .I0(n15812[13]), .I1(n1108_adj_4772), 
            .CO(n40070));
    SB_LUT4 add_6541_10_lut (.I0(GND_net), .I1(n19451[7]), .I2(n697), 
            .I3(n39605), .O(n19252[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_10 (.CI(n39605), .I0(n19451[7]), .I1(n697), .CO(n39606));
    SB_LUT4 add_6289_15_lut (.I0(GND_net), .I1(n15812[12]), .I2(n1035_adj_4746), 
            .I3(n40068), .O(n15091[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6541_9_lut (.I0(GND_net), .I1(n19451[6]), .I2(n624), .I3(n39604), 
            .O(n19252[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_9 (.CI(n39604), .I0(n19451[6]), .I1(n624), .CO(n39605));
    SB_LUT4 add_6541_8_lut (.I0(GND_net), .I1(n19451[5]), .I2(n551), .I3(n39603), 
            .O(n19252[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_8 (.CI(n39603), .I0(n19451[5]), .I1(n551), .CO(n39604));
    SB_LUT4 add_6541_7_lut (.I0(GND_net), .I1(n19451[4]), .I2(n478), .I3(n39602), 
            .O(n19252[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_7 (.CI(n39602), .I0(n19451[4]), .I1(n478), .CO(n39603));
    SB_LUT4 add_6541_6_lut (.I0(GND_net), .I1(n19451[3]), .I2(n405), .I3(n39601), 
            .O(n19252[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_6 (.CI(n39601), .I0(n19451[3]), .I1(n405), .CO(n39602));
    SB_LUT4 add_6541_5_lut (.I0(GND_net), .I1(n19451[2]), .I2(n332), .I3(n39600), 
            .O(n19252[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_5 (.CI(n39600), .I0(n19451[2]), .I1(n332), .CO(n39601));
    SB_LUT4 add_6541_4_lut (.I0(GND_net), .I1(n19451[1]), .I2(n259_adj_4744), 
            .I3(n39599), .O(n19252[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_4 (.CI(n39599), .I0(n19451[1]), .I1(n259_adj_4744), 
            .CO(n39600));
    SB_LUT4 add_6541_3_lut (.I0(GND_net), .I1(n19451[0]), .I2(n186_adj_4743), 
            .I3(n39598), .O(n19252[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_3 (.CI(n39598), .I0(n19451[0]), .I1(n186_adj_4743), 
            .CO(n39599));
    SB_LUT4 add_6541_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n19252[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6541_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6541_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n39598));
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n39281), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25539_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4887), 
            .I3(n19956[1]), .O(n6_adj_4888));   // verilog/motorControl.v(34[16:22])
    defparam i25539_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_6289_15 (.CI(n40068), .I0(n15812[12]), .I1(n1035_adj_4746), 
            .CO(n40069));
    SB_LUT4 add_6270_20_lut (.I0(GND_net), .I1(n15452[17]), .I2(GND_net), 
            .I3(n39589), .O(n14692[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_19_lut (.I0(GND_net), .I1(n15452[16]), .I2(GND_net), 
            .I3(n39588), .O(n14692[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_19 (.CI(n39588), .I0(n15452[16]), .I1(GND_net), 
            .CO(n39589));
    SB_LUT4 add_6270_18_lut (.I0(GND_net), .I1(n15452[15]), .I2(GND_net), 
            .I3(n39587), .O(n14692[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_18 (.CI(n39587), .I0(n15452[15]), .I1(GND_net), 
            .CO(n39588));
    SB_LUT4 add_6270_17_lut (.I0(GND_net), .I1(n15452[14]), .I2(GND_net), 
            .I3(n39586), .O(n14692[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_17 (.CI(n39586), .I0(n15452[14]), .I1(GND_net), 
            .CO(n39587));
    SB_LUT4 add_6270_16_lut (.I0(GND_net), .I1(n15452[13]), .I2(n1108), 
            .I3(n39585), .O(n14692[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_16 (.CI(n39585), .I0(n15452[13]), .I1(n1108), .CO(n39586));
    SB_LUT4 add_6270_15_lut (.I0(GND_net), .I1(n15452[12]), .I2(n1035), 
            .I3(n39584), .O(n14692[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_15 (.CI(n39584), .I0(n15452[12]), .I1(n1035), .CO(n39585));
    SB_LUT4 add_904_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n4096[5]), .I3(n39210), .O(\PID_CONTROLLER.integral_23__N_3672 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_14_lut (.I0(GND_net), .I1(n15452[11]), .I2(n962_adj_4735), 
            .I3(n39583), .O(n14692[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25407_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n19972[0]), 
            .O(n4_adj_4753));   // verilog/motorControl.v(34[25:36])
    defparam i25407_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_6289_14_lut (.I0(GND_net), .I1(n15812[11]), .I2(n962), 
            .I3(n40067), .O(n15091[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_14 (.CI(n39583), .I0(n15452[11]), .I1(n962_adj_4735), 
            .CO(n39584));
    SB_LUT4 add_6270_13_lut (.I0(GND_net), .I1(n15452[10]), .I2(n889_adj_4733), 
            .I3(n39582), .O(n14692[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_13 (.CI(n39582), .I0(n15452[10]), .I1(n889_adj_4733), 
            .CO(n39583));
    SB_LUT4 add_6270_12_lut (.I0(GND_net), .I1(n15452[9]), .I2(n816_adj_4732), 
            .I3(n39581), .O(n14692[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_12 (.CI(n39581), .I0(n15452[9]), .I1(n816_adj_4732), 
            .CO(n39582));
    SB_LUT4 add_6270_11_lut (.I0(GND_net), .I1(n15452[8]), .I2(n743_adj_4731), 
            .I3(n39580), .O(n14692[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_11 (.CI(n39580), .I0(n15452[8]), .I1(n743_adj_4731), 
            .CO(n39581));
    SB_CARRY add_6289_14 (.CI(n40067), .I0(n15812[11]), .I1(n962), .CO(n40068));
    SB_LUT4 add_6270_10_lut (.I0(GND_net), .I1(n15452[7]), .I2(n670_adj_4724), 
            .I3(n39579), .O(n14692[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_10 (.CI(n39579), .I0(n15452[7]), .I1(n670_adj_4724), 
            .CO(n39580));
    SB_LUT4 add_6270_9_lut (.I0(GND_net), .I1(n15452[6]), .I2(n597_adj_4723), 
            .I3(n39578), .O(n14692[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1526 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n19956[1]), 
            .I3(n4_adj_4887), .O(n19907[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1526.LUT_INIT = 16'h8778;
    SB_LUT4 add_6289_13_lut (.I0(GND_net), .I1(n15812[10]), .I2(n889), 
            .I3(n40066), .O(n15091[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_9 (.CI(n39578), .I0(n15452[6]), .I1(n597_adj_4723), 
            .CO(n39579));
    SB_CARRY add_904_7 (.CI(n39210), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n4096[5]), .CO(n39211));
    SB_LUT4 add_6270_8_lut (.I0(GND_net), .I1(n15452[5]), .I2(n524_adj_4722), 
            .I3(n39577), .O(n14692[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_8 (.CI(n39577), .I0(n15452[5]), .I1(n524_adj_4722), 
            .CO(n39578));
    SB_CARRY add_6289_13 (.CI(n40066), .I0(n15812[10]), .I1(n889), .CO(n40067));
    SB_LUT4 add_6270_7_lut (.I0(GND_net), .I1(n15452[4]), .I2(n451_adj_4721), 
            .I3(n39576), .O(n14692[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_4 (.CI(n39281), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n39282));
    SB_LUT4 i2_3_lut_4_lut_adj_1527 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n19956[0]), 
            .I3(n39013), .O(n19907[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1527.LUT_INIT = 16'h8778;
    SB_LUT4 i25531_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n39013), 
            .I3(n19956[0]), .O(n4_adj_4887));   // verilog/motorControl.v(34[16:22])
    defparam i25531_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_6270_7 (.CI(n39576), .I0(n15452[4]), .I1(n451_adj_4721), 
            .CO(n39577));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n39280), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n4096[4]), .I3(n39209), .O(\PID_CONTROLLER.integral_23__N_3672 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6270_6_lut (.I0(GND_net), .I1(n15452[3]), .I2(n378_adj_4691), 
            .I3(n39575), .O(n14692[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_6 (.CI(n39575), .I0(n15452[3]), .I1(n378_adj_4691), 
            .CO(n39576));
    SB_LUT4 add_6270_5_lut (.I0(GND_net), .I1(n15452[2]), .I2(n305_adj_4686), 
            .I3(n39574), .O(n14692[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_5 (.CI(n39574), .I0(n15452[2]), .I1(n305_adj_4686), 
            .CO(n39575));
    SB_LUT4 add_6270_4_lut (.I0(GND_net), .I1(n15452[1]), .I2(n232_adj_4685), 
            .I3(n39573), .O(n14692[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_4 (.CI(n39573), .I0(n15452[1]), .I1(n232_adj_4685), 
            .CO(n39574));
    SB_CARRY add_904_6 (.CI(n39209), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n4096[4]), .CO(n39210));
    SB_LUT4 add_6270_3_lut (.I0(GND_net), .I1(n15452[0]), .I2(n159_adj_4676), 
            .I3(n39572), .O(n14692[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_12_lut (.I0(GND_net), .I1(n15812[9]), .I2(n816), 
            .I3(n40065), .O(n15091[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n4096[3]), .I3(n39208), .O(\PID_CONTROLLER.integral_23__N_3672 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n39280), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n39281));
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n39280));
    SB_CARRY add_6270_3 (.CI(n39572), .I0(n15452[0]), .I1(n159_adj_4676), 
            .CO(n39573));
    SB_CARRY add_6289_12 (.CI(n40065), .I0(n15812[9]), .I1(n816), .CO(n40066));
    SB_LUT4 add_6270_2_lut (.I0(GND_net), .I1(n17_adj_4663), .I2(n86_adj_4662), 
            .I3(GND_net), .O(n14692[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6270_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6270_2 (.CI(GND_net), .I0(n17_adj_4663), .I1(n86_adj_4662), 
            .CO(n39572));
    SB_LUT4 add_6307_19_lut (.I0(GND_net), .I1(n16136[16]), .I2(GND_net), 
            .I3(n39571), .O(n15452[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_18_lut (.I0(GND_net), .I1(n16136[15]), .I2(GND_net), 
            .I3(n39570), .O(n15452[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_18 (.CI(n39570), .I0(n16136[15]), .I1(GND_net), 
            .CO(n39571));
    SB_LUT4 i25356_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n19972[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25356_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_904_5 (.CI(n39208), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n4096[3]), .CO(n39209));
    SB_LUT4 add_6307_17_lut (.I0(GND_net), .I1(n16136[14]), .I2(GND_net), 
            .I3(n39569), .O(n15452[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_11_lut (.I0(GND_net), .I1(n15812[8]), .I2(n743), 
            .I3(n40064), .O(n15091[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_17 (.CI(n39569), .I0(n16136[14]), .I1(GND_net), 
            .CO(n39570));
    SB_CARRY add_6289_11 (.CI(n40064), .I0(n15812[8]), .I1(n743), .CO(n40065));
    SB_LUT4 add_6307_16_lut (.I0(GND_net), .I1(n16136[13]), .I2(n1111), 
            .I3(n39568), .O(n15452[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_16 (.CI(n39568), .I0(n16136[13]), .I1(n1111), .CO(n39569));
    SB_LUT4 add_6307_15_lut (.I0(GND_net), .I1(n16136[12]), .I2(n1038), 
            .I3(n39567), .O(n15452[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_15 (.CI(n39567), .I0(n16136[12]), .I1(n1038), .CO(n39568));
    SB_LUT4 add_6307_14_lut (.I0(GND_net), .I1(n16136[11]), .I2(n965), 
            .I3(n39566), .O(n15452[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_14 (.CI(n39566), .I0(n16136[11]), .I1(n965), .CO(n39567));
    SB_LUT4 add_6289_10_lut (.I0(GND_net), .I1(n15812[7]), .I2(n670), 
            .I3(n40063), .O(n15091[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_13_lut (.I0(GND_net), .I1(n16136[10]), .I2(n892), 
            .I3(n39565), .O(n15452[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_13 (.CI(n39565), .I0(n16136[10]), .I1(n892), .CO(n39566));
    SB_LUT4 add_6307_12_lut (.I0(GND_net), .I1(n16136[9]), .I2(n819), 
            .I3(n39564), .O(n15452[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n4096[2]), .I3(n39207), .O(\PID_CONTROLLER.integral_23__N_3672 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_904_4 (.CI(n39207), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n4096[2]), .CO(n39208));
    SB_CARRY add_6307_12 (.CI(n39564), .I0(n16136[9]), .I1(n819), .CO(n39565));
    SB_LUT4 add_6307_11_lut (.I0(GND_net), .I1(n16136[8]), .I2(n746), 
            .I3(n39563), .O(n15452[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_11 (.CI(n39563), .I0(n16136[8]), .I1(n746), .CO(n39564));
    SB_LUT4 add_6307_10_lut (.I0(GND_net), .I1(n16136[7]), .I2(n673), 
            .I3(n39562), .O(n15452[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_10 (.CI(n39562), .I0(n16136[7]), .I1(n673), .CO(n39563));
    SB_CARRY add_6289_10 (.CI(n40063), .I0(n15812[7]), .I1(n670), .CO(n40064));
    SB_LUT4 add_6307_9_lut (.I0(GND_net), .I1(n16136[6]), .I2(n600), .I3(n39561), 
            .O(n15452[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_9 (.CI(n39561), .I0(n16136[6]), .I1(n600), .CO(n39562));
    SB_LUT4 add_6289_9_lut (.I0(GND_net), .I1(n15812[6]), .I2(n597), .I3(n40062), 
            .O(n15091[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_8_lut (.I0(GND_net), .I1(n16136[5]), .I2(n527), .I3(n39560), 
            .O(n15452[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_8 (.CI(n39560), .I0(n16136[5]), .I1(n527), .CO(n39561));
    SB_LUT4 add_6307_7_lut (.I0(GND_net), .I1(n16136[4]), .I2(n454), .I3(n39559), 
            .O(n15452[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_9 (.CI(n40062), .I0(n15812[6]), .I1(n597), .CO(n40063));
    SB_CARRY add_6307_7 (.CI(n39559), .I0(n16136[4]), .I1(n454), .CO(n39560));
    SB_LUT4 add_6289_8_lut (.I0(GND_net), .I1(n15812[5]), .I2(n524), .I3(n40061), 
            .O(n15091[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6307_6_lut (.I0(GND_net), .I1(n16136[3]), .I2(n381), .I3(n39558), 
            .O(n15452[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_8 (.CI(n40061), .I0(n15812[5]), .I1(n524), .CO(n40062));
    SB_LUT4 add_6289_7_lut (.I0(GND_net), .I1(n15812[4]), .I2(n451), .I3(n40060), 
            .O(n15091[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25358_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n38836));   // verilog/motorControl.v(34[25:36])
    defparam i25358_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_6307_6 (.CI(n39558), .I0(n16136[3]), .I1(n381), .CO(n39559));
    SB_CARRY add_6289_7 (.CI(n40060), .I0(n15812[4]), .I1(n451), .CO(n40061));
    SB_LUT4 add_6307_5_lut (.I0(GND_net), .I1(n16136[2]), .I2(n308), .I3(n39557), 
            .O(n15452[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_13_lut (.I0(GND_net), .I1(n19011[10]), .I2(n910_adj_4642), 
            .I3(n39914), .O(n18724[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_5 (.CI(n39557), .I0(n16136[2]), .I1(n308), .CO(n39558));
    SB_LUT4 add_6307_4_lut (.I0(GND_net), .I1(n16136[1]), .I2(n235), .I3(n39556), 
            .O(n15452[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_4 (.CI(n39556), .I0(n16136[1]), .I1(n235), .CO(n39557));
    SB_LUT4 add_6307_3_lut (.I0(GND_net), .I1(n16136[0]), .I2(n162), .I3(n39555), 
            .O(n15452[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_3 (.CI(n39555), .I0(n16136[0]), .I1(n162), .CO(n39556));
    SB_LUT4 add_6307_2_lut (.I0(GND_net), .I1(n20_adj_4641), .I2(n89), 
            .I3(GND_net), .O(n15452[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6307_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6307_2 (.CI(GND_net), .I0(n20_adj_4641), .I1(n89), .CO(n39555));
    SB_LUT4 add_6559_10_lut (.I0(GND_net), .I1(n19612[7]), .I2(n700), 
            .I3(n39554), .O(n19451[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6559_9_lut (.I0(GND_net), .I1(n19612[6]), .I2(n627), .I3(n39553), 
            .O(n19451[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_9 (.CI(n39553), .I0(n19612[6]), .I1(n627), .CO(n39554));
    SB_LUT4 add_6289_6_lut (.I0(GND_net), .I1(n15812[3]), .I2(n378), .I3(n40059), 
            .O(n15091[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n4096[1]), .I3(n39206), .O(\PID_CONTROLLER.integral_23__N_3672 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6559_8_lut (.I0(GND_net), .I1(n19612[5]), .I2(n554), .I3(n39552), 
            .O(n19451[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_8 (.CI(n39552), .I0(n19612[5]), .I1(n554), .CO(n39553));
    SB_CARRY add_904_3 (.CI(n39206), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n4096[1]), .CO(n39207));
    SB_LUT4 add_6499_12_lut (.I0(GND_net), .I1(n19011[9]), .I2(n837_adj_4640), 
            .I3(n39913), .O(n18724[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6559_7_lut (.I0(GND_net), .I1(n19612[4]), .I2(n481), .I3(n39551), 
            .O(n19451[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_7 (.CI(n39551), .I0(n19612[4]), .I1(n481), .CO(n39552));
    SB_LUT4 add_6559_6_lut (.I0(GND_net), .I1(n19612[3]), .I2(n408), .I3(n39550), 
            .O(n19451[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_6 (.CI(n39550), .I0(n19612[3]), .I1(n408), .CO(n39551));
    SB_LUT4 add_6559_5_lut (.I0(GND_net), .I1(n19612[2]), .I2(n335), .I3(n39549), 
            .O(n19451[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_5 (.CI(n39549), .I0(n19612[2]), .I1(n335), .CO(n39550));
    SB_LUT4 add_6559_4_lut (.I0(GND_net), .I1(n19612[1]), .I2(n262_adj_4639), 
            .I3(n39548), .O(n19451[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6559_4 (.CI(n39548), .I0(n19612[1]), .I1(n262_adj_4639), 
            .CO(n39549));
    SB_LUT4 i25518_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n19907[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25518_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_6559_3_lut (.I0(GND_net), .I1(n19612[0]), .I2(n189), .I3(n39547), 
            .O(n19451[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_6 (.CI(n40059), .I0(n15812[3]), .I1(n378), .CO(n40060));
    SB_CARRY add_6559_3 (.CI(n39547), .I0(n19612[0]), .I1(n189), .CO(n39548));
    SB_LUT4 add_6559_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n19451[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6559_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6289_5_lut (.I0(GND_net), .I1(n15812[2]), .I2(n305), .I3(n40058), 
            .O(n15091[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_5 (.CI(n40058), .I0(n15812[2]), .I1(n305), .CO(n40059));
    SB_CARRY add_6499_12 (.CI(n39913), .I0(n19011[9]), .I1(n837_adj_4640), 
            .CO(n39914));
    SB_CARRY add_6559_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n39547));
    SB_LUT4 add_6342_18_lut (.I0(GND_net), .I1(n16748[15]), .I2(GND_net), 
            .I3(n39546), .O(n16136[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_17_lut (.I0(GND_net), .I1(n16748[14]), .I2(GND_net), 
            .I3(n39545), .O(n16136[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_11_lut (.I0(GND_net), .I1(n19011[8]), .I2(n764_adj_4637), 
            .I3(n39912), .O(n18724[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_904_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n4096[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3672 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_904_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_17 (.CI(n39545), .I0(n16748[14]), .I1(GND_net), 
            .CO(n39546));
    SB_LUT4 add_6342_16_lut (.I0(GND_net), .I1(n16748[13]), .I2(n1114), 
            .I3(n39544), .O(n16136[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_16 (.CI(n39544), .I0(n16748[13]), .I1(n1114), .CO(n39545));
    SB_LUT4 add_6342_15_lut (.I0(GND_net), .I1(n16748[12]), .I2(n1041), 
            .I3(n39543), .O(n16136[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_15 (.CI(n39543), .I0(n16748[12]), .I1(n1041), .CO(n39544));
    SB_LUT4 add_6342_14_lut (.I0(GND_net), .I1(n16748[11]), .I2(n968), 
            .I3(n39542), .O(n16136[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_14 (.CI(n39542), .I0(n16748[11]), .I1(n968), .CO(n39543));
    SB_LUT4 add_6342_13_lut (.I0(GND_net), .I1(n16748[10]), .I2(n895), 
            .I3(n39541), .O(n16136[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_13 (.CI(n39541), .I0(n16748[10]), .I1(n895), .CO(n39542));
    SB_CARRY add_904_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n4096[0]), .CO(n39206));
    SB_LUT4 add_6289_4_lut (.I0(GND_net), .I1(n15812[1]), .I2(n232), .I3(n40057), 
            .O(n15091[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n10322[0]), .I2(n9791[0]), 
            .I3(n39205), .O(duty_23__N_3772[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25520_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n39013));   // verilog/motorControl.v(34[16:22])
    defparam i25520_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_6289_4 (.CI(n40057), .I0(n15812[1]), .I1(n232), .CO(n40058));
    SB_LUT4 add_6342_12_lut (.I0(GND_net), .I1(n16748[9]), .I2(n822), 
            .I3(n39540), .O(n16136[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_11 (.CI(n39912), .I0(n19011[8]), .I1(n764_adj_4637), 
            .CO(n39913));
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n39204), .O(duty_23__N_3772[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_12 (.CI(n39540), .I0(n16748[9]), .I1(n822), .CO(n39541));
    SB_LUT4 add_6289_3_lut (.I0(GND_net), .I1(n15812[0]), .I2(n159), .I3(n40056), 
            .O(n15091[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_11_lut (.I0(GND_net), .I1(n16748[8]), .I2(n749_adj_4636), 
            .I3(n39539), .O(n16136[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_10_lut (.I0(GND_net), .I1(n19011[7]), .I2(n691_adj_4635), 
            .I3(n39911), .O(n18724[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6289_3 (.CI(n40056), .I0(n15812[0]), .I1(n159), .CO(n40057));
    SB_CARRY add_6342_11 (.CI(n39539), .I0(n16748[8]), .I1(n749_adj_4636), 
            .CO(n39540));
    SB_LUT4 add_6342_10_lut (.I0(GND_net), .I1(n16748[7]), .I2(n676_adj_4634), 
            .I3(n39538), .O(n16136[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_10 (.CI(n39538), .I0(n16748[7]), .I1(n676_adj_4634), 
            .CO(n39539));
    SB_LUT4 add_6342_9_lut (.I0(GND_net), .I1(n16748[6]), .I2(n603_adj_4633), 
            .I3(n39537), .O(n16136[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_9 (.CI(n39537), .I0(n16748[6]), .I1(n603_adj_4633), 
            .CO(n39538));
    SB_LUT4 add_6342_8_lut (.I0(GND_net), .I1(n16748[5]), .I2(n530_adj_4632), 
            .I3(n39536), .O(n16136[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_8 (.CI(n39536), .I0(n16748[5]), .I1(n530_adj_4632), 
            .CO(n39537));
    SB_LUT4 add_6342_7_lut (.I0(GND_net), .I1(n16748[4]), .I2(n457_adj_4631), 
            .I3(n39535), .O(n16136[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_7 (.CI(n39535), .I0(n16748[4]), .I1(n457_adj_4631), 
            .CO(n39536));
    SB_LUT4 add_6342_6_lut (.I0(GND_net), .I1(n16748[3]), .I2(n384_adj_4630), 
            .I3(n39534), .O(n16136[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_6 (.CI(n39534), .I0(n16748[3]), .I1(n384_adj_4630), 
            .CO(n39535));
    SB_LUT4 add_6342_5_lut (.I0(GND_net), .I1(n16748[2]), .I2(n311_adj_4629), 
            .I3(n39533), .O(n16136[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_5 (.CI(n39533), .I0(n16748[2]), .I1(n311_adj_4629), 
            .CO(n39534));
    SB_LUT4 add_6342_4_lut (.I0(GND_net), .I1(n16748[1]), .I2(n238_adj_4628), 
            .I3(n39532), .O(n16136[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4885));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6342_4 (.CI(n39532), .I0(n16748[1]), .I1(n238_adj_4628), 
            .CO(n39533));
    SB_LUT4 add_6342_3_lut (.I0(GND_net), .I1(n16748[0]), .I2(n165_adj_4627), 
            .I3(n39531), .O(n16136[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6342_3 (.CI(n39531), .I0(n16748[0]), .I1(n165_adj_4627), 
            .CO(n39532));
    SB_LUT4 add_6289_2_lut (.I0(GND_net), .I1(n17_adj_4626), .I2(n86), 
            .I3(GND_net), .O(n15091[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6289_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6342_2_lut (.I0(GND_net), .I1(n23_adj_4624), .I2(n92_adj_4623), 
            .I3(GND_net), .O(n16136[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6342_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_10 (.CI(n39911), .I0(n19011[7]), .I1(n691_adj_4635), 
            .CO(n39912));
    SB_CARRY add_6342_2 (.CI(GND_net), .I0(n23_adj_4624), .I1(n92_adj_4623), 
            .CO(n39531));
    SB_LUT4 add_6499_9_lut (.I0(GND_net), .I1(n19011[6]), .I2(n618_adj_4622), 
            .I3(n39910), .O(n18724[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_17_lut (.I0(GND_net), .I1(n17292[14]), .I2(GND_net), 
            .I3(n39530), .O(n16748[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_16_lut (.I0(GND_net), .I1(n17292[13]), .I2(n1117_adj_4621), 
            .I3(n39529), .O(n16748[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_16 (.CI(n39529), .I0(n17292[13]), .I1(n1117_adj_4621), 
            .CO(n39530));
    SB_LUT4 add_6375_15_lut (.I0(GND_net), .I1(n17292[12]), .I2(n1044_adj_4620), 
            .I3(n39528), .O(n16748[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_15 (.CI(n39528), .I0(n17292[12]), .I1(n1044_adj_4620), 
            .CO(n39529));
    SB_LUT4 add_6375_14_lut (.I0(GND_net), .I1(n17292[11]), .I2(n971_adj_4619), 
            .I3(n39527), .O(n16748[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_14 (.CI(n39527), .I0(n17292[11]), .I1(n971_adj_4619), 
            .CO(n39528));
    SB_LUT4 add_6375_13_lut (.I0(GND_net), .I1(n17292[10]), .I2(n898_adj_4618), 
            .I3(n39526), .O(n16748[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_13 (.CI(n39526), .I0(n17292[10]), .I1(n898_adj_4618), 
            .CO(n39527));
    SB_LUT4 add_6375_12_lut (.I0(GND_net), .I1(n17292[9]), .I2(n825_adj_4617), 
            .I3(n39525), .O(n16748[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_12 (.CI(n39525), .I0(n17292[9]), .I1(n825_adj_4617), 
            .CO(n39526));
    SB_LUT4 add_6375_11_lut (.I0(GND_net), .I1(n17292[8]), .I2(n752_adj_4616), 
            .I3(n39524), .O(n16748[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_9 (.CI(n39910), .I0(n19011[6]), .I1(n618_adj_4622), 
            .CO(n39911));
    SB_CARRY add_6289_2 (.CI(GND_net), .I0(n17_adj_4626), .I1(n86), .CO(n40056));
    SB_CARRY add_6375_11 (.CI(n39524), .I0(n17292[8]), .I1(n752_adj_4616), 
            .CO(n39525));
    SB_LUT4 add_6375_10_lut (.I0(GND_net), .I1(n17292[7]), .I2(n679), 
            .I3(n39523), .O(n16748[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_10 (.CI(n39523), .I0(n17292[7]), .I1(n679), .CO(n39524));
    SB_LUT4 add_6499_8_lut (.I0(GND_net), .I1(n19011[5]), .I2(n545_adj_4615), 
            .I3(n39909), .O(n18724[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_9_lut (.I0(GND_net), .I1(n17292[6]), .I2(n606), .I3(n39522), 
            .O(n16748[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_9 (.CI(n39522), .I0(n17292[6]), .I1(n606), .CO(n39523));
    SB_CARRY add_6499_8 (.CI(n39909), .I0(n19011[5]), .I1(n545_adj_4615), 
            .CO(n39910));
    SB_LUT4 add_6375_8_lut (.I0(GND_net), .I1(n17292[5]), .I2(n533), .I3(n39521), 
            .O(n16748[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_8 (.CI(n39521), .I0(n17292[5]), .I1(n533), .CO(n39522));
    SB_LUT4 add_6499_7_lut (.I0(GND_net), .I1(n19011[4]), .I2(n472_adj_4613), 
            .I3(n39908), .O(n18724[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_7_lut (.I0(GND_net), .I1(n17292[4]), .I2(n460), .I3(n39520), 
            .O(n16748[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_24 (.CI(n39204), .I0(n106[22]), .I1(n155[22]), .CO(n39205));
    SB_CARRY add_6375_7 (.CI(n39520), .I0(n17292[4]), .I1(n460), .CO(n39521));
    SB_CARRY add_6499_7 (.CI(n39908), .I0(n19011[4]), .I1(n472_adj_4613), 
            .CO(n39909));
    SB_LUT4 add_6375_6_lut (.I0(GND_net), .I1(n17292[3]), .I2(n387), .I3(n39519), 
            .O(n16748[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_6 (.CI(n39519), .I0(n17292[3]), .I1(n387), .CO(n39520));
    SB_LUT4 add_6375_5_lut (.I0(GND_net), .I1(n17292[2]), .I2(n314), .I3(n39518), 
            .O(n16748[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_6_lut (.I0(GND_net), .I1(n19011[3]), .I2(n399_adj_4612), 
            .I3(n39907), .O(n18724[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_5 (.CI(n39518), .I0(n17292[2]), .I1(n314), .CO(n39519));
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n39203), .O(duty_23__N_3772[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6375_4_lut (.I0(GND_net), .I1(n17292[1]), .I2(n241), .I3(n39517), 
            .O(n16748[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_6 (.CI(n39907), .I0(n19011[3]), .I1(n399_adj_4612), 
            .CO(n39908));
    SB_CARRY add_6375_4 (.CI(n39517), .I0(n17292[1]), .I1(n241), .CO(n39518));
    SB_LUT4 add_6375_3_lut (.I0(GND_net), .I1(n17292[0]), .I2(n168), .I3(n39516), 
            .O(n16748[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_3 (.CI(n39516), .I0(n17292[0]), .I1(n168), .CO(n39517));
    SB_LUT4 add_6375_2_lut (.I0(GND_net), .I1(n26_adj_4611), .I2(n95), 
            .I3(GND_net), .O(n16748[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6375_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6375_2 (.CI(GND_net), .I0(n26_adj_4611), .I1(n95), .CO(n39516));
    SB_LUT4 add_6575_9_lut (.I0(GND_net), .I1(n19739[6]), .I2(n630), .I3(n39515), 
            .O(n19612[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6575_8_lut (.I0(GND_net), .I1(n19739[5]), .I2(n557), .I3(n39514), 
            .O(n19612[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_5_lut (.I0(GND_net), .I1(n19011[2]), .I2(n326_adj_4610), 
            .I3(n39906), .O(n18724[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_5 (.CI(n39906), .I0(n19011[2]), .I1(n326_adj_4610), 
            .CO(n39907));
    SB_CARRY add_6575_8 (.CI(n39514), .I0(n19739[5]), .I1(n557), .CO(n39515));
    SB_LUT4 add_6575_7_lut (.I0(GND_net), .I1(n19739[4]), .I2(n484), .I3(n39513), 
            .O(n19612[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6575_7 (.CI(n39513), .I0(n19739[4]), .I1(n484), .CO(n39514));
    SB_LUT4 add_6575_6_lut (.I0(GND_net), .I1(n19739[3]), .I2(n411), .I3(n39512), 
            .O(n19612[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6575_6 (.CI(n39512), .I0(n19739[3]), .I1(n411), .CO(n39513));
    SB_LUT4 add_6575_5_lut (.I0(GND_net), .I1(n19739[2]), .I2(n338), .I3(n39511), 
            .O(n19612[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_4_lut (.I0(GND_net), .I1(n19011[1]), .I2(n253_adj_4609), 
            .I3(n39905), .O(n18724[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_4 (.CI(n39905), .I0(n19011[1]), .I1(n253_adj_4609), 
            .CO(n39906));
    SB_CARRY add_12_23 (.CI(n39203), .I0(n106[21]), .I1(n155[21]), .CO(n39204));
    SB_CARRY add_6575_5 (.CI(n39511), .I0(n19739[2]), .I1(n338), .CO(n39512));
    SB_LUT4 add_6575_4_lut (.I0(GND_net), .I1(n19739[1]), .I2(n265_adj_4608), 
            .I3(n39510), .O(n19612[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6575_4 (.CI(n39510), .I0(n19739[1]), .I1(n265_adj_4608), 
            .CO(n39511));
    SB_LUT4 add_6499_3_lut (.I0(GND_net), .I1(n19011[0]), .I2(n180_adj_4607), 
            .I3(n39904), .O(n18724[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6575_3_lut (.I0(GND_net), .I1(n19739[0]), .I2(n192), .I3(n39509), 
            .O(n19612[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6575_3 (.CI(n39509), .I0(n19739[0]), .I1(n192), .CO(n39510));
    SB_LUT4 add_6575_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n19612[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6575_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6575_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n39509));
    SB_LUT4 add_6406_16_lut (.I0(GND_net), .I1(n17772[13]), .I2(n1120), 
            .I3(n39508), .O(n17292[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6499_3 (.CI(n39904), .I0(n19011[0]), .I1(n180_adj_4607), 
            .CO(n39905));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n39202), .O(duty_23__N_3772[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6406_15_lut (.I0(GND_net), .I1(n17772[12]), .I2(n1047), 
            .I3(n39507), .O(n17292[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6499_2_lut (.I0(GND_net), .I1(n38_adj_4605), .I2(n107_adj_4604), 
            .I3(GND_net), .O(n18724[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6499_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_15 (.CI(n39507), .I0(n17772[12]), .I1(n1047), .CO(n39508));
    SB_LUT4 add_6406_14_lut (.I0(GND_net), .I1(n17772[11]), .I2(n974), 
            .I3(n39506), .O(n17292[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_14 (.CI(n39506), .I0(n17772[11]), .I1(n974), .CO(n39507));
    SB_LUT4 add_6406_13_lut (.I0(GND_net), .I1(n17772[10]), .I2(n901), 
            .I3(n39505), .O(n17292[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_13 (.CI(n39505), .I0(n17772[10]), .I1(n901), .CO(n39506));
    SB_LUT4 add_6406_12_lut (.I0(GND_net), .I1(n17772[9]), .I2(n828), 
            .I3(n39504), .O(n17292[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_12 (.CI(n39504), .I0(n17772[9]), .I1(n828), .CO(n39505));
    SB_CARRY add_6499_2 (.CI(GND_net), .I0(n38_adj_4605), .I1(n107_adj_4604), 
            .CO(n39904));
    SB_CARRY add_12_22 (.CI(n39202), .I0(n106[20]), .I1(n155[20]), .CO(n39203));
    SB_LUT4 add_6406_11_lut (.I0(GND_net), .I1(n17772[8]), .I2(n755), 
            .I3(n39503), .O(n17292[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n39201), .O(duty_23__N_3772[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_11 (.CI(n39503), .I0(n17772[8]), .I1(n755), .CO(n39504));
    SB_LUT4 add_6406_10_lut (.I0(GND_net), .I1(n17772[7]), .I2(n682), 
            .I3(n39502), .O(n17292[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_10 (.CI(n39502), .I0(n17772[7]), .I1(n682), .CO(n39503));
    SB_LUT4 add_6406_9_lut (.I0(GND_net), .I1(n17772[6]), .I2(n609), .I3(n39501), 
            .O(n17292[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_21 (.CI(n39201), .I0(n106[19]), .I1(n155[19]), .CO(n39202));
    SB_CARRY add_6406_9 (.CI(n39501), .I0(n17772[6]), .I1(n609), .CO(n39502));
    SB_LUT4 add_6406_8_lut (.I0(GND_net), .I1(n17772[5]), .I2(n536), .I3(n39500), 
            .O(n17292[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_8 (.CI(n39500), .I0(n17772[5]), .I1(n536), .CO(n39501));
    SB_LUT4 add_6406_7_lut (.I0(GND_net), .I1(n17772[4]), .I2(n463), .I3(n39499), 
            .O(n17292[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_7 (.CI(n39499), .I0(n17772[4]), .I1(n463), .CO(n39500));
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886_adj_4883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4881));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6406_6_lut (.I0(GND_net), .I1(n17772[3]), .I2(n390), .I3(n39498), 
            .O(n17292[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_6 (.CI(n39498), .I0(n17772[3]), .I1(n390), .CO(n39499));
    SB_LUT4 add_6406_5_lut (.I0(GND_net), .I1(n17772[2]), .I2(n317), .I3(n39497), 
            .O(n17292[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n39200), .O(duty_23__N_3772[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_20 (.CI(n39200), .I0(n106[18]), .I1(n155[18]), .CO(n39201));
    SB_CARRY add_6406_5 (.CI(n39497), .I0(n17772[2]), .I1(n317), .CO(n39498));
    SB_LUT4 add_6406_4_lut (.I0(GND_net), .I1(n17772[1]), .I2(n244), .I3(n39496), 
            .O(n17292[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_4 (.CI(n39496), .I0(n17772[1]), .I1(n244), .CO(n39497));
    SB_LUT4 add_6406_3_lut (.I0(GND_net), .I1(n17772[0]), .I2(n171), .I3(n39495), 
            .O(n17292[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_3 (.CI(n39495), .I0(n17772[0]), .I1(n171), .CO(n39496));
    SB_LUT4 add_6406_2_lut (.I0(GND_net), .I1(n29_adj_4573), .I2(n98), 
            .I3(GND_net), .O(n17292[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6406_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n39199), .O(duty_23__N_3772[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6406_2 (.CI(GND_net), .I0(n29_adj_4573), .I1(n98), .CO(n39495));
    SB_CARRY add_12_19 (.CI(n39199), .I0(n106[17]), .I1(n155[17]), .CO(n39200));
    SB_LUT4 add_6435_15_lut (.I0(GND_net), .I1(n18192[12]), .I2(n1050), 
            .I3(n39494), .O(n17772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6435_14_lut (.I0(GND_net), .I1(n18192[11]), .I2(n977), 
            .I3(n39493), .O(n17772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_14 (.CI(n39493), .I0(n18192[11]), .I1(n977), .CO(n39494));
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n39198), .O(duty_23__N_3772[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6435_13_lut (.I0(GND_net), .I1(n18192[10]), .I2(n904), 
            .I3(n39492), .O(n17772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_13 (.CI(n39492), .I0(n18192[10]), .I1(n904), .CO(n39493));
    SB_LUT4 add_6435_12_lut (.I0(GND_net), .I1(n18192[9]), .I2(n831), 
            .I3(n39491), .O(n17772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_18 (.CI(n39198), .I0(n106[16]), .I1(n155[16]), .CO(n39199));
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n39197), .O(duty_23__N_3772[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_12 (.CI(n39491), .I0(n18192[9]), .I1(n831), .CO(n39492));
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4873));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4870));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6435_11_lut (.I0(GND_net), .I1(n18192[8]), .I2(n758), 
            .I3(n39490), .O(n17772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_17 (.CI(n39197), .I0(n106[15]), .I1(n155[15]), .CO(n39198));
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n39196), .O(duty_23__N_3772[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_11 (.CI(n39490), .I0(n18192[8]), .I1(n758), .CO(n39491));
    SB_CARRY add_12_16 (.CI(n39196), .I0(n106[14]), .I1(n155[14]), .CO(n39197));
    SB_LUT4 add_6435_10_lut (.I0(GND_net), .I1(n18192[7]), .I2(n685), 
            .I3(n39489), .O(n17772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n39195), .O(duty_23__N_3772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_10 (.CI(n39489), .I0(n18192[7]), .I1(n685), .CO(n39490));
    SB_CARRY add_12_15 (.CI(n39195), .I0(n106[13]), .I1(n155[13]), .CO(n39196));
    SB_LUT4 add_6435_9_lut (.I0(GND_net), .I1(n18192[6]), .I2(n612), .I3(n39488), 
            .O(n17772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_9 (.CI(n39488), .I0(n18192[6]), .I1(n612), .CO(n39489));
    SB_LUT4 add_6435_8_lut (.I0(GND_net), .I1(n18192[5]), .I2(n539), .I3(n39487), 
            .O(n17772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_8 (.CI(n39487), .I0(n18192[5]), .I1(n539), .CO(n39488));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n39194), .O(duty_23__N_3772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6435_7_lut (.I0(GND_net), .I1(n18192[4]), .I2(n466), .I3(n39486), 
            .O(n17772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n39194), .I0(n106[12]), .I1(n155[12]), .CO(n39195));
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n39193), .O(duty_23__N_3772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_7 (.CI(n39486), .I0(n18192[4]), .I1(n466), .CO(n39487));
    SB_LUT4 add_6435_6_lut (.I0(GND_net), .I1(n18192[3]), .I2(n393), .I3(n39485), 
            .O(n17772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_6 (.CI(n39485), .I0(n18192[3]), .I1(n393), .CO(n39486));
    SB_LUT4 add_6435_5_lut (.I0(GND_net), .I1(n18192[2]), .I2(n320), .I3(n39484), 
            .O(n17772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_5 (.CI(n39484), .I0(n18192[2]), .I1(n320), .CO(n39485));
    SB_LUT4 add_6435_4_lut (.I0(GND_net), .I1(n18192[1]), .I2(n247), .I3(n39483), 
            .O(n17772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6435_4 (.CI(n39483), .I0(n18192[1]), .I1(n247), .CO(n39484));
    SB_LUT4 add_6435_3_lut (.I0(GND_net), .I1(n18192[0]), .I2(n174), .I3(n39482), 
            .O(n17772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_13 (.CI(n39193), .I0(n106[11]), .I1(n155[11]), .CO(n39194));
    SB_CARRY add_6435_3 (.CI(n39482), .I0(n18192[0]), .I1(n174), .CO(n39483));
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n39192), .O(duty_23__N_3772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6435_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n17772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6435_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n39192), .I0(n106[10]), .I1(n155[10]), .CO(n39193));
    SB_CARRY add_6435_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n39482));
    SB_LUT4 add_6325_19_lut (.I0(GND_net), .I1(n16459[16]), .I2(GND_net), 
            .I3(n40032), .O(n15812[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n39191), 
            .O(duty_23__N_3772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6589_8_lut (.I0(GND_net), .I1(n19836[5]), .I2(n560), .I3(n39481), 
            .O(n19739[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6589_7_lut (.I0(GND_net), .I1(n19836[4]), .I2(n487), .I3(n39480), 
            .O(n19739[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n39191), .I0(n106[9]), .I1(n155[9]), .CO(n39192));
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_6589_7 (.CI(n39480), .I0(n19836[4]), .I1(n487), .CO(n39481));
    SB_LUT4 add_6589_6_lut (.I0(GND_net), .I1(n19836[3]), .I2(n414), .I3(n39479), 
            .O(n19739[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6589_6 (.CI(n39479), .I0(n19836[3]), .I1(n414), .CO(n39480));
    SB_LUT4 add_6589_5_lut (.I0(GND_net), .I1(n19836[2]), .I2(n341), .I3(n39478), 
            .O(n19739[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6589_5 (.CI(n39478), .I0(n19836[2]), .I1(n341), .CO(n39479));
    SB_LUT4 add_6589_4_lut (.I0(GND_net), .I1(n19836[1]), .I2(n268), .I3(n39477), 
            .O(n19739[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6589_4 (.CI(n39477), .I0(n19836[1]), .I1(n268), .CO(n39478));
    SB_LUT4 add_6589_3_lut (.I0(GND_net), .I1(n19836[0]), .I2(n195), .I3(n39476), 
            .O(n19739[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6589_3 (.CI(n39476), .I0(n19836[0]), .I1(n195), .CO(n39477));
    SB_LUT4 add_6589_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n19739[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6589_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6589_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n39476));
    SB_LUT4 add_6462_14_lut (.I0(GND_net), .I1(n18556[11]), .I2(n980), 
            .I3(n39475), .O(n18192[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6462_13_lut (.I0(GND_net), .I1(n18556[10]), .I2(n907), 
            .I3(n39474), .O(n18192[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_13 (.CI(n39474), .I0(n18556[10]), .I1(n907), .CO(n39475));
    SB_LUT4 add_6462_12_lut (.I0(GND_net), .I1(n18556[9]), .I2(n834), 
            .I3(n39473), .O(n18192[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_12 (.CI(n39473), .I0(n18556[9]), .I1(n834), .CO(n39474));
    SB_LUT4 add_6462_11_lut (.I0(GND_net), .I1(n18556[8]), .I2(n761), 
            .I3(n39472), .O(n18192[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_11 (.CI(n39472), .I0(n18556[8]), .I1(n761), .CO(n39473));
    SB_LUT4 add_6462_10_lut (.I0(GND_net), .I1(n18556[7]), .I2(n688), 
            .I3(n39471), .O(n18192[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_10 (.CI(n39471), .I0(n18556[7]), .I1(n688), .CO(n39472));
    SB_LUT4 add_6462_9_lut (.I0(GND_net), .I1(n18556[6]), .I2(n615), .I3(n39470), 
            .O(n18192[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_9 (.CI(n39470), .I0(n18556[6]), .I1(n615), .CO(n39471));
    SB_LUT4 add_6462_8_lut (.I0(GND_net), .I1(n18556[5]), .I2(n542), .I3(n39469), 
            .O(n18192[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_8 (.CI(n39469), .I0(n18556[5]), .I1(n542), .CO(n39470));
    SB_LUT4 add_6462_7_lut (.I0(GND_net), .I1(n18556[4]), .I2(n469), .I3(n39468), 
            .O(n18192[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_7 (.CI(n39468), .I0(n18556[4]), .I1(n469), .CO(n39469));
    SB_LUT4 add_6462_6_lut (.I0(GND_net), .I1(n18556[3]), .I2(n396), .I3(n39467), 
            .O(n18192[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_6 (.CI(n39467), .I0(n18556[3]), .I1(n396), .CO(n39468));
    SB_LUT4 add_6462_5_lut (.I0(GND_net), .I1(n18556[2]), .I2(n323), .I3(n39466), 
            .O(n18192[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_5 (.CI(n39466), .I0(n18556[2]), .I1(n323), .CO(n39467));
    SB_LUT4 add_6462_4_lut (.I0(GND_net), .I1(n18556[1]), .I2(n250), .I3(n39465), 
            .O(n18192[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_4 (.CI(n39465), .I0(n18556[1]), .I1(n250), .CO(n39466));
    SB_LUT4 add_6462_3_lut (.I0(GND_net), .I1(n18556[0]), .I2(n177), .I3(n39464), 
            .O(n18192[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_3 (.CI(n39464), .I0(n18556[0]), .I1(n177), .CO(n39465));
    SB_LUT4 add_6462_2_lut (.I0(GND_net), .I1(n35_adj_4535), .I2(n104), 
            .I3(GND_net), .O(n18192[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6462_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6462_2 (.CI(GND_net), .I0(n35_adj_4535), .I1(n104), .CO(n39464));
    SB_LUT4 add_6487_13_lut (.I0(GND_net), .I1(n18868[10]), .I2(n910), 
            .I3(n39463), .O(n18556[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6487_12_lut (.I0(GND_net), .I1(n18868[9]), .I2(n837), 
            .I3(n39462), .O(n18556[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_12 (.CI(n39462), .I0(n18868[9]), .I1(n837), .CO(n39463));
    SB_LUT4 add_6487_11_lut (.I0(GND_net), .I1(n18868[8]), .I2(n764), 
            .I3(n39461), .O(n18556[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_11 (.CI(n39461), .I0(n18868[8]), .I1(n764), .CO(n39462));
    SB_LUT4 add_6487_10_lut (.I0(GND_net), .I1(n18868[7]), .I2(n691), 
            .I3(n39460), .O(n18556[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_10 (.CI(n39460), .I0(n18868[7]), .I1(n691), .CO(n39461));
    SB_LUT4 add_6487_9_lut (.I0(GND_net), .I1(n18868[6]), .I2(n618), .I3(n39459), 
            .O(n18556[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_9 (.CI(n39459), .I0(n18868[6]), .I1(n618), .CO(n39460));
    SB_LUT4 add_6487_8_lut (.I0(GND_net), .I1(n18868[5]), .I2(n545), .I3(n39458), 
            .O(n18556[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_8 (.CI(n39458), .I0(n18868[5]), .I1(n545), .CO(n39459));
    SB_LUT4 add_6487_7_lut (.I0(GND_net), .I1(n18868[4]), .I2(n472), .I3(n39457), 
            .O(n18556[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_7 (.CI(n39457), .I0(n18868[4]), .I1(n472), .CO(n39458));
    SB_LUT4 add_6487_6_lut (.I0(GND_net), .I1(n18868[3]), .I2(n399), .I3(n39456), 
            .O(n18556[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_6 (.CI(n39456), .I0(n18868[3]), .I1(n399), .CO(n39457));
    SB_LUT4 add_6325_18_lut (.I0(GND_net), .I1(n16459[15]), .I2(GND_net), 
            .I3(n40031), .O(n15812[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6487_5_lut (.I0(GND_net), .I1(n18868[2]), .I2(n326), .I3(n39455), 
            .O(n18556[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_5 (.CI(n39455), .I0(n18868[2]), .I1(n326), .CO(n39456));
    SB_LUT4 add_6487_4_lut (.I0(GND_net), .I1(n18868[1]), .I2(n253), .I3(n39454), 
            .O(n18556[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_4 (.CI(n39454), .I0(n18868[1]), .I1(n253), .CO(n39455));
    SB_LUT4 add_6487_3_lut (.I0(GND_net), .I1(n18868[0]), .I2(n180), .I3(n39453), 
            .O(n18556[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6487_3 (.CI(n39453), .I0(n18868[0]), .I1(n180), .CO(n39454));
    SB_CARRY add_6325_18 (.CI(n40031), .I0(n16459[15]), .I1(GND_net), 
            .CO(n40032));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n39190), 
            .O(duty_23__N_3772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n39190), .I0(n106[8]), .I1(n155[8]), .CO(n39191));
    SB_LUT4 add_6487_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n18556[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6487_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_17_lut (.I0(GND_net), .I1(n16459[14]), .I2(GND_net), 
            .I3(n40030), .O(n15812[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_17 (.CI(n40030), .I0(n16459[14]), .I1(GND_net), 
            .CO(n40031));
    SB_CARRY add_6487_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n39453));
    SB_LUT4 add_6601_7_lut (.I0(GND_net), .I1(n45940), .I2(n490_adj_4889), 
            .I3(n39452), .O(n19836[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6601_6_lut (.I0(GND_net), .I1(n19907[3]), .I2(n417_adj_4890), 
            .I3(n39451), .O(n19836[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_16_lut (.I0(GND_net), .I1(n16459[13]), .I2(n1111_adj_4891), 
            .I3(n40029), .O(n15812[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_6 (.CI(n39451), .I0(n19907[3]), .I1(n417_adj_4890), 
            .CO(n39452));
    SB_LUT4 add_6601_5_lut (.I0(GND_net), .I1(n19907[2]), .I2(n344_adj_4892), 
            .I3(n39450), .O(n19836[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_5 (.CI(n39450), .I0(n19907[2]), .I1(n344_adj_4892), 
            .CO(n39451));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n39189), 
            .O(duty_23__N_3772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6601_4_lut (.I0(GND_net), .I1(n19907[1]), .I2(n271_adj_4893), 
            .I3(n39449), .O(n19836[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_4 (.CI(n39449), .I0(n19907[1]), .I1(n271_adj_4893), 
            .CO(n39450));
    SB_CARRY add_6325_16 (.CI(n40029), .I0(n16459[13]), .I1(n1111_adj_4891), 
            .CO(n40030));
    SB_LUT4 add_6601_3_lut (.I0(GND_net), .I1(n19907[0]), .I2(n198_adj_4894), 
            .I3(n39448), .O(n19836[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_3 (.CI(n39448), .I0(n19907[0]), .I1(n198_adj_4894), 
            .CO(n39449));
    SB_LUT4 add_6601_2_lut (.I0(GND_net), .I1(n56_adj_4895), .I2(n125_adj_4896), 
            .I3(GND_net), .O(n19836[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6601_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6601_2 (.CI(GND_net), .I0(n56_adj_4895), .I1(n125_adj_4896), 
            .CO(n39448));
    SB_LUT4 add_6510_12_lut (.I0(GND_net), .I1(n19132[9]), .I2(n840_adj_4897), 
            .I3(n39440), .O(n18868[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6510_11_lut (.I0(GND_net), .I1(n19132[8]), .I2(n767_adj_4898), 
            .I3(n39439), .O(n18868[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_11 (.CI(n39439), .I0(n19132[8]), .I1(n767_adj_4898), 
            .CO(n39440));
    SB_LUT4 add_6510_10_lut (.I0(GND_net), .I1(n19132[7]), .I2(n694_adj_4899), 
            .I3(n39438), .O(n18868[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_10 (.CI(n39438), .I0(n19132[7]), .I1(n694_adj_4899), 
            .CO(n39439));
    SB_LUT4 add_6510_9_lut (.I0(GND_net), .I1(n19132[6]), .I2(n621_adj_4900), 
            .I3(n39437), .O(n18868[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_9 (.CI(n39437), .I0(n19132[6]), .I1(n621_adj_4900), 
            .CO(n39438));
    SB_LUT4 add_6510_8_lut (.I0(GND_net), .I1(n19132[5]), .I2(n548_adj_4901), 
            .I3(n39436), .O(n18868[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_8 (.CI(n39436), .I0(n19132[5]), .I1(n548_adj_4901), 
            .CO(n39437));
    SB_LUT4 add_6510_7_lut (.I0(GND_net), .I1(n19132[4]), .I2(n475_adj_4902), 
            .I3(n39435), .O(n18868[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_7 (.CI(n39435), .I0(n19132[4]), .I1(n475_adj_4902), 
            .CO(n39436));
    SB_LUT4 add_6510_6_lut (.I0(GND_net), .I1(n19132[3]), .I2(n402_adj_4903), 
            .I3(n39434), .O(n18868[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_6 (.CI(n39434), .I0(n19132[3]), .I1(n402_adj_4903), 
            .CO(n39435));
    SB_LUT4 add_6510_5_lut (.I0(GND_net), .I1(n19132[2]), .I2(n329_adj_4904), 
            .I3(n39433), .O(n18868[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_5 (.CI(n39433), .I0(n19132[2]), .I1(n329_adj_4904), 
            .CO(n39434));
    SB_LUT4 add_6510_4_lut (.I0(GND_net), .I1(n19132[1]), .I2(n256_adj_4905), 
            .I3(n39432), .O(n18868[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_4 (.CI(n39432), .I0(n19132[1]), .I1(n256_adj_4905), 
            .CO(n39433));
    SB_LUT4 add_6510_3_lut (.I0(GND_net), .I1(n19132[0]), .I2(n183_adj_4906), 
            .I3(n39431), .O(n18868[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_3 (.CI(n39431), .I0(n19132[0]), .I1(n183_adj_4906), 
            .CO(n39432));
    SB_LUT4 add_6510_2_lut (.I0(GND_net), .I1(n41_adj_4907), .I2(n110_adj_4908), 
            .I3(GND_net), .O(n18868[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6510_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6510_2 (.CI(GND_net), .I0(n41_adj_4907), .I1(n110_adj_4908), 
            .CO(n39431));
    SB_CARRY add_12_9 (.CI(n39189), .I0(n106[7]), .I1(n155[7]), .CO(n39190));
    SB_LUT4 add_6531_11_lut (.I0(GND_net), .I1(n19352[8]), .I2(n770_adj_4909), 
            .I3(n39417), .O(n19132[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_10_lut (.I0(GND_net), .I1(n19352[7]), .I2(n697_adj_4910), 
            .I3(n39416), .O(n19132[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_10 (.CI(n39416), .I0(n19352[7]), .I1(n697_adj_4910), 
            .CO(n39417));
    SB_LUT4 add_6531_9_lut (.I0(GND_net), .I1(n19352[6]), .I2(n624_adj_4911), 
            .I3(n39415), .O(n19132[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_9 (.CI(n39415), .I0(n19352[6]), .I1(n624_adj_4911), 
            .CO(n39416));
    SB_LUT4 add_6531_8_lut (.I0(GND_net), .I1(n19352[5]), .I2(n551_adj_4912), 
            .I3(n39414), .O(n19132[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_8 (.CI(n39414), .I0(n19352[5]), .I1(n551_adj_4912), 
            .CO(n39415));
    SB_LUT4 add_6531_7_lut (.I0(GND_net), .I1(n19352[4]), .I2(n478_adj_4913), 
            .I3(n39413), .O(n19132[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_7 (.CI(n39413), .I0(n19352[4]), .I1(n478_adj_4913), 
            .CO(n39414));
    SB_LUT4 add_6531_6_lut (.I0(GND_net), .I1(n19352[3]), .I2(n405_adj_4914), 
            .I3(n39412), .O(n19132[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_15_lut (.I0(GND_net), .I1(n16459[12]), .I2(n1038_adj_4915), 
            .I3(n40028), .O(n15812[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_6 (.CI(n39412), .I0(n19352[3]), .I1(n405_adj_4914), 
            .CO(n39413));
    SB_LUT4 add_6531_5_lut (.I0(GND_net), .I1(n19352[2]), .I2(n332_adj_4916), 
            .I3(n39411), .O(n19132[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_15 (.CI(n40028), .I0(n16459[12]), .I1(n1038_adj_4915), 
            .CO(n40029));
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n39188), 
            .O(duty_23__N_3772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_5 (.CI(n39411), .I0(n19352[2]), .I1(n332_adj_4916), 
            .CO(n39412));
    SB_LUT4 add_6531_4_lut (.I0(GND_net), .I1(n19352[1]), .I2(n259_adj_4917), 
            .I3(n39410), .O(n19132[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_4 (.CI(n39410), .I0(n19352[1]), .I1(n259_adj_4917), 
            .CO(n39411));
    SB_LUT4 add_6531_3_lut (.I0(GND_net), .I1(n19352[0]), .I2(n186_adj_4918), 
            .I3(n39409), .O(n19132[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_3 (.CI(n39409), .I0(n19352[0]), .I1(n186_adj_4918), 
            .CO(n39410));
    SB_LUT4 add_6325_14_lut (.I0(GND_net), .I1(n16459[11]), .I2(n965_adj_4919), 
            .I3(n40027), .O(n15812[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6531_2_lut (.I0(GND_net), .I1(n44_adj_4920), .I2(n113_adj_4921), 
            .I3(GND_net), .O(n19132[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6531_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6531_2 (.CI(GND_net), .I0(n44_adj_4920), .I1(n113_adj_4921), 
            .CO(n39409));
    SB_CARRY add_6325_14 (.CI(n40027), .I0(n16459[11]), .I1(n965_adj_4919), 
            .CO(n40028));
    SB_LUT4 add_6521_12_lut (.I0(GND_net), .I1(n19252[9]), .I2(n840), 
            .I3(n39882), .O(n19011[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_10_lut (.I0(GND_net), .I1(n19532[7]), .I2(n700_adj_4875), 
            .I3(n39408), .O(n19352[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_9_lut (.I0(GND_net), .I1(n19532[6]), .I2(n627_adj_4872), 
            .I3(n39407), .O(n19352[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_9 (.CI(n39407), .I0(n19532[6]), .I1(n627_adj_4872), 
            .CO(n39408));
    SB_CARRY add_12_8 (.CI(n39188), .I0(n106[6]), .I1(n155[6]), .CO(n39189));
    SB_LUT4 add_6521_11_lut (.I0(GND_net), .I1(n19252[8]), .I2(n767), 
            .I3(n39881), .O(n19011[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_8_lut (.I0(GND_net), .I1(n19532[5]), .I2(n554_adj_4866), 
            .I3(n39406), .O(n19352[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_8 (.CI(n39406), .I0(n19532[5]), .I1(n554_adj_4866), 
            .CO(n39407));
    SB_LUT4 add_6325_13_lut (.I0(GND_net), .I1(n16459[10]), .I2(n892_adj_4857), 
            .I3(n40026), .O(n15812[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_13 (.CI(n40026), .I0(n16459[10]), .I1(n892_adj_4857), 
            .CO(n40027));
    SB_CARRY add_6521_11 (.CI(n39881), .I0(n19252[8]), .I1(n767), .CO(n39882));
    SB_LUT4 add_6521_10_lut (.I0(GND_net), .I1(n19252[7]), .I2(n694), 
            .I3(n39880), .O(n19011[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n39187), 
            .O(duty_23__N_3772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_7_lut (.I0(GND_net), .I1(n19532[4]), .I2(n481_adj_4848), 
            .I3(n39405), .O(n19352[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_7 (.CI(n39405), .I0(n19532[4]), .I1(n481_adj_4848), 
            .CO(n39406));
    SB_LUT4 add_6550_6_lut (.I0(GND_net), .I1(n19532[3]), .I2(n408_adj_4844), 
            .I3(n39404), .O(n19352[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_12_lut (.I0(GND_net), .I1(n16459[9]), .I2(n819_adj_4843), 
            .I3(n40025), .O(n15812[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_12 (.CI(n40025), .I0(n16459[9]), .I1(n819_adj_4843), 
            .CO(n40026));
    SB_CARRY add_6550_6 (.CI(n39404), .I0(n19532[3]), .I1(n408_adj_4844), 
            .CO(n39405));
    SB_LUT4 add_6550_5_lut (.I0(GND_net), .I1(n19532[2]), .I2(n335_adj_4842), 
            .I3(n39403), .O(n19352[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_10 (.CI(n39880), .I0(n19252[7]), .I1(n694), .CO(n39881));
    SB_LUT4 add_6521_9_lut (.I0(GND_net), .I1(n19252[6]), .I2(n621), .I3(n39879), 
            .O(n19011[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n39187), .I0(n106[5]), .I1(n155[5]), .CO(n39188));
    SB_CARRY add_6550_5 (.CI(n39403), .I0(n19532[2]), .I1(n335_adj_4842), 
            .CO(n39404));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n39186), 
            .O(duty_23__N_3772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_4_lut (.I0(GND_net), .I1(n19532[1]), .I2(n262_adj_4839), 
            .I3(n39402), .O(n19352[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_4 (.CI(n39402), .I0(n19532[1]), .I1(n262_adj_4839), 
            .CO(n39403));
    SB_LUT4 add_6325_11_lut (.I0(GND_net), .I1(n16459[8]), .I2(n746_adj_4838), 
            .I3(n40024), .O(n15812[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_9 (.CI(n39879), .I0(n19252[6]), .I1(n621), .CO(n39880));
    SB_CARRY add_12_6 (.CI(n39186), .I0(n106[4]), .I1(n155[4]), .CO(n39187));
    SB_LUT4 add_6550_3_lut (.I0(GND_net), .I1(n19532[0]), .I2(n189_adj_4830), 
            .I3(n39401), .O(n19352[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_11 (.CI(n40024), .I0(n16459[8]), .I1(n746_adj_4838), 
            .CO(n40025));
    SB_LUT4 add_6521_8_lut (.I0(GND_net), .I1(n19252[5]), .I2(n548), .I3(n39878), 
            .O(n19011[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6550_3 (.CI(n39401), .I0(n19532[0]), .I1(n189_adj_4830), 
            .CO(n39402));
    SB_LUT4 add_6325_10_lut (.I0(GND_net), .I1(n16459[7]), .I2(n673_adj_4821), 
            .I3(n40023), .O(n15812[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6521_8 (.CI(n39878), .I0(n19252[5]), .I1(n548), .CO(n39879));
    SB_LUT4 add_6521_7_lut (.I0(GND_net), .I1(n19252[4]), .I2(n475), .I3(n39877), 
            .O(n19011[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6521_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n39185), 
            .O(duty_23__N_3772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6550_2_lut (.I0(GND_net), .I1(n47_adj_4812), .I2(n116_adj_4811), 
            .I3(GND_net), .O(n19352[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6550_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_10 (.CI(n40023), .I0(n16459[7]), .I1(n673_adj_4821), 
            .CO(n40024));
    SB_CARRY add_6550_2 (.CI(GND_net), .I0(n47_adj_4812), .I1(n116_adj_4811), 
            .CO(n39401));
    SB_LUT4 add_6567_9_lut (.I0(GND_net), .I1(n19676[6]), .I2(n630_adj_4810), 
            .I3(n39400), .O(n19532[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6567_8_lut (.I0(GND_net), .I1(n19676[5]), .I2(n557_adj_4809), 
            .I3(n39399), .O(n19532[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_8 (.CI(n39399), .I0(n19676[5]), .I1(n557_adj_4809), 
            .CO(n39400));
    SB_LUT4 add_6567_7_lut (.I0(GND_net), .I1(n19676[4]), .I2(n484_adj_4808), 
            .I3(n39398), .O(n19532[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_9_lut (.I0(GND_net), .I1(n16459[6]), .I2(n600_adj_4805), 
            .I3(n40022), .O(n15812[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_7 (.CI(n39398), .I0(n19676[4]), .I1(n484_adj_4808), 
            .CO(n39399));
    SB_CARRY add_12_5 (.CI(n39185), .I0(n106[3]), .I1(n155[3]), .CO(n39186));
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n39184), 
            .O(duty_23__N_3772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_9 (.CI(n40022), .I0(n16459[6]), .I1(n600_adj_4805), 
            .CO(n40023));
    SB_LUT4 add_6567_6_lut (.I0(GND_net), .I1(n19676[3]), .I2(n411_adj_4803), 
            .I3(n39397), .O(n19532[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_6 (.CI(n39397), .I0(n19676[3]), .I1(n411_adj_4803), 
            .CO(n39398));
    SB_CARRY add_12_4 (.CI(n39184), .I0(n106[2]), .I1(n155[2]), .CO(n39185));
    SB_LUT4 add_6567_5_lut (.I0(GND_net), .I1(n19676[2]), .I2(n338_adj_4796), 
            .I3(n39396), .O(n19532[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_5 (.CI(n39396), .I0(n19676[2]), .I1(n338_adj_4796), 
            .CO(n39397));
    SB_LUT4 add_6567_4_lut (.I0(GND_net), .I1(n19676[1]), .I2(n265_adj_4795), 
            .I3(n39395), .O(n19532[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_4 (.CI(n39395), .I0(n19676[1]), .I1(n265_adj_4795), 
            .CO(n39396));
    SB_LUT4 add_6567_3_lut (.I0(GND_net), .I1(n19676[0]), .I2(n192_adj_4792), 
            .I3(n39394), .O(n19532[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6325_8_lut (.I0(GND_net), .I1(n16459[5]), .I2(n527_adj_4790), 
            .I3(n40021), .O(n15812[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_3 (.CI(n39394), .I0(n19676[0]), .I1(n192_adj_4792), 
            .CO(n39395));
    SB_CARRY add_6325_8 (.CI(n40021), .I0(n16459[5]), .I1(n527_adj_4790), 
            .CO(n40022));
    SB_LUT4 add_6567_2_lut (.I0(GND_net), .I1(n50_adj_4789), .I2(n119_adj_4788), 
            .I3(GND_net), .O(n19532[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6567_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6567_2 (.CI(GND_net), .I0(n50_adj_4789), .I1(n119_adj_4788), 
            .CO(n39394));
    SB_LUT4 add_6325_7_lut (.I0(GND_net), .I1(n16459[4]), .I2(n454_adj_4786), 
            .I3(n40020), .O(n15812[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6582_8_lut (.I0(GND_net), .I1(n19788[5]), .I2(n560_adj_4785), 
            .I3(n39393), .O(n19676[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6582_7_lut (.I0(GND_net), .I1(n19788[4]), .I2(n487_adj_4784), 
            .I3(n39392), .O(n19676[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_7 (.CI(n39392), .I0(n19788[4]), .I1(n487_adj_4784), 
            .CO(n39393));
    SB_LUT4 add_6582_6_lut (.I0(GND_net), .I1(n19788[3]), .I2(n414_adj_4783), 
            .I3(n39391), .O(n19676[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_6 (.CI(n39391), .I0(n19788[3]), .I1(n414_adj_4783), 
            .CO(n39392));
    SB_LUT4 add_6582_5_lut (.I0(GND_net), .I1(n19788[2]), .I2(n341_adj_4781), 
            .I3(n39390), .O(n19676[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_7 (.CI(n40020), .I0(n16459[4]), .I1(n454_adj_4786), 
            .CO(n40021));
    SB_CARRY add_6582_5 (.CI(n39390), .I0(n19788[2]), .I1(n341_adj_4781), 
            .CO(n39391));
    SB_LUT4 add_6325_6_lut (.I0(GND_net), .I1(n16459[3]), .I2(n381_adj_4777), 
            .I3(n40019), .O(n15812[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n39183), 
            .O(duty_23__N_3772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6582_4_lut (.I0(GND_net), .I1(n19788[1]), .I2(n268_adj_4774), 
            .I3(n39389), .O(n19676[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_4 (.CI(n39389), .I0(n19788[1]), .I1(n268_adj_4774), 
            .CO(n39390));
    SB_LUT4 add_6582_3_lut (.I0(GND_net), .I1(n19788[0]), .I2(n195_adj_4773), 
            .I3(n39388), .O(n19676[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_3 (.CI(n39388), .I0(n19788[0]), .I1(n195_adj_4773), 
            .CO(n39389));
    SB_LUT4 add_6582_2_lut (.I0(GND_net), .I1(n53_adj_4768), .I2(n122_adj_4767), 
            .I3(GND_net), .O(n19676[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6582_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6582_2 (.CI(GND_net), .I0(n53_adj_4768), .I1(n122_adj_4767), 
            .CO(n39388));
    SB_CARRY add_6325_6 (.CI(n40019), .I0(n16459[3]), .I1(n381_adj_4777), 
            .CO(n40020));
    SB_CARRY add_12_3 (.CI(n39183), .I0(n106[1]), .I1(n155[1]), .CO(n39184));
    SB_LUT4 add_6595_7_lut (.I0(GND_net), .I1(n45611), .I2(n490), .I3(n39387), 
            .O(n19788[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6595_6_lut (.I0(GND_net), .I1(n19872[3]), .I2(n417), .I3(n39386), 
            .O(n19788[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_6 (.CI(n39386), .I0(n19872[3]), .I1(n417), .CO(n39387));
    SB_LUT4 add_6595_5_lut (.I0(GND_net), .I1(n19872[2]), .I2(n344), .I3(n39385), 
            .O(n19788[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_5 (.CI(n39385), .I0(n19872[2]), .I1(n344), .CO(n39386));
    SB_LUT4 add_6325_5_lut (.I0(GND_net), .I1(n16459[2]), .I2(n308_adj_4739), 
            .I3(n40018), .O(n15812[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6595_4_lut (.I0(GND_net), .I1(n19872[1]), .I2(n271_adj_4738), 
            .I3(n39384), .O(n19788[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_4 (.CI(n39384), .I0(n19872[1]), .I1(n271_adj_4738), 
            .CO(n39385));
    SB_LUT4 add_6595_3_lut (.I0(GND_net), .I1(n19872[0]), .I2(n198), .I3(n39383), 
            .O(n19788[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_3 (.CI(n39383), .I0(n19872[0]), .I1(n198), .CO(n39384));
    SB_LUT4 add_6595_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n19788[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6595_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6595_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n39383));
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n39183));
    SB_CARRY add_6325_5 (.CI(n40018), .I0(n16459[2]), .I1(n308_adj_4739), 
            .CO(n40019));
    SB_LUT4 add_6325_4_lut (.I0(GND_net), .I1(n16459[1]), .I2(n235_adj_4730), 
            .I3(n40017), .O(n15812[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_4 (.CI(n40017), .I0(n16459[1]), .I1(n235_adj_4730), 
            .CO(n40018));
    SB_LUT4 add_6325_3_lut (.I0(GND_net), .I1(n16459[0]), .I2(n162_adj_4727), 
            .I3(n40016), .O(n15812[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_3 (.CI(n40016), .I0(n16459[0]), .I1(n162_adj_4727), 
            .CO(n40017));
    SB_LUT4 add_6325_2_lut (.I0(GND_net), .I1(n20_adj_4720), .I2(n89_adj_4719), 
            .I3(GND_net), .O(n15812[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6325_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6325_2 (.CI(GND_net), .I0(n20_adj_4720), .I1(n89_adj_4719), 
            .CO(n40016));
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[23]), 
            .I3(n39348), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[22]), 
            .I3(n39347), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n39347), .I0(GND_net), .I1(n1_adj_4929[22]), 
            .CO(n39348));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[21]), 
            .I3(n39346), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n39346), .I0(GND_net), .I1(n1_adj_4929[21]), 
            .CO(n39347));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[20]), 
            .I3(n39345), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_18_lut (.I0(GND_net), .I1(n17036[15]), .I2(GND_net), 
            .I3(n40015), .O(n16459[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n39345), .I0(GND_net), .I1(n1_adj_4929[20]), 
            .CO(n39346));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[19]), 
            .I3(n39344), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n39344), .I0(GND_net), .I1(n1_adj_4929[19]), 
            .CO(n39345));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[18]), 
            .I3(n39343), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n39343), .I0(GND_net), .I1(n1_adj_4929[18]), 
            .CO(n39344));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[17]), 
            .I3(n39342), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n39342), .I0(GND_net), .I1(n1_adj_4929[17]), 
            .CO(n39343));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[16]), 
            .I3(n39341), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_17_lut (.I0(GND_net), .I1(n17036[14]), .I2(GND_net), 
            .I3(n40014), .O(n16459[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_17 (.CI(n40014), .I0(n17036[14]), .I1(GND_net), 
            .CO(n40015));
    SB_CARRY unary_minus_16_add_3_18 (.CI(n39341), .I0(GND_net), .I1(n1_adj_4929[16]), 
            .CO(n39342));
    SB_LUT4 add_6359_16_lut (.I0(GND_net), .I1(n17036[13]), .I2(n1114_adj_4707), 
            .I3(n40013), .O(n16459[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[15]), 
            .I3(n39340), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_16 (.CI(n40013), .I0(n17036[13]), .I1(n1114_adj_4707), 
            .CO(n40014));
    SB_CARRY unary_minus_16_add_3_17 (.CI(n39340), .I0(GND_net), .I1(n1_adj_4929[15]), 
            .CO(n39341));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[14]), 
            .I3(n39339), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n39339), .I0(GND_net), .I1(n1_adj_4929[14]), 
            .CO(n39340));
    SB_LUT4 add_6359_15_lut (.I0(GND_net), .I1(n17036[12]), .I2(n1041_adj_4703), 
            .I3(n40012), .O(n16459[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[13]), 
            .I3(n39338), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n39338), .I0(GND_net), .I1(n1_adj_4929[13]), 
            .CO(n39339));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[12]), 
            .I3(n39337), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n39337), .I0(GND_net), .I1(n1_adj_4929[12]), 
            .CO(n39338));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[11]), 
            .I3(n39336), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_15 (.CI(n40012), .I0(n17036[12]), .I1(n1041_adj_4703), 
            .CO(n40013));
    SB_LUT4 add_6359_14_lut (.I0(GND_net), .I1(n17036[11]), .I2(n968_adj_4695), 
            .I3(n40011), .O(n16459[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n39336), .I0(GND_net), .I1(n1_adj_4929[11]), 
            .CO(n39337));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[10]), 
            .I3(n39335), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n39335), .I0(GND_net), .I1(n1_adj_4929[10]), 
            .CO(n39336));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[9]), 
            .I3(n39334), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n39334), .I0(GND_net), .I1(n1_adj_4929[9]), 
            .CO(n39335));
    SB_CARRY add_6359_14 (.CI(n40011), .I0(n17036[11]), .I1(n968_adj_4695), 
            .CO(n40012));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[8]), 
            .I3(n39333), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n39333), .I0(GND_net), .I1(n1_adj_4929[8]), 
            .CO(n39334));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[7]), 
            .I3(n39332), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n39332), .I0(GND_net), .I1(n1_adj_4929[7]), 
            .CO(n39333));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[6]), 
            .I3(n39331), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n39331), .I0(GND_net), .I1(n1_adj_4929[6]), 
            .CO(n39332));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[5]), 
            .I3(n39330), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n39330), .I0(GND_net), .I1(n1_adj_4929[5]), 
            .CO(n39331));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[4]), 
            .I3(n39329), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_13_lut (.I0(GND_net), .I1(n17036[10]), .I2(n895_adj_4665), 
            .I3(n40010), .O(n16459[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n39329), .I0(GND_net), .I1(n1_adj_4929[4]), 
            .CO(n39330));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[3]), 
            .I3(n39328), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n39328), .I0(GND_net), .I1(n1_adj_4929[3]), 
            .CO(n39329));
    SB_CARRY add_6359_13 (.CI(n40010), .I0(n17036[10]), .I1(n895_adj_4665), 
            .CO(n40011));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[2]), 
            .I3(n39327), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n39327), .I0(GND_net), .I1(n1_adj_4929[2]), 
            .CO(n39328));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[1]), 
            .I3(n39326), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n39326), .I0(GND_net), .I1(n1_adj_4929[1]), 
            .CO(n39327));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4929[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6359_12_lut (.I0(GND_net), .I1(n17036[9]), .I2(n822_adj_4644), 
            .I3(n40009), .O(n16459[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6359_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4929[0]), 
            .CO(n39326));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4928[23]), 
            .I3(n39325), .O(\PID_CONTROLLER.integral_23__N_3723 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6359_12 (.CI(n40009), .I0(n17036[9]), .I1(n822_adj_4644), 
            .CO(n40010));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4928[22]), .I3(n39324), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n39324), .I0(GND_net), .I1(n1_adj_4928[22]), 
            .CO(n39325));
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4921));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959_adj_4859));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4858));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032_adj_4856));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4855));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4920));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4919));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_4918));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4854));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105_adj_4853));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_4917));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4845));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21891_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21891_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21890_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21890_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_4916));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4915));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_4914));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4841));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4840));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4836));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4835));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4833));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4832));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4829));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4827));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4823));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4818));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4817));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4815));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4814));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4813));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4806));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4802));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4801));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21889_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21889_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4800));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_4913));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_4912));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4799));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4798));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4797));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_4911));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4794));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_4910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_4909));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4793));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4791));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34548_3_lut_4_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3772[2]), .O(n49985));   // verilog/motorControl.v(38[19:35])
    defparam i34548_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4598));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4787));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4908));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4782));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4906));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4780));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4905));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4779));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4778));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4776));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34587_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(PWMLimit[2]), .O(n50024));   // verilog/motorControl.v(36[10:25])
    defparam i34587_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4775));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_4904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_4903));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_4902));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4771));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_4901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4766));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_4900));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_4899));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4765));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_4898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_4897));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4763));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(GND_net), .O(n6_adj_4569));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4762));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4896));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4894));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4893));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4750));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4748));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4745));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4742));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4741));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21888_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21888_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4728));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4726));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4725));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21887_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21887_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4716));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4715));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4713));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4705));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3772[1]), .I1(n257[1]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3747[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3772[2]), .I1(n257[2]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3747[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3747[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3747[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3747[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3747[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3747[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3747[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3747[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3747[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3747[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3747[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3747[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3747[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3747[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3747[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3747[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3747[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3747[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3747[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3747[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3747[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3772[23]), .I1(n257[23]), .I2(n256_adj_4602), 
            .I3(GND_net), .O(duty_23__N_3747[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3747[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4699));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4698));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4891));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4890));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1528 (.I0(n6_adj_4888), .I1(\Kp[4] ), .I2(n19956[2]), 
            .I3(n1[18]), .O(n19907[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1528.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25394_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .O(n19932[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25394_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4684));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4683));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4680));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4677));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21886_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21886_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4675));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4674));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4672));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4671));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4669));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34515_2_lut_4_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(duty_23__N_3772[9]), .I3(n257[9]), .O(n49952));
    defparam i34515_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i34525_2_lut_4_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(duty_23__N_3772[7]), .I3(n257[7]), .O(n49962));
    defparam i34525_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i34550_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3772[9]), .O(n49987));
    defparam i34550_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4668));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4666));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34560_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3772[7]), .O(n49997));
    defparam i34560_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4660));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25379_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n20004[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25379_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_1529 (.I0(n4_adj_4886), .I1(\Kp[3] ), .I2(n19987[1]), 
            .I3(n1[19]), .O(n19956[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1529.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1530 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_4922));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1530.LUT_INIT = 16'h9c50;
    SB_LUT4 i25547_4_lut (.I0(n19956[2]), .I1(\Kp[4] ), .I2(n6_adj_4888), 
            .I3(n1[18]), .O(n8_adj_4923));   // verilog/motorControl.v(34[16:22])
    defparam i25547_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i21885_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21885_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4654));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1531 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), 
            .I3(n1[21]), .O(n11_adj_4924));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut_adj_1531.LUT_INIT = 16'h6ca0;
    SB_LUT4 i25508_4_lut (.I0(n19987[1]), .I1(\Kp[3] ), .I2(n4_adj_4886), 
            .I3(n1[19]), .O(n6_adj_4925));   // verilog/motorControl.v(34[16:22])
    defparam i25508_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4522));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25381_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n38861));   // verilog/motorControl.v(34[16:22])
    defparam i25381_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4652));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4651));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1532 (.I0(n6_adj_4925), .I1(n11_adj_4924), .I2(n8_adj_4923), 
            .I3(n12_adj_4922), .O(n18_adj_4926));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1533 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), 
            .I3(n1[22]), .O(n13_adj_4927));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut_adj_1533.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1534 (.I0(n13_adj_4927), .I1(n18_adj_4926), .I2(n38861), 
            .I3(n4_adj_4869), .O(n45940));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4928[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21884_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4096[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i21884_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module coms
//

module coms (\data_in_frame[1] , \data_in_frame[3] , CLK_c, GND_net, 
            n29756, control_mode, n25135, \data_in_frame[2] , \data_out_frame[14] , 
            \data_out_frame[15] , \data_out_frame[12] , \data_out_frame[13] , 
            n29755, \FRAME_MATCHER.i_31__N_2622 , n29754, \FRAME_MATCHER.state_31__N_2660[2] , 
            \FRAME_MATCHER.i_31__N_2626 , n4452, n7, rx_data, n771, 
            n29753, n29752, n45880, n3303, \data_in[2] , \data_in[0] , 
            \data_in[3] , \data_in[1] , n63, \data_out_frame[8] , \data_out_frame[9] , 
            \data_out_frame[10] , \data_out_frame[11] , n29751, n29750, 
            n29749, PWMLimit, n29748, \data_in_frame[8] , \FRAME_MATCHER.state[0] , 
            n29747, rx_data_ready, setpoint, n29746, \data_in_frame[10] , 
            n29745, \data_in_frame[11] , \data_in_frame[13] , n29744, 
            n29743, n29742, n29741, n29740, n29739, n29738, n29737, 
            n29736, n29735, n29734, n29733, n29732, n29731, n29730, 
            n29729, n29728, n29727, n51593, n51594, \data_in_frame[9] , 
            \data_out_frame[16] , \data_out_frame[17] , \data_out_frame[18] , 
            \data_out_frame[19] , \data_out_frame[23] , \data_out_frame[20] , 
            n14, tx_active, DE_c, LED_c, \data_out_frame[6] , \data_out_frame[7] , 
            \data_out_frame[4] , \data_out_frame[5] , n25063, \data_in_frame[12] , 
            \data_in_frame[4] , \data_in_frame[6] , \data_in_frame[5] , 
            n29310, \data_out_frame[25] , \data_out_frame[24] , \data_out_frame[27][1] , 
            ID, n4, n29176, n41916, n30209, IntegralLimit, n30208, 
            n30207, n30206, n30205, n30204, n30203, n30202, n30201, 
            n30200, n30199, n30198, n30197, n30196, n30195, n30194, 
            n30193, n30192, n30191, n30190, n30189, n30188, n30186, 
            n30185, n30184, n30183, n30182, n30181, n30180, n30179, 
            n30178, n30177, n30176, n30175, n30174, n30173, n30172, 
            n30171, n30170, n30169, n30168, n30167, n30166, n30165, 
            n30164, n30163, n30162, n30161, n30160, n30159, n30158, 
            n30157, n30156, n30155, n30154, \Kp[1] , n30153, \Kp[2] , 
            n30152, \Kp[3] , n30151, \Kp[4] , n30150, \Kp[5] , n30149, 
            \Kp[6] , n30148, \Kp[7] , n30147, \Kp[8] , n30146, \Kp[9] , 
            n30145, \Kp[10] , n30144, \Kp[11] , n30143, \Kp[12] , 
            n30141, \Kp[13] , n30140, \Kp[14] , n30139, \Kp[15] , 
            n30138, \Ki[1] , n30137, \Ki[2] , n30136, \Ki[3] , n30135, 
            \Ki[4] , n30134, \Ki[5] , n30133, \Ki[6] , n30132, \Ki[7] , 
            n30131, \Ki[8] , n30130, \Ki[9] , n30129, \Ki[10] , 
            n30128, \Ki[11] , n30127, \Ki[12] , n30126, \Ki[13] , 
            n30125, \Ki[14] , n30124, \Ki[15] , n30123, n30122, 
            n30121, n30120, n30119, n30118, n30117, n30116, n30115, 
            n30114, n30113, n30112, n30111, n30110, n30109, n30108, 
            n30107, n30106, n30105, n30104, n30103, n30102, n30101, 
            n30100, n30099, n30098, n30097, n30096, n30095, n30094, 
            n30093, n30092, n30091, n30090, n30089, n30088, n30087, 
            n30086, n30085, n30084, n30083, n30082, n30081, n30080, 
            n30079, n30078, n30077, n30076, n30075, n30074, n30073, 
            n30072, n30071, n30070, n30069, n30068, n30067, n30066, 
            n30065, n30064, n30063, n30062, n30061, n30060, n30059, 
            n30058, n30057, n30056, n30055, n30054, n30053, n30052, 
            n30051, n30050, n30049, n30048, n30047, n30046, n30045, 
            n30044, n30043, n30042, n30041, n30040, n30039, n30038, 
            n30037, n30036, n30035, n30034, n30033, n30032, n30031, 
            n30030, n30029, n30028, n30027, n30026, n30025, n30024, 
            n30023, n30022, n30021, n30020, n30019, n30018, n30017, 
            n30016, n30015, n30014, n30013, n30012, n30011, n30009, 
            n30008, n30007, n30006, n30005, n30004, n30003, n30002, 
            n30001, n30000, n29999, n29998, n29997, n29996, n29995, 
            n29994, n29993, n29992, n29991, n29990, n29989, n29988, 
            n29987, n29986, n29985, n29984, n29983, n29982, n29981, 
            n29980, n29979, n29978, n29977, n29976, n29975, n29974, 
            n29973, n29972, n29971, n29970, n29969, n29968, n29967, 
            n29966, n29965, n29964, n29963, n29962, n29961, neopxl_color, 
            n29960, n29959, n29958, n29957, n29956, n29955, n29954, 
            n29953, n29952, n29951, n29950, n29949, n29948, n29947, 
            n29946, n29945, n29944, n29943, n29942, n29941, n29940, 
            n29939, n43483, n29658, n29657, n29654, n29653, \Ki[0] , 
            n29652, \Kp[0] , n29626, n29625, n82, \FRAME_MATCHER.i_31__N_2624 , 
            n45660, \state[0] , \state[2] , \state[3] , n6935, n123, 
            n1, n29234, \r_SM_Main_2__N_3613[1] , r_SM_Main, \r_Bit_Index[0] , 
            tx_o, n44068, n29667, n29662, n51668, VCC_net, n20400, 
            n4_adj_6, tx_enable, n29246, r_Rx_Data, r_SM_Main_adj_14, 
            RX_N_10, \r_Bit_Index[0]_adj_10 , n44059, \r_SM_Main_2__N_3542[2] , 
            n27976, n4_adj_11, n29679, n29672, n43733, n29650, n29649, 
            n29648, n29647, n29646, n29645, n29644, n44138, n4_adj_12, 
            n4_adj_13, n27971, n35414) /* synthesis syn_module_defined=1 */ ;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[3] ;
    input CLK_c;
    input GND_net;
    input n29756;
    output [7:0]control_mode;
    output n25135;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[13] ;
    input n29755;
    output \FRAME_MATCHER.i_31__N_2622 ;
    input n29754;
    output \FRAME_MATCHER.state_31__N_2660[2] ;
    output \FRAME_MATCHER.i_31__N_2626 ;
    output n4452;
    output n7;
    output [7:0]rx_data;
    output n771;
    input n29753;
    input n29752;
    output n45880;
    output n3303;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[1] ;
    output n63;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[11] ;
    input n29751;
    input n29750;
    input n29749;
    output [23:0]PWMLimit;
    input n29748;
    output [7:0]\data_in_frame[8] ;
    output \FRAME_MATCHER.state[0] ;
    input n29747;
    output rx_data_ready;
    output [23:0]setpoint;
    input n29746;
    output [7:0]\data_in_frame[10] ;
    input n29745;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[13] ;
    input n29744;
    input n29743;
    input n29742;
    input n29741;
    input n29740;
    input n29739;
    input n29738;
    input n29737;
    input n29736;
    input n29735;
    input n29734;
    input n29733;
    input n29732;
    input n29731;
    input n29730;
    input n29729;
    input n29728;
    input n29727;
    input n51593;
    input n51594;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[20] ;
    output n14;
    output tx_active;
    output DE_c;
    output LED_c;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[5] ;
    output n25063;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[5] ;
    output n29310;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[24] ;
    output \data_out_frame[27][1] ;
    input [7:0]ID;
    output n4;
    output n29176;
    output n41916;
    input n30209;
    output [23:0]IntegralLimit;
    input n30208;
    input n30207;
    input n30206;
    input n30205;
    input n30204;
    input n30203;
    input n30202;
    input n30201;
    input n30200;
    input n30199;
    input n30198;
    input n30197;
    input n30196;
    input n30195;
    input n30194;
    input n30193;
    input n30192;
    input n30191;
    input n30190;
    input n30189;
    input n30188;
    input n30186;
    input n30185;
    input n30184;
    input n30183;
    input n30182;
    input n30181;
    input n30180;
    input n30179;
    input n30178;
    input n30177;
    input n30176;
    input n30175;
    input n30174;
    input n30173;
    input n30172;
    input n30171;
    input n30170;
    input n30169;
    input n30168;
    input n30167;
    input n30166;
    input n30165;
    input n30164;
    input n30163;
    input n30162;
    input n30161;
    input n30160;
    input n30159;
    input n30158;
    input n30157;
    input n30156;
    input n30155;
    input n30154;
    output \Kp[1] ;
    input n30153;
    output \Kp[2] ;
    input n30152;
    output \Kp[3] ;
    input n30151;
    output \Kp[4] ;
    input n30150;
    output \Kp[5] ;
    input n30149;
    output \Kp[6] ;
    input n30148;
    output \Kp[7] ;
    input n30147;
    output \Kp[8] ;
    input n30146;
    output \Kp[9] ;
    input n30145;
    output \Kp[10] ;
    input n30144;
    output \Kp[11] ;
    input n30143;
    output \Kp[12] ;
    input n30141;
    output \Kp[13] ;
    input n30140;
    output \Kp[14] ;
    input n30139;
    output \Kp[15] ;
    input n30138;
    output \Ki[1] ;
    input n30137;
    output \Ki[2] ;
    input n30136;
    output \Ki[3] ;
    input n30135;
    output \Ki[4] ;
    input n30134;
    output \Ki[5] ;
    input n30133;
    output \Ki[6] ;
    input n30132;
    output \Ki[7] ;
    input n30131;
    output \Ki[8] ;
    input n30130;
    output \Ki[9] ;
    input n30129;
    output \Ki[10] ;
    input n30128;
    output \Ki[11] ;
    input n30127;
    output \Ki[12] ;
    input n30126;
    output \Ki[13] ;
    input n30125;
    output \Ki[14] ;
    input n30124;
    output \Ki[15] ;
    input n30123;
    input n30122;
    input n30121;
    input n30120;
    input n30119;
    input n30118;
    input n30117;
    input n30116;
    input n30115;
    input n30114;
    input n30113;
    input n30112;
    input n30111;
    input n30110;
    input n30109;
    input n30108;
    input n30107;
    input n30106;
    input n30105;
    input n30104;
    input n30103;
    input n30102;
    input n30101;
    input n30100;
    input n30099;
    input n30098;
    input n30097;
    input n30096;
    input n30095;
    input n30094;
    input n30093;
    input n30092;
    input n30091;
    input n30090;
    input n30089;
    input n30088;
    input n30087;
    input n30086;
    input n30085;
    input n30084;
    input n30083;
    input n30082;
    input n30081;
    input n30080;
    input n30079;
    input n30078;
    input n30077;
    input n30076;
    input n30075;
    input n30074;
    input n30073;
    input n30072;
    input n30071;
    input n30070;
    input n30069;
    input n30068;
    input n30067;
    input n30066;
    input n30065;
    input n30064;
    input n30063;
    input n30062;
    input n30061;
    input n30060;
    input n30059;
    input n30058;
    input n30057;
    input n30056;
    input n30055;
    input n30054;
    input n30053;
    input n30052;
    input n30051;
    input n30050;
    input n30049;
    input n30048;
    input n30047;
    input n30046;
    input n30045;
    input n30044;
    input n30043;
    input n30042;
    input n30041;
    input n30040;
    input n30039;
    input n30038;
    input n30037;
    input n30036;
    input n30035;
    input n30034;
    input n30033;
    input n30032;
    input n30031;
    input n30030;
    input n30029;
    input n30028;
    input n30027;
    input n30026;
    input n30025;
    input n30024;
    input n30023;
    input n30022;
    input n30021;
    input n30020;
    input n30019;
    input n30018;
    input n30017;
    input n30016;
    input n30015;
    input n30014;
    input n30013;
    input n30012;
    input n30011;
    input n30009;
    input n30008;
    input n30007;
    input n30006;
    input n30005;
    input n30004;
    input n30003;
    input n30002;
    input n30001;
    input n30000;
    input n29999;
    input n29998;
    input n29997;
    input n29996;
    input n29995;
    input n29994;
    input n29993;
    input n29992;
    input n29991;
    input n29990;
    input n29989;
    input n29988;
    input n29987;
    input n29986;
    input n29985;
    input n29984;
    input n29983;
    input n29982;
    input n29981;
    input n29980;
    input n29979;
    input n29978;
    input n29977;
    input n29976;
    input n29975;
    input n29974;
    input n29973;
    input n29972;
    input n29971;
    input n29970;
    input n29969;
    input n29968;
    input n29967;
    input n29966;
    input n29965;
    input n29964;
    input n29963;
    input n29962;
    input n29961;
    output [23:0]neopxl_color;
    input n29960;
    input n29959;
    input n29958;
    input n29957;
    input n29956;
    input n29955;
    input n29954;
    input n29953;
    input n29952;
    input n29951;
    input n29950;
    input n29949;
    input n29948;
    input n29947;
    input n29946;
    input n29945;
    input n29944;
    input n29943;
    input n29942;
    input n29941;
    input n29940;
    input n29939;
    input n43483;
    input n29658;
    input n29657;
    input n29654;
    input n29653;
    output \Ki[0] ;
    input n29652;
    output \Kp[0] ;
    input n29626;
    input n29625;
    output n82;
    output \FRAME_MATCHER.i_31__N_2624 ;
    output n45660;
    input \state[0] ;
    input \state[2] ;
    input \state[3] ;
    output n6935;
    output n123;
    output n1;
    output n29234;
    output \r_SM_Main_2__N_3613[1] ;
    output [2:0]r_SM_Main;
    output \r_Bit_Index[0] ;
    output tx_o;
    output n44068;
    input n29667;
    input n29662;
    input n51668;
    input VCC_net;
    output n20400;
    output n4_adj_6;
    output tx_enable;
    output n29246;
    output r_Rx_Data;
    output [2:0]r_SM_Main_adj_14;
    input RX_N_10;
    output \r_Bit_Index[0]_adj_10 ;
    output n44059;
    output \r_SM_Main_2__N_3542[2] ;
    output n27976;
    output n4_adj_11;
    input n29679;
    input n29672;
    input n43733;
    input n29650;
    input n29649;
    input n29648;
    input n29647;
    input n29646;
    input n29645;
    input n29644;
    input n44138;
    output n4_adj_12;
    output n4_adj_13;
    output n27971;
    output n35414;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire Kp_23__N_988;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n29060, n29764;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n29763, n29762, n29761, n29760, n29759, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n2_adj_4211, n39171, n2987, n29758, n29757, n13, 
        n45062;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    wire [31:0]\FRAME_MATCHER.state_31__N_2724 ;
    
    wire n44384;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n48882, n48881, n39172, n4_c, n48504;
    wire [7:0]n8825;
    
    wire n31447, n44825, n2_adj_4212, n39170, n44293, Kp_23__N_974, 
        n44602, n29017, n8, n44156;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n29781, n5, n36241, n6, tx_transmit_N_3513, n27958, n4_adj_4213, 
        n35517, \FRAME_MATCHER.i_31__N_2623 , n31443, n45036, \FRAME_MATCHER.i_31__N_2621 , 
        n2_adj_4214, n39169, n8_adj_4215, n27981, n8_adj_4216, n44134, 
        n29782, n44, n42, n43, n41, n40, n39, n50, n45, n27841, 
        n8_adj_4217, n28032, n20, n27838, n19, n48641, n14_c, 
        n28038, n15, n16, n17, n27968, n10, n14_adj_4218, n9, 
        n18, n20_adj_4219, n15_adj_4220, n63_adj_4221, n16_adj_4222, 
        n17_adj_4223, n63_adj_4224, n20372, n29783, n48848, n48849, 
        n35182, n44163, n29784, n29785, n29786, n29787, n31, n25324, 
        n35205, n44786, n44584, n16_adj_4225, n18_adj_4226, n44596, 
        n44831, n17_adj_4227, n42452;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n24, Kp_23__N_1217, n9_adj_4228, n46131, n41577, n28, n28428, 
        n28837, n28342, n28749, n26, n28313, n28319, n28347, n27, 
        n28736, n28719, n28630, n4_adj_4229, n25, n31_adj_4230, 
        n24773, n36381, n98, n12, n36247, n36029, n29187, n48843, 
        n48842, n48851, n48852;
    wire [0:0]n5426;
    wire [2:0]r_SM_Main_2__N_3616;
    
    wire n44882, \FRAME_MATCHER.rx_data_ready_prev , n48813, n48812, 
        n48854, n48855, n6560, n48753, n48752, n48857, n29788, 
        n48858, n48864, n48863, n6_adj_4231, n48869, n48870, n48723, 
        n48722, n48872, n48873, n48720, n48719, n44444, n44837, 
        n44427, n44684, n36087, n70, n35343, n44367, n28675, n44703, 
        n44553, n44765, n42380;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n8_adj_4232, n35184, n7_adj_4233, n36505, n8_adj_4234, n44431, 
        n44852, n44777, n28445, n16_adj_4235, n17_adj_4236, n49730, 
        n49729, n16_adj_4237, n17_adj_4238, n49727, n49726, n16_adj_4240, 
        n7_adj_4241, n17_adj_4242, n49724, n49723, n2_adj_4243, n39168, 
        n16_adj_4244, n17_adj_4245, n49721, n49720, n2_adj_4246, n39167, 
        n16_adj_4247, n17_adj_4248, n49718, n49717, n16_adj_4249, 
        n2_adj_4250, n39166, n17_adj_4251, n49712, n49711, n2_adj_4252, 
        n39165, n16_adj_4253, n17_adj_4254, n49709, n49708, n16_adj_4255, 
        n17_adj_4256, n49706, n49705, n2_adj_4257, n39164, n28612, 
        n10_adj_4258, n2_adj_4259, n39163, n44393, n27601, n6_adj_4260, 
        n88, n46735, n46530, n29452, n46541, n46485, n2_adj_4261, 
        n39162, n48780, n48781, n48779, n28618, n51528, n49728, 
        n6583, n2_adj_4262, n39161, n6582, n6581, n6580, n6579, 
        n6578, n6577, n6576, n6575, n6574, n6573, n6572, n6571, 
        n6570, n6569, n6568, n6567, n6566, n6565, n6564, n6563, 
        n48823, n6562, n48821, n6561, n43669, n43539, n169, Kp_23__N_1426, 
        n44700;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n8_adj_4263, n41670, n10_adj_4264, n46645, n41549, n42122, 
        n44521, n44447, n6_adj_4265, n42345, n44424, n28235, n44505, 
        n44756, n2_adj_4266, n39160;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n10_adj_4267, n44846;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n14_adj_4268, n42356, n46063, n44818;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n44569, n44572, n28941, n44530, n42368, n42408, n44780, 
        n44540, n28264, n44774, n46396, n42341, n10_adj_4269, n27552, 
        n44671, n28796, n12_adj_4270, n41819, n28160, n44410, n38, 
        n44252, n52, n56, n44544, n44524, n44364, n54, n44279, 
        n55, n44849, n44637, n44792, n53, n44486, n50_adj_4271, 
        n44578, n58, n62, n44346, n49, n2_adj_4272, n39159, n42347, 
        n14_adj_4273, n15_adj_4274, Kp_23__N_1536, n42343, n44599, 
        n44611, n44205, n24_adj_4275, n44664, n44224, n42413, n22, 
        n18_adj_4276, n26_adj_4277, n28289, n44759, n28655, n6_adj_4278, 
        n44233, n44810, n41622, n29057, n8_adj_4279, n44325, Kp_23__N_1228, 
        n44716, n44587, n20_adj_4280, n44399, n44658, n19_adj_4281, 
        n44316, n28624, n21, Kp_23__N_1306, n43667, n43543, n44246, 
        n41553, n42082, n14_adj_4282, n44337, n15_adj_4283, n44413, 
        n44208, n28171, n44349, n28_adj_4284, n32, n43665, n43547, 
        n43663, n43551, n43661, n43555, n7_adj_4285, n8_adj_4286, 
        n43659, n43559, n7_adj_4287, n8_adj_4288, n43657, n43563, 
        n43655, n43567, n43653, n43571, n35190, n36044, n43651, 
        n43575, n43649, n43579, n43647, n43583, n7_adj_4289, n8_adj_4290, 
        n43645, n43587, n43643, n43591, n43641, n43595, n43639, 
        n43513, n44236, n30, n31_adj_4291, n29, n28890, n28494, 
        n6_adj_4292, n43637, n43505, n43635, n43493, n42398, n43633, 
        n43599, n43631, n43509, n43629, n43603, n43627, n43607, 
        n43625, n43611, n43623, n43489, n43485, n43691, n44547, 
        n6_adj_4293, n44813, n28705, n44453, n44652, n10_adj_4294, 
        n2_adj_4295, n39158, Kp_23__N_981, n28840, n46112;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n44713, n44789, n45837, n45838, n45552, n45583, n44577, 
        n28794, n45554;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n46786, n45780, n46761, n46120, n45896, n46218, n46058, 
        n44227, n10_adj_4296, Kp_23__N_977, Kp_23__N_993, n44402, 
        Kp_23__N_1096, n44396, n6_adj_4297, n28843, n28114, n10_adj_4298, 
        n51372, n49725, n51567, n51468, n7_adj_4299;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n51378, n49722, n51561, n51462, n7_adj_4300, n51384, n49719, 
        n51555, n51456, n7_adj_4301, n51390, n49713, n51549, n51450, 
        n7_adj_4302, n51396, n49710, n51543, n51444, n7_adj_4303, 
        n51402, n49707, n51537, n51438, n7_adj_4304, n51408, n49704, 
        n51531, n2_adj_4305, n3_adj_4306, n2_adj_4307, n3_adj_4308, 
        n2_adj_4309, n3_adj_4310, n2_adj_4311, n3_adj_4312, n3_adj_4313, 
        n3_adj_4314, n3_adj_4315, n3_adj_4316, n3_adj_4317, n3_adj_4318, 
        n3_adj_4319, n3_adj_4320, n3_adj_4321, n3_adj_4322, n3_adj_4323, 
        n3_adj_4324, n3_adj_4325, n3_adj_4326, n2_adj_4327, n3_adj_4328, 
        n2_adj_4329, n3_adj_4330, n2_adj_4331, n3_adj_4332, n2_adj_4333, 
        n3_adj_4334, n2_adj_4335, n3_adj_4336, n2_adj_4337, n3_adj_4338, 
        n2_adj_4339, n3_adj_4340, n2_adj_4341, n3_adj_4342, n2_adj_4343, 
        n3_adj_4344, n2_adj_4345, n3_adj_4346, n2_adj_4347, n3_adj_4348, 
        n2_adj_4349, n3_adj_4350, n2_adj_4351, n3_adj_4352, n44690, 
        n44239, n44306, n39157, n28238, n44834, n44199, n44741, 
        n44495, n28615, n28156, n10_adj_4353, n28204, n39156, n44352, 
        n39155, n26_adj_4354, n36, n44256, n34, n44605, n40_adj_4355, 
        n38_adj_4356, n39_adj_4357, n37, Kp_23__N_1020, n44482, n6_adj_4358, 
        n39154, n51432, n7_adj_4359, n51525, n51519, n51522, n51513, 
        n51516, n51507, n51510, n51501, n51504, n51495, n51498, 
        n51489, n51492, n51483, n51486, n51366, n51477, n51426, 
        n7_adj_4360, n44622, n10_adj_4361, n44744, n44608, n14_adj_4362, 
        n28753, n39153, n44416, n12_adj_4363, n44355, n41565, n46102, 
        n39152, n44218, n6_adj_4364, n39151, n44296, n12_adj_4365, 
        n39150, n6_adj_4366, n28349, n28716, n44343, n28956, n10_adj_4367, 
        n44771, n48817, n190, n44183, n12_adj_4368, n10_adj_4369, 
        n11, n48815, n9_adj_4370, n8_adj_4371, n44661, n16_adj_4372, 
        n18_adj_4373, n48807, n48808, n48806, n6_adj_4374, n14_adj_4375, 
        n46262, n48801, n48802, n48800, n6_adj_4376, n16_adj_4377, 
        n17_adj_4378;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n8_adj_4379, n46883, n13_adj_4380, n16_adj_4381, n48795, 
        n48796, n12_adj_4382, n10_adj_4383, n14_adj_4384, n46244, 
        n10_adj_4385, n6_adj_4386, n46339, n12_adj_4387, n13_adj_4388, 
        n12_adj_4389, n48794, n46324, n48581, n48789, n48790, n48788, 
        n11_adj_4390, n46425, n22_adj_4391, n28_adj_4392, n46724, 
        n6_adj_4393, n48784, n12_adj_4394, n45599, n6_adj_4395, n46374, 
        n48782, n39149, n45835, n46136, n48583, n48585, n30_adj_4396, 
        n25_adj_4397, n39148, n188, n39147, n39146, n39145, n161, 
        n51465, n51459, n51453, n51447, n51441, n27874, n44408, 
        n44722, n44456, n44390, n44498, n28588, n12_adj_4399, n45883, 
        n44753, n45973, n41591, n44312, n14_adj_4400, n44710, n44640, 
        n15_adj_4401, n42428, n28583, n44489, n44437, n8_adj_4402, 
        n29773, n44434, n6_adj_4403, n41584, n28856, n51435, n29774, 
        n28849, n28855, n41638, n29775, n27608, n44340, n28096, 
        n44643, n29776, n14_adj_4404, n29777, n10_adj_4405, n29778, 
        n8_adj_4406, n29779, n41575, n27564, n42364, n18_adj_4407, 
        n42394, n44494, n44590, n20_adj_4408, n44550, n15_adj_4409, 
        n42403, n46040, n44518, n41659, n28468, n44282, n10_adj_4410, 
        n44798, n44707, n6_adj_4411, n41655, n44373, n44768, n26_adj_4412, 
        n44750, n29_adj_4413, n41571, n27722, n28_adj_4414, n32_adj_4415, 
        n44581, n26118, n28646, n27_adj_4416, n44215, n7_adj_4417, 
        n8_adj_4418, n29780, n27588, n41601, n27652, n42439, n10_adj_4419, 
        n46263, n44533, n41331, n41611, n6_adj_4420, n8_adj_4421, 
        n29765, n46085, n29766, n46780, n28776, n42360, n44565, 
        n28201, n28490, n44361, n12_adj_4422, n51429, n44655, n44287, 
        n44463, n12_adj_4423, n28884, n44728, n29767, n44628, n10_adj_4424, 
        n44271, n10_adj_4425, n14_adj_4426, n18_adj_4427, n44450, 
        n44631, n10_adj_4428, n44387, n44242, n6_adj_4429, n44319, 
        n44646, n29768, n44512, n28392, n27665, n26043, n41609, 
        n29931, n29930, n44840, n29929, n29928, n44804, n44290, 
        n10_adj_4430, n4_adj_4431, n103, n29769, n44843, n15_adj_4432, 
        n14_adj_4433, n28658, n48837, n48836, n48884, n48885, n51423, 
        n48834, n48833, n29770, n44719, n29656, n29927, n44221, 
        n44405, n12_adj_4434, n29926, n29925, n29924, n29923, n29922, 
        n29921, n29920, n29919, n29918, n29917, n29916, n29915, 
        n29914, n29913, n29912, n29911, n29910, n29909, n29908, 
        n29907, n29906, n29905, n29904, n29903, n29902, n29901, 
        n29900, n29899, n29898, n29897, n29771, n46787, n29772, 
        n44687, n1519, n28078, n29896, n29895, n29894, n29893, 
        n29892, n29891, n29890, n29889, n29888, n29887, n29886, 
        n29885, n29884, n29883, n29882, n29881, n29880, n29879, 
        n29878, n29877, n29876, n29875, n29874, n29873, n29872, 
        n29871, n29870, n29869, n29868, n29867, n29866, n29865, 
        n29864, n29863, n29862, n29861, n29860, n29859, n29858, 
        n29857, n29856, n29855, n29854, n29853, n29852, n29851, 
        n29850, n29849, n29848, n29847, n29846, n29845, n29844, 
        n29843, n29842, n29841, n29840, n29839, n29838, n29837, 
        n29836, n29835, n29834, n29833, n29832, n29831, n29830, 
        n29829, n29828, n29827, n29826, n29825, n29824, n29823, 
        n29822, n29821, n29820, n29819, n29818, n29817, n29816, 
        n29815, n29814, n29813, n29812, n29811, n29810, n29809, 
        n29808, n29807, n29806, n29805, n29804, n29803, n29802, 
        n29801, n29800, n29799, n29798, n29797, n29796, n29795, 
        n29794, n29793, n29792, n29791, n29790, n29789, n44169, 
        n30_adj_4435, n28874, n44556, n34_adj_4436, n41545, n32_adj_4437, 
        n44249, n44334, n42180, n33, n28531, n44309, n1516, n44807, 
        n31_adj_4438, n46648, n22_adj_4439, n44625, n21_adj_4440, 
        n41791, n14_adj_4441, n23, n15_adj_4442, n28713, n19_adj_4443, 
        n44725, n44559, n22_adj_4444, n44509, n18_adj_4445, n44731, 
        n10_adj_4446, n44259, n44828, n44502, n14_adj_4447, n10_adj_4448, 
        n41541, n28141, n45757, n44492, n44795, n44615, n44230, 
        n44473, n44265, n42433, n6_adj_4449, n39182, n44537, n24_adj_4450, 
        n39181, n41636, n41940, n39180, n10_adj_4451, n22_adj_4452, 
        n39179, n26_adj_4453, n39178, n10_adj_4454, n1510, n1513, 
        n39177, n39176, n10_adj_4455, n44459, n27572, n28388, n14_adj_4456, 
        n44380, n27866, n4_adj_4457, n8_adj_4458, n39175, n39174, 
        n39173, n44696, n44681, n15_adj_4459, n44268, n14_adj_4460, 
        n44735, n1673, n10_adj_4461, n41531, n44693, n44420, n1191, 
        n28041, n31_adj_4462, n44634, n44262, n14_adj_4463, n10_adj_4464, 
        n44649, n44322, n29039, n6_adj_4465, n25_adj_4466, n8_adj_4467, 
        n29054, n44476, n44470, n10_adj_4468, n28045, n6_adj_4469, 
        n10_adj_4470, n51405, n29027, n52_adj_4471, n44678, n50_adj_4472, 
        n28104, n51, n49_adj_4473, n32_adj_4474, n44328, n48, n44668, 
        n47, n58_adj_4475, n53_adj_4476, n27574, n41523, n44377, 
        n10_adj_4477, n103_adj_4478, n4_adj_4479, n51399, n44738, 
        n44358, n12_adj_4480, n15_adj_4481, n12_adj_4482, n28805, 
        n12_adj_4483, n14_adj_4484, n10_adj_4485, n12_adj_4486, n44762, 
        n45615, n44186, n45105, n44062, n51393, n44176, n11_adj_4487, 
        n51387, n1_c, n44331, n44934, n28904, n2_adj_4488, n51381, 
        n51375, n51369, n51363, n18_adj_4490, n21_adj_4491, n20_adj_4492, 
        n30_adj_4493, n28_adj_4494, n29_adj_4495, n27_adj_4496, n45066, 
        n15_adj_4497, n4_adj_4498, n45024, n45517;
    
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_988), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[0] [6]), .O(n29060));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n29764));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n29763));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n29762));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n29761));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n29760));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n29759));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_29_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n39171), .O(n2_adj_4211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n29758));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n29757));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n29756));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut (.I0(n13), .I1(n45062), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state_31__N_2724 [3]), .O(n25135));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_988), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [7]), .O(n44384));   // verilog/coms.v(70[16:27])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33445_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48882));
    defparam i33445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33444_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48881));
    defparam i33444_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_29 (.CI(n39171), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n39172));
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n29755));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33140_3_lut_4_lut (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [6]), .I3(n4_c), .O(n48504));   // verilog/coms.v(77[16:27])
    defparam i33140_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n31447), .D(n8825[1]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
            .E(n31447), .D(n8825[2]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
            .E(n31447), .D(n8825[3]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
            .E(n31447), .D(n8825[4]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n29754));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n44825));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_28_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n39170), .O(n2_adj_4212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_28 (.CI(n39170), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n39171));
    SB_LUT4 i2_3_lut_4_lut_adj_870 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [5]), .I3(n44293), .O(Kp_23__N_988));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_871 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [4]), .I3(Kp_23__N_974), .O(n44602));
    defparam i2_3_lut_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 select_650_Select_2_i7_3_lut (.I0(\FRAME_MATCHER.state_31__N_2660[2] ), 
            .I1(\FRAME_MATCHER.i_31__N_2626 ), .I2(n4452), .I3(GND_net), 
            .O(n7));
    defparam select_650_Select_2_i7_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_3_lut_adj_872 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n29017));
    defparam i1_2_lut_3_lut_adj_872.LUT_INIT = 16'h9696;
    SB_LUT4 i16254_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n29781));
    defparam i16254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21949_4_lut (.I0(n5), .I1(\FRAME_MATCHER.i [31]), .I2(\FRAME_MATCHER.i [2]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i21949_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i35219_2_lut (.I0(n36241), .I1(n6), .I2(GND_net), .I3(GND_net), 
            .O(tx_transmit_N_3513));
    defparam i35219_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n27958), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4213));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i17917_4_lut (.I0(n35517), .I1(\FRAME_MATCHER.i_31__N_2623 ), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n4_adj_4213), .O(n31443));   // verilog/coms.v(112[11:16])
    defparam i17917_4_lut.LUT_INIT = 16'hc5c0;
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n29753));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n45036), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2621 ));   // verilog/coms.v(127[12] 300[6])
    defparam i2_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_43_27_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n39169), .O(n2_adj_4214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n29752));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_27 (.CI(n39169), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n39170));
    SB_LUT4 i21953_4_lut (.I0(n8_adj_4215), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27981), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i21953_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i3_3_lut (.I0(\FRAME_MATCHER.i_31__N_2622 ), .I1(\FRAME_MATCHER.i_31__N_2621 ), 
            .I2(n31443), .I3(GND_net), .O(n8_adj_4216));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n8_adj_4216), .I2(n2987), 
            .I3(n44134), .O(n45880));
    defparam i4_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i16255_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n29782));
    defparam i16255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n27981));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_873 (.I0(\FRAME_MATCHER.i [4]), .I1(n27981), .I2(GND_net), 
            .I3(GND_net), .O(n27841));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_873.LUT_INIT = 16'heeee;
    SB_LUT4 i21950_4_lut (.I0(n8_adj_4217), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n27841), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i21950_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i8_4_lut (.I0(\data_in[2] [6]), .I1(\data_in[2] [0]), .I2(n28032), 
            .I3(\data_in[0] [5]), .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut (.I0(n27838), .I1(\data_in[3] [7]), .I2(\data_in[1] [6]), 
            .I3(\data_in[2] [5]), .O(n19));
    defparam i7_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33276_4_lut (.I0(\data_in[1] [2]), .I1(\data_in[1] [3]), .I2(\data_in[0] [1]), 
            .I3(\data_in[3] [2]), .O(n48641));
    defparam i33276_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i11_3_lut (.I0(n48641), .I1(n19), .I2(n20), .I3(GND_net), 
            .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i5_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[2] [4]), .I2(\data_in[3] [0]), 
            .I3(GND_net), .O(n14_c));
    defparam i5_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut (.I0(\data_in[1] [4]), .I1(\data_in[0] [6]), .I2(n28038), 
            .I3(\data_in[1] [5]), .O(n15));
    defparam i6_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_874 (.I0(n15), .I1(\data_in[1] [0]), .I2(n14_c), 
            .I3(\data_in[2] [2]), .O(n27838));
    defparam i8_4_lut_adj_874.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_875 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16));
    defparam i6_4_lut_adj_875.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_876 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17));
    defparam i7_4_lut_adj_876.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_in[1] [6]), .I2(n16), .I3(\data_in[3] [7]), 
            .O(n27968));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_877 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10));
    defparam i4_4_lut_adj_877.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_878 (.I0(\data_in[3] [4]), .I1(n10), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n28038));
    defparam i5_3_lut_adj_878.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_879 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4218));
    defparam i6_4_lut_adj_879.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_880 (.I0(\data_in[3] [5]), .I1(\data_in[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n9));
    defparam i1_2_lut_adj_880.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_881 (.I0(n9), .I1(n14_adj_4218), .I2(\data_in[3] [6]), 
            .I3(\data_in[2] [1]), .O(n28032));
    defparam i7_4_lut_adj_881.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_882 (.I0(\data_in[2] [4]), .I1(n28032), .I2(\data_in[1] [5]), 
            .I3(n28038), .O(n18));
    defparam i7_4_lut_adj_882.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_883 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n27968), .O(n20_adj_4219));
    defparam i9_4_lut_adj_883.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4220));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n15_adj_4220), .I1(n20_adj_4219), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_adj_4221));
    defparam i10_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_884 (.I0(\data_in[3] [6]), .I1(n27838), .I2(\data_in[2] [1]), 
            .I3(\data_in[0] [7]), .O(n16_adj_4222));
    defparam i6_4_lut_adj_884.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_885 (.I0(n27968), .I1(\data_in[3] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[2] [3]), .O(n17_adj_4223));
    defparam i7_4_lut_adj_885.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_886 (.I0(n17_adj_4223), .I1(\data_in[3] [1]), .I2(n16_adj_4222), 
            .I3(\data_in[3] [5]), .O(n63_adj_4224));
    defparam i9_4_lut_adj_886.LUT_INIT = 16'hfbff;
    SB_LUT4 i6990_2_lut (.I0(n63), .I1(n771), .I2(GND_net), .I3(GND_net), 
            .O(n20372));   // verilog/coms.v(157[6] 159[9])
    defparam i6990_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16256_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n29783));
    defparam i16256_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33411_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48848));
    defparam i33411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33412_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48849));
    defparam i33412_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n29751));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n29750));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n29749));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_887 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n35182), .O(n44163));
    defparam i2_3_lut_4_lut_adj_887.LUT_INIT = 16'hf7ff;
    SB_LUT4 i16257_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n29784));
    defparam i16257_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16258_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n29785));
    defparam i16258_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16259_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n29786));
    defparam i16259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n29748));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16260_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n29787));
    defparam i16260_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21695_2_lut (.I0(n31), .I1(n25324), .I2(GND_net), .I3(GND_net), 
            .O(n35205));
    defparam i21695_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_888 (.I0(n4_c), .I1(\data_in_frame[8] [1]), .I2(n44786), 
            .I3(n44584), .O(n16_adj_4225));
    defparam i6_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(\data_in_frame[3] [6]), .I1(n16_adj_4225), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(n18_adj_4226));
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_889 (.I0(\data_in_frame[3] [5]), .I1(n44596), .I2(n44831), 
            .I3(n29017), .O(n17_adj_4227));
    defparam i7_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_890 (.I0(n17_adj_4227), .I1(n42452), .I2(n18_adj_4226), 
            .I3(\data_in_frame[7] [7]), .O(n24));
    defparam i8_4_lut_adj_890.LUT_INIT = 16'hde7b;
    SB_LUT4 equal_2054_i9_2_lut (.I0(Kp_23__N_1217), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4228));   // verilog/coms.v(236[9:81])
    defparam equal_2054_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut (.I0(n46131), .I1(n24), .I2(n41577), .I3(\data_in_frame[8] [0]), 
            .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hdfef;
    SB_LUT4 i10_4_lut_adj_891 (.I0(n28428), .I1(n28837), .I2(n28342), 
            .I3(n28749), .O(n26));
    defparam i10_4_lut_adj_891.LUT_INIT = 16'hffef;
    SB_LUT4 i11_4_lut (.I0(n28313), .I1(n9_adj_4228), .I2(n28319), .I3(n28347), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_892 (.I0(n28736), .I1(n28719), .I2(n28630), .I3(n4_adj_4229), 
            .O(n25));
    defparam i9_4_lut_adj_892.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_893 (.I0(n25), .I1(n27), .I2(n26), .I3(n28), 
            .O(n31));
    defparam i15_4_lut_adj_893.LUT_INIT = 16'hfffe;
    SB_LUT4 i8103_3_lut (.I0(n31_adj_4230), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n24773));   // verilog/coms.v(145[4] 299[11])
    defparam i8103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(n25324), .I1(n36381), .I2(n98), .I3(n24773), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i35203_4_lut (.I0(n36247), .I1(n12), .I2(n36029), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n29187));
    defparam i35203_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i33406_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48843));
    defparam i33406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33405_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48842));
    defparam i33405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33414_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48851));
    defparam i33414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33415_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48852));
    defparam i33415_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n29747));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
            .E(n31447), .D(n8825[5]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3616[0]), .C(CLK_c), .D(n5426[0]), 
            .R(n44882));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33376_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48813));
    defparam i33376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33375_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48812));
    defparam i33375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33417_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48854));
    defparam i33417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33418_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48855));
    defparam i33418_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n29187), .D(n6560));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33316_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48753));
    defparam i33316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33315_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48752));
    defparam i33315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33420_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48857));
    defparam i33420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16261_3_lut_4_lut (.I0(n8), .I1(n44156), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n29788));
    defparam i16261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n29746));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33421_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48858));
    defparam i33421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33427_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48864));
    defparam i33427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33426_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48863));
    defparam i33426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_894 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[10] [3]), .I3(GND_net), .O(n6_adj_4231));
    defparam i1_2_lut_3_lut_adj_894.LUT_INIT = 16'h9696;
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n29745));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33432_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48869));
    defparam i33432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33433_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48870));
    defparam i33433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33286_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48723));
    defparam i33286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33285_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48722));
    defparam i33285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33435_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48872));
    defparam i33435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33436_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48873));
    defparam i33436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33283_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48720));
    defparam i33283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33282_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48719));
    defparam i33282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_895 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[8] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n44444));
    defparam i1_2_lut_3_lut_adj_895.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_896 (.I0(\data_in_frame[11] [1]), .I1(n44837), 
            .I2(\data_in_frame[10] [7]), .I3(\data_in_frame[13] [3]), .O(n44427));
    defparam i2_3_lut_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n29744));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
            .E(n31447), .D(n8825[6]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n29743));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n29742));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n29741));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n29740));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n29739));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
            .E(n31447), .D(n8825[7]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2660_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4215));
    defparam i2660_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n29738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n29737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n29736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n29735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n29734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n29733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n29732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n29731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n29730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n29729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n29728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n29727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(CLK_c), 
           .D(n51593));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(CLK_c), 
           .D(n51594));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_897 (.I0(\data_in_frame[9] [0]), .I1(n28736), 
            .I2(\data_in_frame[9] [7]), .I3(GND_net), .O(n44684));
    defparam i1_2_lut_3_lut_adj_897.LUT_INIT = 16'h9696;
    SB_LUT4 i22571_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n36087));
    defparam i22571_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n36087), .I3(byte_transmit_counter[2]), .O(n36241));
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i2_3_lut (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n6));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n70));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h8888;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
            .E(n31447), .D(n8825[0]), .R(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_899 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n35343));
    defparam i1_2_lut_adj_899.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_900 (.I0(\data_in_frame[9] [0]), .I1(n28736), 
            .I2(n28428), .I3(GND_net), .O(n44367));
    defparam i1_2_lut_3_lut_adj_900.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_901 (.I0(n28675), .I1(n44703), .I2(n44553), 
            .I3(n44765), .O(n42380));
    defparam i2_3_lut_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut (.I0(n28675), .I1(n44703), .I2(\data_in_frame[13] [5]), 
            .I3(\data_in_frame[16] [0]), .O(n8_adj_4232));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_902 (.I0(n36241), .I1(n35184), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4233));
    defparam i2_2_lut_adj_902.LUT_INIT = 16'heeee;
    SB_LUT4 mux_1330_i1_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n7_adj_4233), 
            .I2(n36505), .I3(n8_adj_4234), .O(n5426[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_1330_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i1_2_lut_3_lut_adj_903 (.I0(\data_in_frame[11] [4]), .I1(n44431), 
            .I2(n44852), .I3(GND_net), .O(n44777));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_904 (.I0(\data_in_frame[11] [4]), .I1(n44431), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n44703));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_904.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_905 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n28445));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_905.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4235));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4236));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34434_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49730));
    defparam i34434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34432_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49729));
    defparam i34432_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4237));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4238));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_906 (.I0(tx_transmit_N_3513), .I1(n35184), 
            .I2(\FRAME_MATCHER.i_31__N_2623 ), .I3(GND_net), .O(n14));   // verilog/coms.v(213[6] 220[9])
    defparam i1_2_lut_3_lut_adj_906.LUT_INIT = 16'he0e0;
    SB_LUT4 i34465_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49727));
    defparam i34465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34467_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49726));
    defparam i34467_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4240));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21675_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), .I2(GND_net), 
            .I3(GND_net), .O(n35184));
    defparam i21675_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_907 (.I0(\FRAME_MATCHER.state [3]), .I1(n7_adj_4241), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2622 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4242));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34468_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49724));
    defparam i34468_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34470_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49723));
    defparam i34470_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_43_26_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n39168), .O(n2_adj_4243)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4244));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n35184), .I1(\FRAME_MATCHER.i_31__N_2622 ), .I2(\FRAME_MATCHER.i_31__N_2623 ), 
            .I3(GND_net), .O(n31447));
    defparam i1_3_lut.LUT_INIT = 16'hdcdc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4245));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34472_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49721));
    defparam i34472_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34474_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49720));
    defparam i34474_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_26 (.CI(n39168), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n39169));
    SB_LUT4 add_43_25_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n39167), .O(n2_adj_4246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4247));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4248));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_25 (.CI(n39167), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n39168));
    SB_LUT4 i34475_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49718));
    defparam i34475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34387_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49717));
    defparam i34387_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4249));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_24_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n39166), .O(n2_adj_4250)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n39166), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n39167));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4251));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34478_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49712));
    defparam i34478_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34480_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49711));
    defparam i34480_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_43_23_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n39165), .O(n2_adj_4252)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4253));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4254));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34481_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49709));
    defparam i34481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34483_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49708));
    defparam i34483_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4255));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4256));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34484_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49706));
    defparam i34484_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34486_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49705));
    defparam i34486_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_23 (.CI(n39165), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n39166));
    SB_LUT4 add_43_22_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n39164), .O(n2_adj_4257)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(n28612), .I3(n10_adj_4258), .O(Kp_23__N_1217));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_43_22 (.CI(n39164), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n39165));
    SB_LUT4 add_43_21_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n39163), .O(n2_adj_4259)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_908 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n44393));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_908.LUT_INIT = 16'h9696;
    SB_CARRY add_43_21 (.CI(n39163), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n39164));
    SB_LUT4 i1_2_lut_3_lut_adj_909 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(n27601), .I3(GND_net), .O(n6_adj_4260));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_909.LUT_INIT = 16'h9696;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(CLK_c), .E(n46735), .D(n88), 
            .R(n46530));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR LED_3874 (.Q(LED_c), .C(CLK_c), .E(n46541), .D(n29452), 
            .R(n46485));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_20_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n39162), .O(n2_adj_4261)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n39162), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n39163));
    SB_LUT4 i33343_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48780));
    defparam i33343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33344_4_lut (.I0(n48780), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48781));
    defparam i33344_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i33342_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48779));
    defparam i33342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_910 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n28618));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_910.LUT_INIT = 16'h9696;
    SB_LUT4 i34466_2_lut (.I0(n51528), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49728));
    defparam i34466_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n29187), .D(n6583));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_19_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n39161), .O(n2_adj_4262)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n29187), .D(n6582));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n29187), .D(n6581));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n29187), .D(n6580));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n29187), .D(n6579));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n29187), .D(n6578));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n29187), .D(n6577));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n29187), .D(n6576));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n29187), .D(n6575));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n29187), .D(n6574));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n29187), .D(n6573));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n29187), .D(n6572));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n29187), .D(n6571));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n29187), .D(n6570));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n29187), .D(n6569));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n29187), .D(n6568));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n29187), .D(n6567));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n29187), .D(n6566));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n29187), .D(n6565));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n29187), .D(n6564));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n29187), .D(n6563));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33386_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n48823));
    defparam i33386_4_lut.LUT_INIT = 16'hec2c;
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n29187), .D(n6562));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33384_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48821));
    defparam i33384_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n29187), .D(n6561));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(CLK_c), 
            .D(n43669), .S(n43539));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_19 (.CI(n39161), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n39162));
    SB_LUT4 i1_3_lut_4_lut (.I0(tx_transmit_N_3513), .I1(n35184), .I2(\FRAME_MATCHER.i_31__N_2623 ), 
            .I3(n25063), .O(n169));   // verilog/coms.v(213[6] 220[9])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'he000;
    SB_LUT4 i1_2_lut_adj_911 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_911.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_912 (.I0(Kp_23__N_1426), .I1(\data_in_frame[11] [3]), 
            .I2(n44427), .I3(GND_net), .O(n44700));   // verilog/coms.v(72[16:41])
    defparam i2_3_lut_adj_912.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_913 (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[19] [5]), 
            .I2(\data_in_frame[19] [4]), .I3(GND_net), .O(n8_adj_4263));
    defparam i2_3_lut_adj_913.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_914 (.I0(\data_in_frame[19] [1]), .I1(n8_adj_4263), 
            .I2(n41670), .I3(\data_in_frame[19] [2]), .O(n10_adj_4264));
    defparam i4_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_915 (.I0(\data_in_frame[19] [7]), .I1(n10_adj_4264), 
            .I2(n46645), .I3(\data_in_frame[19] [6]), .O(n41549));
    defparam i5_4_lut_adj_915.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_916 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[18] [6]), 
            .I2(n42122), .I3(\data_in_frame[16] [4]), .O(n44521));   // verilog/coms.v(72[16:41])
    defparam i3_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[18] [7]), .I1(n44447), .I2(n6_adj_4265), 
            .I3(n42345), .O(n44424));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_917 (.I0(n28235), .I1(n44505), .I2(GND_net), 
            .I3(GND_net), .O(n44756));
    defparam i1_2_lut_adj_917.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_18_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n39160), .O(n2_adj_4266)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_adj_918 (.I0(n44703), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4267));
    defparam i2_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_919 (.I0(n44846), .I1(\data_in_frame[17] [6]), 
            .I2(n44427), .I3(\data_in_frame[15] [5]), .O(n14_adj_4268));
    defparam i6_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_920 (.I0(\data_in_frame[16] [0]), .I1(n14_adj_4268), 
            .I2(n10_adj_4267), .I3(n42356), .O(n46063));
    defparam i7_4_lut_adj_920.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_921 (.I0(\data_in_frame[18] [0]), .I1(n44818), 
            .I2(GND_net), .I3(GND_net), .O(n44846));
    defparam i1_2_lut_adj_921.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_922 (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[12] [2]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n44569));
    defparam i2_3_lut_adj_922.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44572));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_924 (.I0(\data_in_frame[16] [3]), .I1(n28941), 
            .I2(GND_net), .I3(GND_net), .O(n44530));
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_925 (.I0(n42368), .I1(n44530), .I2(\data_in_frame[16] [4]), 
            .I3(GND_net), .O(n42408));
    defparam i2_3_lut_adj_925.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_926 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[18] [1]), 
            .I2(\data_in_frame[10] [7]), .I3(GND_net), .O(n44780));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_926.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_927 (.I0(\data_in_frame[16] [7]), .I1(n44540), 
            .I2(n28264), .I3(\data_in_frame[16] [6]), .O(n44774));
    defparam i3_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_928 (.I0(n44774), .I1(\data_in_frame[17] [0]), 
            .I2(n42345), .I3(GND_net), .O(n46396));
    defparam i2_3_lut_adj_928.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_929 (.I0(\data_in_frame[12] [3]), .I1(n42341), 
            .I2(\data_in_frame[14] [4]), .I3(\data_in_frame[12] [2]), .O(n10_adj_4269));
    defparam i4_4_lut_adj_929.LUT_INIT = 16'h6996;
    SB_CARRY add_43_18 (.CI(n39160), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n39161));
    SB_LUT4 i5_3_lut_adj_930 (.I0(\data_in_frame[10] [0]), .I1(n10_adj_4269), 
            .I2(n27552), .I3(GND_net), .O(n42345));
    defparam i5_3_lut_adj_930.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_931 (.I0(n44569), .I1(n44671), .I2(\data_in_frame[10] [1]), 
            .I3(n28796), .O(n12_adj_4270));
    defparam i5_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_932 (.I0(n41819), .I1(n12_adj_4270), .I2(n44684), 
            .I3(n28160), .O(n42368));
    defparam i6_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_933 (.I0(n42368), .I1(\data_in_frame[16] [5]), 
            .I2(n42345), .I3(GND_net), .O(n44447));
    defparam i2_3_lut_adj_933.LUT_INIT = 16'h9696;
    SB_LUT4 i6_3_lut (.I0(\data_in_frame[18] [5]), .I1(n44410), .I2(\data_in_frame[18] [4]), 
            .I3(GND_net), .O(n38));
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i20_4_lut (.I0(n44252), .I1(\data_in_frame[18] [3]), .I2(\data_in_frame[12] [5]), 
            .I3(n46396), .O(n52));
    defparam i20_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i24_4_lut_adj_934 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[18] [2]), .I3(n42408), .O(n56));
    defparam i24_4_lut_adj_934.LUT_INIT = 16'h9669;
    SB_LUT4 i22_4_lut (.I0(n44544), .I1(n44447), .I2(n44524), .I3(n44364), 
            .O(n54));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n44279), .I1(n42341), .I2(\data_in_frame[10] [5]), 
            .I3(\data_in_frame[17] [6]), .O(n55));
    defparam i23_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i21_4_lut (.I0(n44849), .I1(n44637), .I2(n44792), .I3(n44572), 
            .O(n53));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_935 (.I0(n44780), .I1(n28749), .I2(n44486), 
            .I3(\data_in_frame[18] [7]), .O(n50_adj_4271));
    defparam i18_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(n44837), .I1(n52), .I2(n38), .I3(n44578), 
            .O(n58));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n53), .I1(n55), .I2(n54), .I3(n56), .O(n62));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_936 (.I0(\data_in_frame[17] [5]), .I1(n44569), 
            .I2(n44346), .I3(\data_in_frame[14] [1]), .O(n49));
    defparam i17_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_17_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n39159), .O(n2_adj_4272)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i31_4_lut (.I0(n49), .I1(n62), .I2(n58), .I3(n50_adj_4271), 
            .O(n42347));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_937 (.I0(n42122), .I1(n41670), .I2(\data_in_frame[13] [4]), 
            .I3(\data_in_frame[16] [0]), .O(n14_adj_4273));
    defparam i5_4_lut_adj_937.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_938 (.I0(n44852), .I1(n42347), .I2(n44530), .I3(n44846), 
            .O(n15_adj_4274));
    defparam i6_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_939 (.I0(n15_adj_4274), .I1(n44765), .I2(n14_adj_4273), 
            .I3(Kp_23__N_1536), .O(n46645));
    defparam i8_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_940 (.I0(n46645), .I1(n42347), .I2(GND_net), 
            .I3(GND_net), .O(n42343));
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_941 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44599));   // verilog/coms.v(70[16:62])
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_942 (.I0(n44611), .I1(n44205), .I2(n44393), 
            .I3(n41577), .O(n24_adj_4275));
    defparam i10_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_943 (.I0(n44664), .I1(n44224), .I2(n42413), .I3(\data_in_frame[14] [1]), 
            .O(n22));
    defparam i8_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_944 (.I0(n44599), .I1(n24_adj_4275), .I2(n18_adj_4276), 
            .I3(\data_in_frame[4] [3]), .O(n26_adj_4277));
    defparam i12_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[6] [7]), .I1(n26_adj_4277), .I2(n22), 
            .I3(\data_in_frame[11] [5]), .O(n28941));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_945 (.I0(n42356), .I1(n28941), .I2(\data_in_frame[16] [2]), 
            .I3(GND_net), .O(n44553));
    defparam i2_3_lut_adj_945.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_946 (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44765));
    defparam i1_2_lut_adj_946.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_947 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[9] [7]), .I3(n6_adj_4231), .O(n44410));
    defparam i4_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_948 (.I0(n28289), .I1(n44410), .I2(n28428), .I3(GND_net), 
            .O(n28235));
    defparam i2_3_lut_adj_948.LUT_INIT = 16'h9696;
    SB_CARRY add_43_17 (.CI(n39159), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n39160));
    SB_LUT4 i2_3_lut_adj_949 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[14] [5]), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n44505));
    defparam i2_3_lut_adj_949.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_950 (.I0(\data_in_frame[15] [0]), .I1(n44759), 
            .I2(n44505), .I3(\data_in_frame[17] [1]), .O(n44346));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_951 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44759));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_951.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_952 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[11] [2]), 
            .I2(n28719), .I3(n28655), .O(n44818));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_952.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_in_frame[18] [2]), .I1(n44818), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4278));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_954 (.I0(\data_in_frame[13] [7]), .I1(n28675), 
            .I2(n44777), .I3(n6_adj_4278), .O(n44233));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_954.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44810));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_956 (.I0(\data_in_frame[14] [2]), .I1(n44810), 
            .I2(\data_in_frame[9] [5]), .I3(\data_in_frame[11] [7]), .O(n44792));   // verilog/coms.v(70[16:62])
    defparam i3_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_in_frame[9] [3]), .I1(n41577), .I2(GND_net), 
            .I3(GND_net), .O(n44279));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_958 (.I0(n27601), .I1(n44684), .I2(n44393), .I3(n41622), 
            .O(n41819));
    defparam i3_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_959 (.I0(\data_in_frame[7] [3]), .I1(n29057), .I2(n8_adj_4279), 
            .I3(n44325), .O(n41577));
    defparam i1_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\data_in_frame[7] [1]), .I1(Kp_23__N_1228), 
            .I2(GND_net), .I3(GND_net), .O(n28630));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_961 (.I0(\data_in_frame[8] [5]), .I1(n44716), .I2(n41577), 
            .I3(n44587), .O(n20_adj_4280));
    defparam i8_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_962 (.I0(n44399), .I1(\data_in_frame[7] [0]), .I2(n28630), 
            .I3(n44658), .O(n19_adj_4281));
    defparam i7_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_963 (.I0(n44316), .I1(n28342), .I2(n28624), .I3(\data_in_frame[8] [7]), 
            .O(n21));
    defparam i9_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_964 (.I0(n21), .I1(n19_adj_4281), .I2(n20_adj_4280), 
            .I3(GND_net), .O(n27601));
    defparam i11_3_lut_adj_964.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1306));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(CLK_c), 
            .D(n43667), .S(n43543));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_965 (.I0(Kp_23__N_1306), .I1(\data_in_frame[9] [3]), 
            .I2(n44246), .I3(n6_adj_4260), .O(n44671));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_966 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44716));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_967 (.I0(n44671), .I1(n44367), .I2(n27552), .I3(GND_net), 
            .O(n41553));
    defparam i2_3_lut_adj_967.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_968 (.I0(n42082), .I1(\data_in_frame[8] [6]), .I2(n44444), 
            .I3(GND_net), .O(n14_adj_4282));
    defparam i5_3_lut_adj_968.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_969 (.I0(n44825), .I1(n41553), .I2(n44337), .I3(n44716), 
            .O(n15_adj_4283));
    defparam i6_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_970 (.I0(n15_adj_4283), .I1(n44413), .I2(n14_adj_4282), 
            .I3(n44208), .O(n42413));
    defparam i8_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_971 (.I0(n28171), .I1(n44349), .I2(\data_in_frame[11] [6]), 
            .I3(n42413), .O(n28_adj_4284));
    defparam i10_4_lut_adj_971.LUT_INIT = 16'h9669;
    SB_LUT4 i14_3_lut (.I0(n28618), .I1(n28_adj_4284), .I2(n44524), .I3(GND_net), 
            .O(n32));
    defparam i14_3_lut.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(CLK_c), 
            .D(n43665), .S(n43547));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(CLK_c), 
            .D(n43663), .S(n43551));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(CLK_c), 
            .D(n43661), .S(n43555));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(CLK_c), 
            .D(n7_adj_4285), .S(n8_adj_4286));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(CLK_c), 
            .D(n43659), .S(n43559));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(CLK_c), 
            .D(n7_adj_4287), .S(n8_adj_4288));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(CLK_c), 
            .D(n43657), .S(n43563));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(CLK_c), 
            .D(n43655), .S(n43567));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(CLK_c), 
            .D(n43653), .S(n43571));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(CLK_c), 
            .D(n35190), .S(n36044));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(CLK_c), 
            .D(n43651), .S(n43575));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(CLK_c), 
            .D(n43649), .S(n43579));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(CLK_c), 
            .D(n43647), .S(n43583));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(CLK_c), 
            .D(n7_adj_4289), .S(n8_adj_4290));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(CLK_c), 
            .D(n43645), .S(n43587));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(CLK_c), 
            .D(n43643), .S(n43591));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(CLK_c), 
            .D(n43641), .S(n43595));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(CLK_c), 
            .D(n43639), .S(n43513));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_972 (.I0(n41819), .I1(n44236), .I2(n44611), 
            .I3(\data_in_frame[4] [7]), .O(n30));
    defparam i12_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_973 (.I0(\data_in_frame[12] [1]), .I1(n29060), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[5] [0]), .O(n31_adj_4291));
    defparam i13_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_974 (.I0(n44792), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[0] [2]), .I3(\data_in_frame[4] [6]), .O(n29));
    defparam i11_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_975 (.I0(n29), .I1(n31_adj_4291), .I2(n30), 
            .I3(n32), .O(n42122));
    defparam i17_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_976 (.I0(\data_in_frame[5] [2]), .I1(n28890), .I2(\data_in_frame[7] [4]), 
            .I3(n28494), .O(n44349));
    defparam i3_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_977 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44246));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_977.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_978 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4292));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_978.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_979 (.I0(n28342), .I1(n28749), .I2(n44246), .I3(n6_adj_4292), 
            .O(n44852));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_979.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(CLK_c), 
            .D(n43637), .S(n43505));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(CLK_c), 
            .D(n43635), .S(n43493));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1536));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_980 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [3]), 
            .I2(n42122), .I3(GND_net), .O(n44544));
    defparam i2_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_981 (.I0(n44544), .I1(n44777), .I2(Kp_23__N_1536), 
            .I3(GND_net), .O(n42398));
    defparam i2_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_982 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44224));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_983 (.I0(\data_in_frame[15] [4]), .I1(n28655), 
            .I2(\data_in_frame[13] [3]), .I3(GND_net), .O(n44849));
    defparam i2_3_lut_adj_983.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(CLK_c), 
            .D(n43633), .S(n43599));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(CLK_c), 
            .D(n43631), .S(n43509));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(CLK_c), 
            .D(n43629), .S(n43603));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(CLK_c), 
            .D(n43627), .S(n43607));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(CLK_c), 
            .D(n43625), .S(n43611));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(CLK_c), 
            .D(n43623), .S(n43489));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n43485), .S(n43691));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_984 (.I0(n44849), .I1(n28319), .I2(\data_in_frame[11] [2]), 
            .I3(\data_in_frame[11] [0]), .O(n44547));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_984.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4293));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_986 (.I0(n44547), .I1(\data_in_frame[13] [1]), 
            .I2(n44813), .I3(n6_adj_4293), .O(n41670));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_987 (.I0(\data_in_frame[14] [7]), .I1(n28264), 
            .I2(GND_net), .I3(GND_net), .O(n28705));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_988 (.I0(n44453), .I1(\data_in_frame[6] [7]), .I2(\data_in_frame[2] [6]), 
            .I3(n44652), .O(n10_adj_4294));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_989 (.I0(\data_in_frame[4] [7]), .I1(n10_adj_4294), 
            .I2(\data_in_frame[4] [5]), .I3(GND_net), .O(Kp_23__N_1228));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_adj_989.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_990 (.I0(Kp_23__N_1228), .I1(n28618), .I2(n28837), 
            .I3(GND_net), .O(Kp_23__N_1426));   // verilog/coms.v(72[16:41])
    defparam i2_3_lut_adj_990.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_16_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n39158), .O(n2_adj_4295)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_991 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n44364));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_991.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_0__5__I_0_2_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_981));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_0__5__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_992 (.I0(\data_in_frame[5] [0]), .I1(n29057), .I2(\data_in_frame[7] [2]), 
            .I3(n28840), .O(n44205));
    defparam i3_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_993 (.I0(n29017), .I1(n44205), .I2(n28445), .I3(\data_in_frame[4] [6]), 
            .O(n28749));
    defparam i3_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n29310), .D(n46112));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_994 (.I0(n44713), .I1(\data_in_frame[2] [4]), .I2(\data_in_frame[0] [0]), 
            .I3(n44789), .O(n10_adj_4258));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_995 (.I0(Kp_23__N_1217), .I1(n28749), .I2(GND_net), 
            .I3(GND_net), .O(n28624));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_996 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28171));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_996.LUT_INIT = 16'h6666;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n29310), .D(n45837));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n29310), .D(n45838));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n29310), .D(n45552));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n29310), .D(n45583));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n29310), .D(n44577));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(CLK_c), 
            .E(n29310), .D(n28794));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n29310), .D(n45554));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n29310), .D(n46786));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n29310), .D(n45780));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n29310), .D(n46761));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n29310), .D(n46120));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n29310), .D(n45896));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n29310), .D(n46218));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n29310), .D(n46058));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_997 (.I0(n44364), .I1(n44431), .I2(Kp_23__N_1426), 
            .I3(GND_net), .O(n28675));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_997.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_998 (.I0(\data_in_frame[8] [6]), .I1(n44227), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[4] [4]), .O(n10_adj_4296));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_999 (.I0(\data_in_frame[4] [3]), .I1(n10_adj_4296), 
            .I2(n4_c), .I3(GND_net), .O(n44399));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_999.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_0__1__I_0_2_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_977));   // verilog/coms.v(72[16:27])
    defparam data_in_frame_0__1__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1000 (.I0(Kp_23__N_993), .I1(n44664), .I2(n44402), 
            .I3(Kp_23__N_977), .O(Kp_23__N_1096));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1001 (.I0(\data_in_frame[8] [5]), .I1(n44396), 
            .I2(Kp_23__N_1096), .I3(\data_in_frame[6] [4]), .O(n28736));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1001.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1002 (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44713));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1003 (.I0(\data_in_frame[2] [1]), .I1(n44713), 
            .I2(\data_in_frame[4] [3]), .I3(\data_in_frame[4] [5]), .O(n44236));
    defparam i3_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4297));
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1005 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [4]), 
            .I2(n44236), .I3(n6_adj_4297), .O(n44658));
    defparam i4_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44337));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in_frame[5] [3]), .I1(n44384), 
            .I2(GND_net), .I3(GND_net), .O(n28494));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1008 (.I0(\data_in_frame[1] [3]), .I1(n28843), 
            .I2(n28494), .I3(n28114), .O(n10_adj_4298));
    defparam i4_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1009 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[3] [1]), 
            .I2(n10_adj_4298), .I3(\data_in_frame[5] [4]), .O(n28428));
    defparam i1_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1010 (.I0(n44367), .I1(n28428), .I2(n28837), 
            .I3(GND_net), .O(n44837));
    defparam i3_3_lut_adj_1010.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n51372), .I2(n49725), .I3(byte_transmit_counter[4]), .O(n51567));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51567_bdd_4_lut (.I0(n51567), .I1(n51468), .I2(n7_adj_4299), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n51567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36092 (.I0(byte_transmit_counter[3]), 
            .I1(n51378), .I2(n49722), .I3(byte_transmit_counter[4]), .O(n51561));
    defparam byte_transmit_counter_3__bdd_4_lut_36092.LUT_INIT = 16'he4aa;
    SB_LUT4 n51561_bdd_4_lut (.I0(n51561), .I1(n51462), .I2(n7_adj_4300), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n51561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36087 (.I0(byte_transmit_counter[3]), 
            .I1(n51384), .I2(n49719), .I3(byte_transmit_counter[4]), .O(n51555));
    defparam byte_transmit_counter_3__bdd_4_lut_36087.LUT_INIT = 16'he4aa;
    SB_LUT4 n51555_bdd_4_lut (.I0(n51555), .I1(n51456), .I2(n7_adj_4301), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n51555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36082 (.I0(byte_transmit_counter[3]), 
            .I1(n51390), .I2(n49713), .I3(byte_transmit_counter[4]), .O(n51549));
    defparam byte_transmit_counter_3__bdd_4_lut_36082.LUT_INIT = 16'he4aa;
    SB_LUT4 n51549_bdd_4_lut (.I0(n51549), .I1(n51450), .I2(n7_adj_4302), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n51549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36077 (.I0(byte_transmit_counter[3]), 
            .I1(n51396), .I2(n49710), .I3(byte_transmit_counter[4]), .O(n51543));
    defparam byte_transmit_counter_3__bdd_4_lut_36077.LUT_INIT = 16'he4aa;
    SB_LUT4 n51543_bdd_4_lut (.I0(n51543), .I1(n51444), .I2(n7_adj_4303), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n51543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36072 (.I0(byte_transmit_counter[3]), 
            .I1(n51402), .I2(n49707), .I3(byte_transmit_counter[4]), .O(n51537));
    defparam byte_transmit_counter_3__bdd_4_lut_36072.LUT_INIT = 16'he4aa;
    SB_LUT4 n51537_bdd_4_lut (.I0(n51537), .I1(n51438), .I2(n7_adj_4304), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n51537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36067 (.I0(byte_transmit_counter[3]), 
            .I1(n51408), .I2(n49704), .I3(byte_transmit_counter[4]), .O(n51531));
    defparam byte_transmit_counter_3__bdd_4_lut_36067.LUT_INIT = 16'he4aa;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_4305), .S(n3_adj_4306));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4307), .S(n3_adj_4308));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4309), .S(n3_adj_4310));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4311), .S(n3_adj_4312));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_4211), .S(n3_adj_4313));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_4212), .S(n3_adj_4314));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_4214), .S(n3_adj_4315));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_4243), .S(n3_adj_4316));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_4246), .S(n3_adj_4317));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_4250), .S(n3_adj_4318));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_4252), .S(n3_adj_4319));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_4257), .S(n3_adj_4320));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_4259), .S(n3_adj_4321));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_4261), .S(n3_adj_4322));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_4262), .S(n3_adj_4323));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_4266), .S(n3_adj_4324));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_4272), .S(n3_adj_4325));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_4295), .S(n3_adj_4326));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_4327), .S(n3_adj_4328));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_4329), .S(n3_adj_4330));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_4331), .S(n3_adj_4332));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_4333), .S(n3_adj_4334));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_4335), .S(n3_adj_4336));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_4337), .S(n3_adj_4338));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4339), .S(n3_adj_4340));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4341), .S(n3_adj_4342));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4343), .S(n3_adj_4344));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4345), .S(n3_adj_4346));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_4347), .S(n3_adj_4348));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4349), .S(n3_adj_4350));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4351), .S(n3_adj_4352));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1011 (.I0(n28719), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[11] [0]), .I3(GND_net), .O(n44690));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1012 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[13] [2]), 
            .I2(n44813), .I3(n44239), .O(n44306));
    defparam i3_4_lut_adj_1012.LUT_INIT = 16'h6996;
    SB_CARRY add_43_16 (.CI(n39158), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n39159));
    SB_LUT4 add_43_15_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n39157), .O(n2_adj_4327)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28114));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(n28238), .I1(n44834), .I2(GND_net), 
            .I3(GND_net), .O(n44199));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1015 (.I0(\data_in_frame[1] [4]), .I1(n44741), 
            .I2(n44495), .I3(\data_in_frame[1] [2]), .O(n46131));
    defparam i3_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1016 (.I0(n28615), .I1(n28156), .I2(\data_in_frame[1] [1]), 
            .I3(n44413), .O(n10_adj_4353));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_CARRY add_43_15 (.CI(n39157), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n39158));
    SB_LUT4 i1_2_lut_adj_1017 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n28612));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1018 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1018.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_0__7__I_0_3901_2_lut (.I0(\data_in_frame[0] [7]), 
            .I1(\data_in_frame[0] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_974));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_0__7__I_0_3901_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1019 (.I0(\data_in_frame[0] [0]), .I1(n44602), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n28204));   // verilog/coms.v(70[16:62])
    defparam i2_3_lut_adj_1019.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_14_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n39156), .O(n2_adj_4329)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44664));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(\data_in_frame[2] [6]), .I1(n44384), 
            .I2(GND_net), .I3(GND_net), .O(n44352));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1022 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[5] [2]), .I3(GND_net), .O(n44325));
    defparam i2_3_lut_adj_1022.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1023 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[1] [0]), .O(n28890));
    defparam i3_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_CARRY add_43_14 (.CI(n39156), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n39157));
    SB_LUT4 add_43_13_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n39155), .O(n2_adj_4331)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1024 (.I0(\data_in_frame[5] [4]), .I1(n28890), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n44834));
    defparam i2_3_lut_adj_1024.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28156));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44402));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44789));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4221), 
            .I2(n63_adj_4224), .I3(n63), .O(\FRAME_MATCHER.state_31__N_2660[2] ));   // verilog/coms.v(112[11:16])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hb300;
    SB_LUT4 i4_2_lut_adj_1028 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4354));   // verilog/coms.v(78[16:27])
    defparam i4_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut_adj_1029 (.I0(n44789), .I1(n44402), .I2(n44495), 
            .I3(n44293), .O(n36));   // verilog/coms.v(78[16:27])
    defparam i14_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1030 (.I0(n44834), .I1(n44453), .I2(n44256), 
            .I3(\data_in_frame[3] [3]), .O(n34));   // verilog/coms.v(78[16:27])
    defparam i12_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1031 (.I0(n44605), .I1(n36), .I2(n26_adj_4354), 
            .I3(n44325), .O(n40_adj_4355));   // verilog/coms.v(78[16:27])
    defparam i18_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1032 (.I0(n44352), .I1(n44664), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[2] [4]), .O(n38_adj_4356));   // verilog/coms.v(78[16:27])
    defparam i16_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i17_3_lut (.I0(\data_in_frame[2] [5]), .I1(n34), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(n39_adj_4357));   // verilog/coms.v(78[16:27])
    defparam i17_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut_adj_1033 (.I0(n28204), .I1(\data_in_frame[5] [3]), 
            .I2(n29060), .I3(\data_in_frame[2] [3]), .O(n37));   // verilog/coms.v(78[16:27])
    defparam i15_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1034 (.I0(n37), .I1(n39_adj_4357), .I2(n38_adj_4356), 
            .I3(n40_adj_4355), .O(n42082));   // verilog/coms.v(78[16:27])
    defparam i21_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\data_in_frame[6] [0]), .I1(n44831), 
            .I2(GND_net), .I3(GND_net), .O(n44208));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(n4_c), .I1(n29017), .I2(GND_net), .I3(GND_net), 
            .O(Kp_23__N_1020));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(\data_in_frame[4] [5]), .I1(n42082), 
            .I2(GND_net), .I3(GND_net), .O(n44786));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44482));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1039 (.I0(n44786), .I1(Kp_23__N_1020), .I2(n44208), 
            .I3(n44596), .O(n44741));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1040 (.I0(\data_in_frame[3] [3]), .I1(n44825), 
            .I2(n44741), .I3(n44482), .O(n42452));
    defparam i3_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4358));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h6666;
    SB_CARRY add_43_13 (.CI(n39155), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n39156));
    SB_LUT4 i4_4_lut_adj_1042 (.I0(n28796), .I1(n46131), .I2(n44199), 
            .I3(n6_adj_4358), .O(n44587));
    defparam i4_4_lut_adj_1042.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_12_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n39154), .O(n2_adj_4333)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n51531_bdd_4_lut (.I0(n51531), .I1(n51432), .I2(n7_adj_4359), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n51531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n51525));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51525_bdd_4_lut (.I0(n51525), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n51528));
    defparam n51525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36057 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27][1] ), 
            .I3(byte_transmit_counter[1]), .O(n51519));
    defparam byte_transmit_counter_0__bdd_4_lut_36057.LUT_INIT = 16'he4aa;
    SB_LUT4 n51519_bdd_4_lut (.I0(n51519), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n51522));
    defparam n51519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36052 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n51513));
    defparam byte_transmit_counter_0__bdd_4_lut_36052.LUT_INIT = 16'he4aa;
    SB_LUT4 n51513_bdd_4_lut (.I0(n51513), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n51516));
    defparam n51513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36047 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n51507));
    defparam byte_transmit_counter_0__bdd_4_lut_36047.LUT_INIT = 16'he4aa;
    SB_LUT4 n51507_bdd_4_lut (.I0(n51507), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n51510));
    defparam n51507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36042 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n51501));
    defparam byte_transmit_counter_0__bdd_4_lut_36042.LUT_INIT = 16'he4aa;
    SB_LUT4 n51501_bdd_4_lut (.I0(n51501), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n51504));
    defparam n51501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36037 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n51495));
    defparam byte_transmit_counter_0__bdd_4_lut_36037.LUT_INIT = 16'he4aa;
    SB_LUT4 n51495_bdd_4_lut (.I0(n51495), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n51498));
    defparam n51495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36032 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n51489));
    defparam byte_transmit_counter_0__bdd_4_lut_36032.LUT_INIT = 16'he4aa;
    SB_LUT4 n51489_bdd_4_lut (.I0(n51489), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n51492));
    defparam n51489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36027 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n51483));
    defparam byte_transmit_counter_0__bdd_4_lut_36027.LUT_INIT = 16'he4aa;
    SB_LUT4 n51483_bdd_4_lut (.I0(n51483), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n51486));
    defparam n51483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36062 (.I0(byte_transmit_counter[3]), 
            .I1(n51366), .I2(n49728), .I3(byte_transmit_counter[4]), .O(n51477));
    defparam byte_transmit_counter_3__bdd_4_lut_36062.LUT_INIT = 16'he4aa;
    SB_LUT4 n51477_bdd_4_lut (.I0(n51477), .I1(n51426), .I2(n7_adj_4360), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n51477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_adj_1043 (.I0(n44622), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4361));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_adj_1043.LUT_INIT = 16'h6666;
    SB_CARRY add_43_12 (.CI(n39154), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n39155));
    SB_LUT4 i6_4_lut_adj_1044 (.I0(n44744), .I1(\data_in_frame[1] [2]), 
            .I2(n44608), .I3(\data_in_frame[4] [0]), .O(n14_adj_4362));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1045 (.I0(\data_in_frame[10] [3]), .I1(n14_adj_4362), 
            .I2(n10_adj_4361), .I3(n44444), .O(n28753));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1046 (.I0(\data_in_frame[10] [2]), .I1(n44587), 
            .I2(n42452), .I3(\data_in_frame[7] [7]), .O(n42341));
    defparam i3_4_lut_adj_1046.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_11_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n39153), .O(n2_adj_4335)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1047 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n44239));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1047.LUT_INIT = 16'h9696;
    SB_CARRY add_43_11 (.CI(n39153), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n39154));
    SB_LUT4 i5_4_lut_adj_1048 (.I0(n44306), .I1(\data_in_frame[13] [0]), 
            .I2(n44690), .I3(n44416), .O(n12_adj_4363));   // verilog/coms.v(76[16:43])
    defparam i5_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1049 (.I0(n44239), .I1(n12_adj_4363), .I2(\data_in_frame[17] [4]), 
            .I3(n44355), .O(n41565));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1050 (.I0(n42341), .I1(n28753), .I2(\data_in_frame[12] [4]), 
            .I3(GND_net), .O(n46102));
    defparam i2_3_lut_adj_1050.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1051 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44227));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1051.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_10_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n39152), .O(n2_adj_4337)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1052 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28615));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1052.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44608));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1054 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n28238));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1054.LUT_INIT = 16'h9696;
    SB_CARRY add_43_10 (.CI(n39152), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n39153));
    SB_LUT4 i3_4_lut_adj_1055 (.I0(n28238), .I1(n44608), .I2(n44218), 
            .I3(n28615), .O(n28160));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\data_in_frame[8] [2]), .I1(n28160), 
            .I2(GND_net), .I3(GND_net), .O(n44316));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_993));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1057 (.I0(n44227), .I1(\data_in_frame[4] [2]), 
            .I2(n44611), .I3(n6_adj_4364), .O(n44396));   // verilog/coms.v(70[16:69])
    defparam i4_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44355));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_9_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n39151), .O(n2_adj_4339)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1059 (.I0(n44296), .I1(n44396), .I2(\data_in_frame[8] [4]), 
            .I3(GND_net), .O(n28319));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1059.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44584));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44218));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44605));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1063 (.I0(\data_in_frame[4] [0]), .I1(n44605), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[1] [6]), .O(n12_adj_4365));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1064 (.I0(\data_in_frame[1] [7]), .I1(n12_adj_4365), 
            .I2(\data_in_frame[6] [2]), .I3(n44218), .O(n44296));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_CARRY add_43_9 (.CI(n39151), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n39152));
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_in_frame[8] [3]), .I1(n44296), 
            .I2(GND_net), .I3(GND_net), .O(n44637));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1066 (.I0(\data_in_frame[1] [4]), .I1(n44622), 
            .I2(n44256), .I3(\data_in_frame[3] [5]), .O(n28289));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_8_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n39150), .O(n2_adj_4341)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1067 (.I0(\data_in_frame[15] [0]), .I1(n28313), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4366));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1067.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1068 (.I0(n28349), .I1(n28319), .I2(n44355), 
            .I3(n6_adj_4366), .O(n28716));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\data_in_frame[10] [5]), .I1(n44343), 
            .I2(GND_net), .I3(GND_net), .O(n28956));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1070 (.I0(n28956), .I1(\data_in_frame[14] [7]), 
            .I2(n28716), .I3(\data_in_frame[13] [0]), .O(n10_adj_4367));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1071 (.I0(n44252), .I1(n10_adj_4367), .I2(\data_in_frame[10] [6]), 
            .I3(GND_net), .O(n44771));   // verilog/coms.v(76[16:43])
    defparam i5_3_lut_adj_1071.LUT_INIT = 16'h9696;
    SB_LUT4 i34508_2_lut (.I0(n51486), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49704));
    defparam i34508_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1072 (.I0(\data_in_frame[17] [2]), .I1(n46102), 
            .I2(n41565), .I3(GND_net), .O(n44486));
    defparam i2_3_lut_adj_1072.LUT_INIT = 16'h6969;
    SB_LUT4 i33380_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n48817));
    defparam i33380_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i1_2_lut_3_lut_adj_1073 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n43611));
    defparam i1_2_lut_3_lut_adj_1073.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1074 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4368));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_1074.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1075 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4369));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_1075.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1076 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_1076.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_2_lut_3_lut_adj_1077 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n43607));
    defparam i1_2_lut_3_lut_adj_1077.LUT_INIT = 16'he0e0;
    SB_LUT4 i33378_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48815));
    defparam i33378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1078 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n43603));
    defparam i1_2_lut_3_lut_adj_1078.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_4_lut_adj_1079 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_4370));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_1079.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1080 (.I0(n9_adj_4370), .I1(n11), .I2(n10_adj_4369), 
            .I3(n12_adj_4368), .O(n25324));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1080.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1081 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n43599));
    defparam i1_2_lut_3_lut_adj_1081.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_3_lut_adj_1082 (.I0(\data_in_frame[14] [6]), .I1(n44486), 
            .I2(n44771), .I3(GND_net), .O(n8_adj_4371));
    defparam i3_3_lut_adj_1082.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1083 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[19] [5]), 
            .I2(n44661), .I3(n44343), .O(n16_adj_4372));
    defparam i6_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i34485_2_lut (.I0(n51492), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49707));
    defparam i34485_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i8_3_lut_adj_1084 (.I0(\data_in_frame[21] [7]), .I1(n16_adj_4372), 
            .I2(n41670), .I3(GND_net), .O(n18_adj_4373));
    defparam i8_3_lut_adj_1084.LUT_INIT = 16'h9696;
    SB_LUT4 i33370_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48807));
    defparam i33370_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33371_4_lut (.I0(n48807), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48808));
    defparam i33371_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i33369_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48806));
    defparam i33369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1085 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n43595));
    defparam i1_2_lut_3_lut_adj_1085.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1086 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n43591));
    defparam i1_2_lut_3_lut_adj_1086.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1087 (.I0(\data_in_frame[18] [5]), .I1(n42398), 
            .I2(\data_in_frame[18] [4]), .I3(GND_net), .O(n6_adj_4374));
    defparam i2_3_lut_adj_1087.LUT_INIT = 16'h9696;
    SB_LUT4 i34482_2_lut (.I0(n51498), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49710));
    defparam i34482_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i9_4_lut_adj_1088 (.I0(\data_in_frame[19] [6]), .I1(n18_adj_4373), 
            .I2(n14_adj_4375), .I3(n44759), .O(n46262));
    defparam i9_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i33364_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48801));
    defparam i33364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33365_4_lut (.I0(n48801), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48802));
    defparam i33365_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i33363_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48800));
    defparam i33363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1089 (.I0(n44233), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[16] [0]), .I3(GND_net), .O(n6_adj_4376));
    defparam i1_3_lut_adj_1089.LUT_INIT = 16'h9696;
    SB_LUT4 i34479_2_lut (.I0(n51504), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49713));
    defparam i34479_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i6_4_lut_adj_1090 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[19] [3]), 
            .I2(n44346), .I3(n28319), .O(n16_adj_4377));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1091 (.I0(\data_in_frame[19] [4]), .I1(n28235), 
            .I2(n44661), .I3(n28956), .O(n17_adj_4378));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1092 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[20] [5]), 
            .I2(n42380), .I3(GND_net), .O(n8_adj_4379));
    defparam i3_3_lut_adj_1092.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1093 (.I0(n17_adj_4378), .I1(\data_in_frame[21] [5]), 
            .I2(n16_adj_4377), .I3(\data_in_frame[16] [7]), .O(n46883));   // verilog/coms.v(75[16:43])
    defparam i9_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1094 (.I0(\data_in_frame[17] [5]), .I1(n41565), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4380));   // verilog/coms.v(85[17:28])
    defparam i4_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_CARRY add_43_8 (.CI(n39150), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n39151));
    SB_LUT4 i7_4_lut_adj_1095 (.I0(n13_adj_4380), .I1(n46063), .I2(\data_in_frame[20] [0]), 
            .I3(n42380), .O(n16_adj_4381));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i33358_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48795));
    defparam i33358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33359_4_lut (.I0(n48795), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n48796));
    defparam i33359_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i1_2_lut_3_lut_adj_1096 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n43587));
    defparam i1_2_lut_3_lut_adj_1096.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_4_lut_adj_1097 (.I0(n44233), .I1(n44572), .I2(\data_in_frame[20] [3]), 
            .I3(n42356), .O(n12_adj_4382));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_1097.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1098 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[19] [2]), .I3(GND_net), .O(n10_adj_4383));
    defparam i2_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1099 (.I0(n44756), .I1(n28716), .I2(n44424), 
            .I3(\data_in_frame[17] [1]), .O(n14_adj_4384));
    defparam i6_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1100 (.I0(\data_in_frame[21] [3]), .I1(n14_adj_4384), 
            .I2(n10_adj_4383), .I3(n28705), .O(n46244));
    defparam i7_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1101 (.I0(n44521), .I1(\data_in_frame[21] [2]), 
            .I2(\data_in_frame[19] [1]), .I3(n44774), .O(n10_adj_4385));
    defparam i4_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1102 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n43583));
    defparam i1_2_lut_3_lut_adj_1102.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1103 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[18] [5]), 
            .I2(n41549), .I3(GND_net), .O(n6_adj_4386));
    defparam i2_3_lut_adj_1103.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1104 (.I0(\data_in_frame[19] [0]), .I1(n10_adj_4385), 
            .I2(\data_in_frame[17] [0]), .I3(GND_net), .O(n46339));
    defparam i5_3_lut_adj_1104.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1105 (.I0(\data_in_frame[13] [4]), .I1(n44572), 
            .I2(n8_adj_4232), .I3(n44700), .O(n12_adj_4387));
    defparam i4_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1106 (.I0(\data_in_frame[20] [1]), .I1(n42398), 
            .I2(n42356), .I3(n42380), .O(n13_adj_4388));
    defparam i5_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1107 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n43579));
    defparam i1_2_lut_3_lut_adj_1107.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_4_lut_adj_1108 (.I0(\data_in_frame[19] [2]), .I1(n44540), 
            .I2(\data_in_frame[21] [4]), .I3(\data_in_frame[17] [2]), .O(n12_adj_4389));
    defparam i5_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i33357_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48794));
    defparam i33357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1109 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n43575));
    defparam i1_2_lut_3_lut_adj_1109.LUT_INIT = 16'he0e0;
    SB_LUT4 i34476_2_lut (.I0(n51510), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49719));
    defparam i34476_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1110 (.I0(\data_in_frame[21] [6]), .I1(n8_adj_4371), 
            .I2(\data_in_frame[19] [5]), .I3(\data_in_frame[19] [4]), .O(n46324));
    defparam i4_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i33216_4_lut (.I0(\data_in_frame[20] [6]), .I1(n46262), .I2(n6_adj_4374), 
            .I3(n42408), .O(n48581));
    defparam i33216_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i1_2_lut_3_lut_adj_1111 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n43571));
    defparam i1_2_lut_3_lut_adj_1111.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1112 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n43567));
    defparam i1_2_lut_3_lut_adj_1112.LUT_INIT = 16'he0e0;
    SB_LUT4 i33352_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48789));
    defparam i33352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33353_4_lut (.I0(n48789), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n48790));
    defparam i33353_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i33351_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48788));
    defparam i33351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_3_lut (.I0(n46396), .I1(n44771), .I2(\data_in_frame[19] [3]), 
            .I3(GND_net), .O(n11_adj_4390));
    defparam i4_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i34473_2_lut (.I0(n51516), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49722));
    defparam i34473_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1113 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[20] [4]), 
            .I2(n44553), .I3(n6_adj_4376), .O(n46425));
    defparam i4_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1114 (.I0(n46883), .I1(\data_in_frame[18] [4]), 
            .I2(n8_adj_4379), .I3(n42398), .O(n22_adj_4391));
    defparam i6_4_lut_adj_1114.LUT_INIT = 16'hebbe;
    SB_LUT4 i12_4_lut_adj_1115 (.I0(n11_adj_4390), .I1(n48581), .I2(n46324), 
            .I3(n12_adj_4389), .O(n28_adj_4392));
    defparam i12_4_lut_adj_1115.LUT_INIT = 16'hf7fb;
    SB_LUT4 i1_2_lut_3_lut_adj_1116 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n43563));
    defparam i1_2_lut_3_lut_adj_1116.LUT_INIT = 16'he0e0;
    SB_LUT4 i7_4_lut_adj_1117 (.I0(n13_adj_4388), .I1(\data_in_frame[19] [7]), 
            .I2(n12_adj_4387), .I3(n42343), .O(n46724));
    defparam i7_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1118 (.I0(n44521), .I1(\data_in_frame[21] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4393));
    defparam i2_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i33347_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n48784));
    defparam i33347_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i8_4_lut_adj_1119 (.I0(n44306), .I1(n16_adj_4381), .I2(n12_adj_4394), 
            .I3(n42398), .O(n45599));   // verilog/coms.v(85[17:28])
    defparam i8_4_lut_adj_1119.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1120 (.I0(n46063), .I1(\data_in_frame[20] [2]), 
            .I2(n44547), .I3(n6_adj_4395), .O(n46374));
    defparam i4_4_lut_adj_1120.LUT_INIT = 16'h9669;
    SB_LUT4 i33345_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48782));
    defparam i33345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_7_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n39149), .O(n2_adj_4343)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1121 (.I0(\data_in_frame[18] [1]), .I1(n12_adj_4382), 
            .I2(n44700), .I3(\data_in_frame[16] [1]), .O(n45835));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i34469_2_lut (.I0(n51522), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49725));
    defparam i34469_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_4_lut_adj_1122 (.I0(\data_in_frame[19] [0]), .I1(n6_adj_4393), 
            .I2(n42345), .I3(n41549), .O(n46136));
    defparam i3_4_lut_adj_1122.LUT_INIT = 16'h9669;
    SB_LUT4 i33218_4_lut (.I0(n46244), .I1(n41549), .I2(n44424), .I3(\data_in_frame[21] [1]), 
            .O(n48583));
    defparam i33218_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i33220_4_lut (.I0(\data_in_frame[20] [7]), .I1(n46339), .I2(n6_adj_4386), 
            .I3(n42408), .O(n48585));
    defparam i33220_4_lut.LUT_INIT = 16'h4884;
    SB_CARRY add_43_7 (.CI(n39149), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n39150));
    SB_LUT4 i14_4_lut_adj_1123 (.I0(n46724), .I1(n28_adj_4392), .I2(n22_adj_4391), 
            .I3(n46425), .O(n30_adj_4396));
    defparam i14_4_lut_adj_1123.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_1124 (.I0(n46136), .I1(n45835), .I2(n46374), 
            .I3(n45599), .O(n25_adj_4397));
    defparam i9_4_lut_adj_1124.LUT_INIT = 16'hfffb;
    SB_LUT4 i15_4_lut_adj_1125 (.I0(n25_adj_4397), .I1(n30_adj_4396), .I2(n48585), 
            .I3(n48583), .O(n31_adj_4230));
    defparam i15_4_lut_adj_1125.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1126 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n43559));
    defparam i1_2_lut_3_lut_adj_1126.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1127 (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4221), 
            .I2(n63_adj_4224), .I3(n20372), .O(n4));   // verilog/coms.v(112[11:16])
    defparam i1_2_lut_4_lut_adj_1127.LUT_INIT = 16'hb300;
    SB_LUT4 add_43_6_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n39148), .O(n2_adj_4345)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1128 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n43555));
    defparam i1_2_lut_3_lut_adj_1128.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_6 (.CI(n39148), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n39149));
    SB_LUT4 i1_2_lut_3_lut_adj_1129 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n43551));
    defparam i1_2_lut_3_lut_adj_1129.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1130 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n43547));
    defparam i1_2_lut_3_lut_adj_1130.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1131 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n43543));
    defparam i1_2_lut_3_lut_adj_1131.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1132 (.I0(n190), .I1(n44183), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n43539));
    defparam i1_2_lut_3_lut_adj_1132.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1133 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n43623));
    defparam i1_2_lut_3_lut_adj_1133.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1134 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n43625));
    defparam i1_2_lut_3_lut_adj_1134.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1135 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n43627));
    defparam i1_2_lut_3_lut_adj_1135.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1136 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n43629));
    defparam i1_2_lut_3_lut_adj_1136.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1137 (.I0(\FRAME_MATCHER.state [1]), .I1(n44134), 
            .I2(n31_adj_4230), .I3(n25324), .O(n29176));
    defparam i3_4_lut_adj_1137.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_3_lut_adj_1138 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n43631));
    defparam i1_2_lut_3_lut_adj_1138.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_5_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n39147), .O(n2_adj_4347)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_5 (.CI(n39147), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n39148));
    SB_LUT4 add_43_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n39146), .O(n2_adj_4349)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_4 (.CI(n39146), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n39147));
    SB_LUT4 add_43_3_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n39145), .O(n2_adj_4351)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_3 (.CI(n39145), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n39146));
    SB_LUT4 add_43_2_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n48719), .I2(n48720), .I3(byte_transmit_counter[2]), .O(n51465));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51465_bdd_4_lut (.I0(n51465), .I1(n48873), .I2(n48872), .I3(byte_transmit_counter[2]), 
            .O(n51468));
    defparam n51465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36010 (.I0(byte_transmit_counter[1]), 
            .I1(n48722), .I2(n48723), .I3(byte_transmit_counter[2]), .O(n51459));
    defparam byte_transmit_counter_1__bdd_4_lut_36010.LUT_INIT = 16'he4aa;
    SB_LUT4 n51459_bdd_4_lut (.I0(n51459), .I1(n48870), .I2(n48869), .I3(byte_transmit_counter[2]), 
            .O(n51462));
    defparam n51459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36005 (.I0(byte_transmit_counter[1]), 
            .I1(n48863), .I2(n48864), .I3(byte_transmit_counter[2]), .O(n51453));
    defparam byte_transmit_counter_1__bdd_4_lut_36005.LUT_INIT = 16'he4aa;
    SB_LUT4 n51453_bdd_4_lut (.I0(n51453), .I1(n48858), .I2(n48857), .I3(byte_transmit_counter[2]), 
            .O(n51456));
    defparam n51453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36000 (.I0(byte_transmit_counter[1]), 
            .I1(n48752), .I2(n48753), .I3(byte_transmit_counter[2]), .O(n51447));
    defparam byte_transmit_counter_1__bdd_4_lut_36000.LUT_INIT = 16'he4aa;
    SB_LUT4 n51447_bdd_4_lut (.I0(n51447), .I1(n48855), .I2(n48854), .I3(byte_transmit_counter[2]), 
            .O(n51450));
    defparam n51447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35995 (.I0(byte_transmit_counter[1]), 
            .I1(n48812), .I2(n48813), .I3(byte_transmit_counter[2]), .O(n51441));
    defparam byte_transmit_counter_1__bdd_4_lut_35995.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1139 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n43633));
    defparam i1_2_lut_3_lut_adj_1139.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1140 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n43635));
    defparam i1_2_lut_3_lut_adj_1140.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1141 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n43637));
    defparam i1_2_lut_3_lut_adj_1141.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1142 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n43639));
    defparam i1_2_lut_3_lut_adj_1142.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n39145));
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\FRAME_MATCHER.state[0] ), .I1(n27958), 
            .I2(GND_net), .I3(GND_net), .O(n27874));   // verilog/coms.v(231[5:23])
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1144 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n43641));
    defparam i1_2_lut_3_lut_adj_1144.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1145 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n43643));
    defparam i1_2_lut_3_lut_adj_1145.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1146 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n43645));
    defparam i1_2_lut_3_lut_adj_1146.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1147 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n7_adj_4289));
    defparam i1_2_lut_3_lut_adj_1147.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1148 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n43647));
    defparam i1_2_lut_3_lut_adj_1148.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1149 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n43649));
    defparam i1_2_lut_3_lut_adj_1149.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1150 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n43651));
    defparam i1_2_lut_3_lut_adj_1150.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_1151 (.I0(n44408), .I1(n44722), .I2(n44456), 
            .I3(\data_out_frame[23] [4]), .O(n46058));
    defparam i3_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1152 (.I0(n44390), .I1(n44498), .I2(\data_out_frame[25] [7]), 
            .I3(n28588), .O(n12_adj_4399));
    defparam i5_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1153 (.I0(n45883), .I1(n12_adj_4399), .I2(n44753), 
            .I3(n45973), .O(n46218));
    defparam i6_4_lut_adj_1153.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1154 (.I0(\data_out_frame[24] [1]), .I1(n41591), 
            .I2(n44312), .I3(GND_net), .O(n14_adj_4400));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_adj_1154.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1155 (.I0(n44710), .I1(\data_out_frame[19] [6]), 
            .I2(\data_out_frame[24] [0]), .I3(n44640), .O(n15_adj_4401));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1156 (.I0(n15_adj_4401), .I1(n42428), .I2(n14_adj_4400), 
            .I3(\data_out_frame[23] [6]), .O(n45896));   // verilog/coms.v(71[16:27])
    defparam i8_4_lut_adj_1156.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1157 (.I0(n28583), .I1(n44489), .I2(n44437), 
            .I3(n41591), .O(n45973));
    defparam i3_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i16246_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n29773));
    defparam i16246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21680_2_lut_3_lut (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n35190));
    defparam i21680_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1158 (.I0(\data_out_frame[24] [2]), .I1(n44434), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4403));
    defparam i1_2_lut_adj_1158.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1159 (.I0(n41584), .I1(n44408), .I2(n28856), 
            .I3(n6_adj_4403), .O(n46761));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1160 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n43653));
    defparam i1_2_lut_3_lut_adj_1160.LUT_INIT = 16'he0e0;
    SB_LUT4 n51441_bdd_4_lut (.I0(n51441), .I1(n48852), .I2(n48851), .I3(byte_transmit_counter[2]), 
            .O(n51444));
    defparam n51441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35990 (.I0(byte_transmit_counter[1]), 
            .I1(n48842), .I2(n48843), .I3(byte_transmit_counter[2]), .O(n51435));
    defparam byte_transmit_counter_1__bdd_4_lut_35990.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1161 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n43655));
    defparam i1_2_lut_3_lut_adj_1161.LUT_INIT = 16'he0e0;
    SB_LUT4 i16247_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n29774));
    defparam i16247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1162 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n43657));
    defparam i1_2_lut_3_lut_adj_1162.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1163 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n7_adj_4287));
    defparam i1_2_lut_3_lut_adj_1163.LUT_INIT = 16'he0e0;
    SB_LUT4 i30_3_lut (.I0(n28849), .I1(n28855), .I2(\data_out_frame[24] [4]), 
            .I3(GND_net), .O(n41638));
    defparam i30_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i16248_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n29775));
    defparam i16248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1164 (.I0(\data_out_frame[17] [4]), .I1(n27608), 
            .I2(n44340), .I3(n28096), .O(n44643));
    defparam i3_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1165 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n43659));
    defparam i1_2_lut_3_lut_adj_1165.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1166 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n7_adj_4285));
    defparam i1_2_lut_3_lut_adj_1166.LUT_INIT = 16'he0e0;
    SB_LUT4 i16249_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n29776));
    defparam i16249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1167 (.I0(n44643), .I1(\data_out_frame[20] [0]), 
            .I2(n42428), .I3(n41638), .O(n14_adj_4404));
    defparam i6_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1168 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n43661));
    defparam i1_2_lut_3_lut_adj_1168.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1169 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n43663));
    defparam i1_2_lut_3_lut_adj_1169.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1170 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n43665));
    defparam i1_2_lut_3_lut_adj_1170.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1171 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n43667));
    defparam i1_2_lut_3_lut_adj_1171.LUT_INIT = 16'he0e0;
    SB_LUT4 i16250_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n29777));
    defparam i16250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1172 (.I0(\data_out_frame[24] [5]), .I1(n14_adj_4404), 
            .I2(n10_adj_4405), .I3(n28588), .O(n46786));
    defparam i7_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i16251_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n29778));
    defparam i16251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1173 (.I0(n169), .I1(n188), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n43669));
    defparam i1_2_lut_3_lut_adj_1173.LUT_INIT = 16'he0e0;
    SB_LUT4 i16230_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n29757));
    defparam i16230_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16252_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n29779));
    defparam i16252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1174 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28588));
    defparam i1_2_lut_adj_1174.LUT_INIT = 16'h6666;
    SB_LUT4 i16231_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n29758));
    defparam i16231_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1175 (.I0(n41575), .I1(n27564), .I2(\data_out_frame[24] [7]), 
            .I3(n42364), .O(n18_adj_4407));
    defparam i7_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1176 (.I0(n42394), .I1(n18_adj_4407), .I2(n44494), 
            .I3(n44590), .O(n20_adj_4408));
    defparam i9_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1177 (.I0(n44550), .I1(n28588), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4409));
    defparam i4_2_lut_adj_1177.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1178 (.I0(n15_adj_4409), .I1(n20_adj_4408), .I2(n42403), 
            .I3(n46040), .O(n45554));
    defparam i10_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44518));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\data_out_frame[23] [6]), .I1(n41659), 
            .I2(GND_net), .I3(GND_net), .O(n44722));
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1181 (.I0(\data_out_frame[25] [7]), .I1(\data_out_frame[25] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44456));
    defparam i1_2_lut_adj_1181.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1182 (.I0(\data_out_frame[15] [4]), .I1(n28468), 
            .I2(n42428), .I3(n44282), .O(n10_adj_4410));
    defparam i4_4_lut_adj_1182.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1183 (.I0(\data_out_frame[15] [3]), .I1(n10_adj_4410), 
            .I2(\data_out_frame[17] [5]), .I3(GND_net), .O(n28855));
    defparam i5_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i16232_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n29759));
    defparam i16232_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16233_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n29760));
    defparam i16233_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(n28855), .I1(n44798), .I2(GND_net), 
            .I3(GND_net), .O(n28856));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i16234_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n29761));
    defparam i16234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16235_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n29762));
    defparam i16235_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_out_frame[20] [5]), .I1(n44390), 
            .I2(GND_net), .I3(GND_net), .O(n28583));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i16236_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n29763));
    defparam i16236_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(n28855), .I1(\data_out_frame[20] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44707));
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1187 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [2]), 
            .I2(n44640), .I3(n6_adj_4411), .O(n45883));
    defparam i4_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1188 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[24] [5]), .I3(n28856), .O(n44550));
    defparam i3_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[23] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44489));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1190 (.I0(n41655), .I1(n44373), .I2(\data_out_frame[24] [0]), 
            .I3(GND_net), .O(n44753));
    defparam i2_3_lut_adj_1190.LUT_INIT = 16'h9696;
    SB_LUT4 i16237_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44156), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n29764));
    defparam i16237_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_3_lut (.I0(\data_out_frame[24] [3]), .I1(n44753), .I2(n44768), 
            .I3(GND_net), .O(n26_adj_4412));
    defparam i9_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i12_4_lut_adj_1191 (.I0(n44750), .I1(n44489), .I2(n44550), 
            .I3(n45883), .O(n29_adj_4413));
    defparam i12_4_lut_adj_1191.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1192 (.I0(n44722), .I1(n41571), .I2(n27722), 
            .I3(\data_out_frame[23] [5]), .O(n28_adj_4414));
    defparam i11_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1193 (.I0(n29_adj_4413), .I1(\data_out_frame[23] [0]), 
            .I2(n26_adj_4412), .I3(\data_out_frame[24] [4]), .O(n32_adj_4415));
    defparam i15_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1194 (.I0(n44581), .I1(n44518), .I2(n26118), 
            .I3(n28646), .O(n27_adj_4416));
    defparam i10_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1195 (.I0(n44215), .I1(n27_adj_4416), .I2(n32_adj_4415), 
            .I3(n28_adj_4414), .O(n7_adj_4417));   // verilog/coms.v(71[16:27])
    defparam i1_4_lut_adj_1195.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1196 (.I0(\data_out_frame[25] [5]), .I1(n7_adj_4417), 
            .I2(\data_out_frame[25] [4]), .I3(n8_adj_4418), .O(n41575));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 n51435_bdd_4_lut (.I0(n51435), .I1(n48849), .I2(n48848), .I3(byte_transmit_counter[2]), 
            .O(n51438));
    defparam n51435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16253_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44156), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n29780));
    defparam i16253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1197 (.I0(n27588), .I1(n41601), .I2(n27652), 
            .I3(n42439), .O(n10_adj_4419));
    defparam i4_4_lut_adj_1197.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1198 (.I0(n46263), .I1(n10_adj_4419), .I2(n41575), 
            .I3(GND_net), .O(n41916));
    defparam i5_3_lut_adj_1198.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1199 (.I0(n28849), .I1(n44798), .I2(GND_net), 
            .I3(GND_net), .O(n27564));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1199.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1200 (.I0(n44533), .I1(n41331), .I2(n41611), 
            .I3(n27564), .O(n44768));
    defparam i3_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1201 (.I0(n44768), .I1(\data_out_frame[20] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4420));
    defparam i2_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1202 (.I0(\data_out_frame[25] [0]), .I1(\data_out_frame[24] [6]), 
            .I2(n6_adj_4420), .I3(n42394), .O(n42364));
    defparam i1_4_lut_adj_1202.LUT_INIT = 16'h9669;
    SB_LUT4 i16238_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n29765));
    defparam i16238_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_out_frame[20] [7]), .I1(n46085), 
            .I2(GND_net), .I3(GND_net), .O(n42394));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h9999;
    SB_LUT4 i16239_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n29766));
    defparam i16239_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1204 (.I0(n44581), .I1(\data_out_frame[24] [7]), 
            .I2(n44494), .I3(GND_net), .O(n44533));
    defparam i2_3_lut_adj_1204.LUT_INIT = 16'h6969;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n30209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n30208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n30207));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n30206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n30205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n30204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n30203));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n30202));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n30201));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n30200));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n30199));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n30198));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n30197));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n30196));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n30195));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n30194));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n30193));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n30192));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n30191));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n30190));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n30189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n30188));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n30186));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n30185));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n30184));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n30183));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n30182));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n30181));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n30180));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n30179));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n30178));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n30177));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n30176));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n30175));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n30174));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n30173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n30172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n30171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n30170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n30169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n30168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n30167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n30166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n30165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n30164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n30163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n30162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n30161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n30160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n30159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n30158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n30157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n30156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n30155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n30154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n30153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n30152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n30151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n30150));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n30149));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n30148));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n30147));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n30146));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n30145));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n30144));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n30143));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n30141));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n30140));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n30139));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1205 (.I0(n46780), .I1(n28776), .I2(GND_net), 
            .I3(GND_net), .O(n44498));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(n42360), .I1(n44565), .I2(GND_net), 
            .I3(GND_net), .O(n28201));
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1207 (.I0(n28490), .I1(n44361), .I2(\data_out_frame[18] [1]), 
            .I3(\data_out_frame[16] [0]), .O(n12_adj_4422));
    defparam i5_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35985 (.I0(byte_transmit_counter[1]), 
            .I1(n48881), .I2(n48882), .I3(byte_transmit_counter[2]), .O(n51429));
    defparam byte_transmit_counter_1__bdd_4_lut_35985.LUT_INIT = 16'he4aa;
    SB_LUT4 i6_4_lut_adj_1208 (.I0(n28201), .I1(n12_adj_4422), .I2(n44655), 
            .I3(\data_out_frame[13] [6]), .O(n28849));
    defparam i6_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n30138));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n30137));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n30136));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n30135));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n30134));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n30133));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n30132));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n30131));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n30130));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1209 (.I0(n44287), .I1(n44463), .I2(\data_out_frame[18] [2]), 
            .I3(\data_out_frame[13] [6]), .O(n12_adj_4423));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1209.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1210 (.I0(n28884), .I1(n12_adj_4423), .I2(n44728), 
            .I3(\data_out_frame[13] [7]), .O(n28776));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n30129));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n30128));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n30127));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n30126));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n30125));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n30124));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n30123));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n30122));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n30121));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n30120));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n30119));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n30118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n30117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n30116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n30115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n30114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n30113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n30112));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n30111));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n30110));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n30109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n30108));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n30107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n30106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n30105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n30104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n30103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n30102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n30101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n30100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n30099));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1211 (.I0(n28776), .I1(n28849), .I2(GND_net), 
            .I3(GND_net), .O(n26118));
    defparam i1_2_lut_adj_1211.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n30098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n30097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n30096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n30095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n30094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n30093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n30092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n30091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n30090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n30089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n30088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n30087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n30086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n30085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n30084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n30083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n30082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n30081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n30080));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16240_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n29767));
    defparam i16240_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1212 (.I0(n44282), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[17] [3]), .I3(n44628), .O(n10_adj_4424));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n30079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n30078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n30077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n30076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n30075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n30074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n30073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n30072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n30071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n30070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n30069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n30068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n30067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n30066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n30065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n30064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n30063));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n30062));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n30061));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n30060));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n30059));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n30058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n30057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n30056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n30055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n30054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n30053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n30052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n30051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n30050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n30049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n30048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n30047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n30046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n30045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n30044));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n30043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n30042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n30041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n30040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n30039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n30038));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n30037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n30036));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n30035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n30034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n30033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n30032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n30031));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n30030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n30029));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n30028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n30027));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n30026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n30025));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n30024));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n30023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n30022));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n30021));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n30020));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n30019));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n30018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n30017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n30016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n30015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n30014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n30013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n30012));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(CLK_c), 
           .D(n30011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(CLK_c), 
           .D(n30009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(CLK_c), 
           .D(n30008));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n30007));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n30006));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n30005));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(CLK_c), 
           .D(n30004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n30003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n30002));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n30001));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n30000));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n29999));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n29998));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n29997));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n29996));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n29995));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(CLK_c), 
           .D(n29994));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(CLK_c), 
           .D(n29993));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n29992));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n29991));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(CLK_c), 
           .D(n29990));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n29989));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n29988));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n29987));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n29986));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n29985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n29984));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n29983));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n29982));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n29981));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n29980));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n29979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n29978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n29977));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n29976));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n29975));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1213 (.I0(\data_out_frame[19] [4]), .I1(n44271), 
            .I2(n10_adj_4424), .I3(\data_out_frame[15] [0]), .O(n44408));
    defparam i1_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n29974));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n29973));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n29972));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n29971));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n29970));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n29969));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_adj_1214 (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4425));
    defparam i2_2_lut_adj_1214.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1215 (.I0(\FRAME_MATCHER.state [8]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [14]), .I3(\FRAME_MATCHER.state [12]), 
            .O(n14_adj_4426));
    defparam i6_4_lut_adj_1215.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n29968));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1216 (.I0(\FRAME_MATCHER.state [10]), .I1(n14_adj_4426), 
            .I2(n10_adj_4425), .I3(\FRAME_MATCHER.state [11]), .O(n36247));
    defparam i7_4_lut_adj_1216.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_2_lut_adj_1217 (.I0(\FRAME_MATCHER.state [26]), .I1(\FRAME_MATCHER.state [29]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4427));
    defparam i4_2_lut_adj_1217.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n29967));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n29966));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n29965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1218 (.I0(n44450), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[13] [3]), .I3(n44631), .O(n10_adj_4428));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n29964));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n29963));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i218 (.Q(\data_out_frame[27][1] ), .C(CLK_c), 
           .D(n29962));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n29961));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n29960));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n29959));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n29958));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n29957));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n29956));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n29955));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n29954));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n29953));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n29952));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n29951));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n29950));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n29949));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n29948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n29947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n29946));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n29945));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n29944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n29943));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n29942));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n29941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n29940));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n29939));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_adj_1219 (.I0(n44387), .I1(n10_adj_4428), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n28468));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1219.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1220 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n44242));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4429));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1222 (.I0(n44319), .I1(\data_out_frame[15] [2]), 
            .I2(n44646), .I3(n6_adj_4429), .O(n44312));
    defparam i4_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i16241_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n29768));
    defparam i16241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[19] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44512));
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1224 (.I0(\data_out_frame[13] [5]), .I1(n28392), 
            .I2(n27665), .I3(n26043), .O(n41609));
    defparam i3_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28096));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1226 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[15] [4]), .I3(\data_out_frame[15] [5]), 
            .O(n44361));
    defparam i3_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n29931));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n29930));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_292_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4406));   // verilog/coms.v(154[7:23])
    defparam equal_292_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i3_4_lut_adj_1227 (.I0(\data_out_frame[7] [0]), .I1(n44840), 
            .I2(\data_out_frame[11] [2]), .I3(\data_out_frame[4] [6]), .O(n44631));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n29929));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n29928));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1228 (.I0(\data_out_frame[13] [4]), .I1(n44804), 
            .I2(n44290), .I3(\data_out_frame[6] [5]), .O(n10_adj_4430));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1229 (.I0(n44631), .I1(n10_adj_4430), .I2(\data_out_frame[8] [6]), 
            .I3(GND_net), .O(n44463));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1230 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[8] [6]), .I3(\data_out_frame[11] [1]), .O(n44450));   // verilog/coms.v(76[16:27])
    defparam i3_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 equal_293_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4421));   // verilog/coms.v(154[7:23])
    defparam equal_293_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44804));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1232 (.I0(n4_adj_4431), .I1(n103), .I2(n190), 
            .I3(\FRAME_MATCHER.state [16]), .O(n8_adj_4290));
    defparam i1_2_lut_4_lut_adj_1232.LUT_INIT = 16'hfe00;
    SB_LUT4 i16242_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n29769));
    defparam i16242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1233 (.I0(n44843), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[4] [4]), .I3(n44804), .O(n15_adj_4432));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1234 (.I0(n15_adj_4432), .I1(n44450), .I2(n14_adj_4433), 
            .I3(\data_out_frame[4] [1]), .O(n28658));   // verilog/coms.v(76[16:27])
    defparam i8_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 n51429_bdd_4_lut (.I0(n51429), .I1(n48837), .I2(n48836), .I3(byte_transmit_counter[2]), 
            .O(n51432));
    defparam n51429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35980 (.I0(byte_transmit_counter[1]), 
            .I1(n48884), .I2(n48885), .I3(byte_transmit_counter[2]), .O(n51423));
    defparam byte_transmit_counter_1__bdd_4_lut_35980.LUT_INIT = 16'he4aa;
    SB_LUT4 n51423_bdd_4_lut (.I0(n51423), .I1(n48834), .I2(n48833), .I3(byte_transmit_counter[2]), 
            .O(n51426));
    defparam n51423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16243_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n29770));
    defparam i16243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1235 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44719));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h6666;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(CLK_c), 
           .D(n43483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n29658));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n29657));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n29656));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n29654));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n29653));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n29652));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n29927));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1236 (.I0(\data_out_frame[12] [7]), .I1(n44719), 
            .I2(n44221), .I3(n44405), .O(n12_adj_4434));
    defparam i5_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n29926));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n29925));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n29924));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n29923));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n29922));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n29921));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n29920));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n29919));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n29918));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n29917));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n29916));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n29915));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n29914));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n29913));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n29912));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n29911));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n29910));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n29909));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n29908));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n29907));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n29906));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n29905));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n29904));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n29903));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n29902));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n29901));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n29900));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n29899));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n29898));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n29897));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16244_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n29771));
    defparam i16244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1237 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n46787));
    defparam i2_3_lut_adj_1237.LUT_INIT = 16'h9696;
    SB_LUT4 i16245_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44156), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n29772));
    defparam i16245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1238 (.I0(n46787), .I1(n12_adj_4434), .I2(\data_out_frame[13] [1]), 
            .I3(n44687), .O(n44282));
    defparam i6_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i22529_2_lut_4_lut (.I0(n4_adj_4431), .I1(n103), .I2(n190), 
            .I3(\FRAME_MATCHER.state [20]), .O(n36044));
    defparam i22529_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_adj_1239 (.I0(n44282), .I1(n1519), .I2(\data_out_frame[14] [7]), 
            .I3(n28078), .O(n44646));
    defparam i3_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1240 (.I0(n4_adj_4431), .I1(n103), .I2(n190), 
            .I3(\FRAME_MATCHER.state [24]), .O(n8_adj_4288));
    defparam i1_2_lut_4_lut_adj_1240.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1241 (.I0(n4_adj_4431), .I1(n103), .I2(n190), 
            .I3(\FRAME_MATCHER.state [26]), .O(n8_adj_4286));
    defparam i1_2_lut_4_lut_adj_1241.LUT_INIT = 16'hfe00;
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n29896));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n29895));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n29894));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n29893));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n29892));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n29891));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n29890));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n29889));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n29888));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n29887));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n29886));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n29885));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n29884));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n29883));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n29882));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n29881));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n29880));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n29879));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n29878));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n29877));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n29876));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n29875));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n29874));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n29873));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n29872));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n29871));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n29870));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n29869));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n29868));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n29867));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n29866));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n29865));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n29864));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n29863));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n29862));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n29861));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n29860));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n29859));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n29858));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n29857));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n29856));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n29855));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n29854));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n29853));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n29852));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n29851));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n29850));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n29849));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n29848));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n29847));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n29846));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n29845));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n29844));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n29843));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n29842));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n29841));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n29840));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n29839));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n29838));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n29837));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n29836));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n29835));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n29834));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\data_out_frame[13] [0]), .I1(n28658), 
            .I2(GND_net), .I3(GND_net), .O(n44340));
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n29833));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n29832));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n29831));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n29830));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n29829));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n29828));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n29827));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n29626));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n29625));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n29826));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n29825));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n29824));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n29823));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n29822));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n29821));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n29820));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n29819));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n29818));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n29817));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n29816));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n29815));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n29814));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n29813));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n29812));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n29811));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n29810));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n29809));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n29808));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n29807));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n29806));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n29805));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n29804));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n29803));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n29802));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n29801));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n29800));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n29799));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n29798));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n29797));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n29796));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n29795));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n29794));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n29793));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n29792));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n29791));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n29790));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n29789));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n29788));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n29787));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n29786));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n29785));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n29784));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n29783));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n29782));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1243 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44287));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1243.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(n41609), .I1(n28468), .I2(GND_net), 
            .I3(GND_net), .O(n44565));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h6666;
    SB_LUT4 i16398_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n29925));
    defparam i16398_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1245 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [1]), 
            .I2(n44565), .I3(\data_out_frame[16] [3]), .O(n30_adj_4435));
    defparam i11_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1246 (.I0(n28874), .I1(n30_adj_4435), .I2(n44556), 
            .I3(\data_out_frame[16] [2]), .O(n34_adj_4436));
    defparam i15_4_lut_adj_1246.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1247 (.I0(n44340), .I1(n41545), .I2(\data_out_frame[13] [5]), 
            .I3(n44646), .O(n32_adj_4437));
    defparam i13_4_lut_adj_1247.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1248 (.I0(n44463), .I1(n44249), .I2(n44334), 
            .I3(n42180), .O(n33));
    defparam i14_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1249 (.I0(n28531), .I1(n44309), .I2(n1516), 
            .I3(n44807), .O(n31_adj_4438));
    defparam i12_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1250 (.I0(n31_adj_4438), .I1(n33), .I2(n32_adj_4437), 
            .I3(n34_adj_4436), .O(n46648));
    defparam i18_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1251 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[17] [4]), 
            .I2(n44361), .I3(n46648), .O(n22_adj_4439));
    defparam i9_4_lut_adj_1251.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1252 (.I0(n28096), .I1(\data_out_frame[17] [6]), 
            .I2(n44625), .I3(\data_out_frame[17] [0]), .O(n21_adj_4440));
    defparam i8_4_lut_adj_1252.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1253 (.I0(n41791), .I1(\data_out_frame[17] [5]), 
            .I2(n41609), .I3(n14_adj_4441), .O(n23));
    defparam i10_4_lut_adj_1253.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1254 (.I0(n44437), .I1(n23), .I2(n21_adj_4440), 
            .I3(n22_adj_4439), .O(n15_adj_4442));
    defparam i3_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1255 (.I0(n44512), .I1(n44312), .I2(n28713), 
            .I3(n44565), .O(n19_adj_4443));
    defparam i7_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1256 (.I0(n19_adj_4443), .I1(n15_adj_4442), .I2(n44725), 
            .I3(n44559), .O(n22_adj_4444));
    defparam i10_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1257 (.I0(n44509), .I1(n22_adj_4444), .I2(n18_adj_4445), 
            .I3(n44408), .O(n46085));
    defparam i11_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(n41659), .I1(n46085), .I2(GND_net), 
            .I3(GND_net), .O(n44731));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h9999;
    SB_LUT4 i16399_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n29926));
    defparam i16399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1259 (.I0(n44559), .I1(\data_out_frame[23] [1]), 
            .I2(\data_out_frame[23] [0]), .I3(n44731), .O(n10_adj_4446));
    defparam i4_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1260 (.I0(\data_out_frame[20] [5]), .I1(n10_adj_4446), 
            .I2(n46040), .I3(GND_net), .O(n27652));
    defparam i5_3_lut_adj_1260.LUT_INIT = 16'h6969;
    SB_LUT4 i16400_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n29927));
    defparam i16400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16129_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n29656));
    defparam i16129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44215));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1262 (.I0(n42439), .I1(n44215), .I2(n27652), 
            .I3(GND_net), .O(n45552));
    defparam i2_3_lut_adj_1262.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1263 (.I0(\data_out_frame[4] [3]), .I1(n44259), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n27665));
    defparam i2_3_lut_adj_1263.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44728));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1265 (.I0(n44828), .I1(\data_out_frame[16] [2]), 
            .I2(n44502), .I3(\data_out_frame[15] [7]), .O(n14_adj_4447));
    defparam i6_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i16401_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n29928));
    defparam i16401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1266 (.I0(\data_out_frame[18] [3]), .I1(n14_adj_4447), 
            .I2(n10_adj_4448), .I3(n28490), .O(n46780));
    defparam i7_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1267 (.I0(\data_out_frame[20] [6]), .I1(n27722), 
            .I2(n42403), .I3(GND_net), .O(n41611));
    defparam i2_3_lut_adj_1267.LUT_INIT = 16'h6969;
    SB_LUT4 i16402_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n29929));
    defparam i16402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16403_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n29930));
    defparam i16403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(n41541), .I1(n46780), .I2(GND_net), 
            .I3(GND_net), .O(n28141));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[23] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44750));
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1270 (.I0(n28141), .I1(n45757), .I2(n41611), 
            .I3(\data_out_frame[20] [5]), .O(n44492));
    defparam i3_4_lut_adj_1270.LUT_INIT = 16'h9669;
    SB_LUT4 i16404_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44169), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n29931));
    defparam i16404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1271 (.I0(\data_out_frame[5] [1]), .I1(n44795), 
            .I2(n44615), .I3(n44230), .O(n26043));
    defparam i3_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1272 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[13] [7]), .I3(GND_net), .O(n44828));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1272.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1273 (.I0(\data_out_frame[14] [0]), .I1(n44473), 
            .I2(n44265), .I3(\data_out_frame[11] [6]), .O(n28884));
    defparam i3_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(n28884), .I1(n44828), .I2(GND_net), 
            .I3(GND_net), .O(n44334));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(\data_out_frame[11] [4]), .I1(n26043), 
            .I2(GND_net), .I3(GND_net), .O(n44655));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1276 (.I0(n42433), .I1(\data_out_frame[16] [2]), 
            .I2(n44334), .I3(n6_adj_4449), .O(n41541));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1276.LUT_INIT = 16'h9669;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n39182), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1277 (.I0(n41541), .I1(n44537), .I2(\data_out_frame[18] [5]), 
            .I3(GND_net), .O(n42403));
    defparam i2_3_lut_adj_1277.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1278 (.I0(\FRAME_MATCHER.state [30]), .I1(\FRAME_MATCHER.state [19]), 
            .I2(\FRAME_MATCHER.state [28]), .I3(\FRAME_MATCHER.state [18]), 
            .O(n24_adj_4450));
    defparam i10_4_lut_adj_1278.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n39181), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1279 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[23] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n28646));
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(\data_out_frame[25] [4]), .I1(n46263), 
            .I2(GND_net), .I3(GND_net), .O(n41636));
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h9999;
    SB_CARRY add_3971_8 (.CI(n39181), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n39182));
    SB_LUT4 i3_4_lut_adj_1281 (.I0(n41636), .I1(n28646), .I2(n41940), 
            .I3(\data_out_frame[25] [5]), .O(n45837));
    defparam i3_4_lut_adj_1281.LUT_INIT = 16'h9669;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n39180), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 equal_290_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4451));   // verilog/coms.v(154[7:23])
    defparam equal_290_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i8_4_lut_adj_1282 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [21]), .I3(\FRAME_MATCHER.state [31]), 
            .O(n22_adj_4452));
    defparam i8_4_lut_adj_1282.LUT_INIT = 16'hfffe;
    SB_CARRY add_3971_7 (.CI(n39180), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n39181));
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n39179), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_6 (.CI(n39179), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n39180));
    SB_LUT4 i12_4_lut_adj_1283 (.I0(\FRAME_MATCHER.state [17]), .I1(n24_adj_4450), 
            .I2(n18_adj_4427), .I3(\FRAME_MATCHER.state [20]), .O(n26_adj_4453));
    defparam i12_4_lut_adj_1283.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n39178), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_5 (.CI(n39178), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n39179));
    SB_LUT4 equal_298_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4454));   // verilog/coms.v(154[7:23])
    defparam equal_298_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n1510), .I1(\data_out_frame[12] [2]), 
            .I2(n1513), .I3(\data_out_frame[12] [3]), .O(n44249));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n39177), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_4 (.CI(n39177), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n39178));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n39176), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_3_lut_4_lut_adj_1284 (.I0(n1510), .I1(\data_out_frame[12] [2]), 
            .I2(n28078), .I3(n10_adj_4455), .O(n44459));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_3 (.CI(n39176), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n39177));
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3513), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_3_lut_4_lut_adj_1285 (.I0(n27572), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[14] [2]), .I3(n28388), .O(n14_adj_4456));
    defparam i5_3_lut_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3513), 
            .CO(n39176));
    SB_LUT4 i1_2_lut_3_lut_adj_1286 (.I0(n44492), .I1(\data_out_frame[23] [1]), 
            .I2(\data_out_frame[23] [2]), .I3(GND_net), .O(n42439));
    defparam i1_2_lut_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1287 (.I0(n27572), .I1(\data_out_frame[12] [1]), 
            .I2(n1519), .I3(n28531), .O(n44380));
    defparam i2_3_lut_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1288 (.I0(\FRAME_MATCHER.state [2]), .I1(n27866), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2626 ));
    defparam i1_2_lut_3_lut_adj_1288.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_4_lut_adj_1289 (.I0(n41659), .I1(n4_adj_4457), .I2(\data_out_frame[20] [7]), 
            .I3(n44492), .O(n44494));
    defparam i1_2_lut_4_lut_adj_1289.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(\FRAME_MATCHER.state [2]), .I1(n27866), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n82));
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n29781));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16390_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n29917));
    defparam i16390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_33_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n39175), .O(n2_adj_4305)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_32_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n39174), .O(n2_adj_4307)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n39174), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n39175));
    SB_LUT4 add_43_31_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n39173), .O(n2_adj_4309)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n39173), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n39174));
    SB_LUT4 i16391_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n29918));
    defparam i16391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16392_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n29919));
    defparam i16392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16393_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n29920));
    defparam i16393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16394_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n29921));
    defparam i16394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16395_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n29922));
    defparam i16395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1291 (.I0(n44696), .I1(\data_out_frame[11] [5]), 
            .I2(\data_out_frame[12] [0]), .I3(n44681), .O(n15_adj_4459));
    defparam i6_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1292 (.I0(n15_adj_4459), .I1(n44268), .I2(n14_adj_4460), 
            .I3(\data_out_frame[5] [3]), .O(n42180));
    defparam i8_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1293 (.I0(n1513), .I1(n42180), .I2(n44735), .I3(n1673), 
            .O(n10_adj_4461));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i16396_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n29923));
    defparam i16396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1294 (.I0(n1519), .I1(n10_adj_4461), .I2(n1516), 
            .I3(GND_net), .O(n44502));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_1294.LUT_INIT = 16'h9696;
    SB_LUT4 i16397_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44169), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n29924));
    defparam i16397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1295 (.I0(\data_out_frame[16] [5]), .I1(n44249), 
            .I2(\data_out_frame[14] [4]), .I3(n41531), .O(n41791));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1296 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(n44693), .I3(n44420), .O(n44268));
    defparam i2_3_lut_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1297 (.I0(\data_out_frame[16] [3]), .I1(n41545), 
            .I2(\data_out_frame[14] [1]), .I3(n42433), .O(n45757));
    defparam i3_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1298 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [3]), .I3(n1191), .O(n28041));
    defparam i2_3_lut_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_30_lut (.I0(n2987), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n39172), .O(n2_adj_4311)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44625));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1300 (.I0(n44420), .I1(n44696), .I2(n28041), 
            .I3(\data_out_frame[11] [5]), .O(n28490));
    defparam i1_2_lut_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44290));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1302 (.I0(n44420), .I1(n44696), .I2(n28041), 
            .I3(n28392), .O(n31_adj_4462));
    defparam i1_2_lut_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1303 (.I0(n44634), .I1(\data_out_frame[8] [3]), 
            .I2(n44262), .I3(\data_out_frame[8] [5]), .O(n14_adj_4463));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1304 (.I0(\data_out_frame[10] [6]), .I1(n14_adj_4463), 
            .I2(n10_adj_4464), .I3(\data_out_frame[4] [3]), .O(n27608));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1305 (.I0(\data_out_frame[5] [7]), .I1(n44649), 
            .I2(n44322), .I3(\data_out_frame[10] [1]), .O(n1513));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n29780));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n29779));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1306 (.I0(\data_out_frame[12] [6]), .I1(n29039), 
            .I2(\data_out_frame[17] [2]), .I3(n6_adj_4465), .O(n44271));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1307 (.I0(\FRAME_MATCHER.state [23]), .I1(n22_adj_4452), 
            .I2(\FRAME_MATCHER.state [27]), .I3(GND_net), .O(n25_adj_4466));
    defparam i11_3_lut_adj_1307.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n29778));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1308 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[16] [7]), 
            .I2(n8_adj_4467), .I3(n44625), .O(n44437));
    defparam i1_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_CARRY add_43_30 (.CI(n39172), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n39173));
    SB_LUT4 i1_4_lut_adj_1309 (.I0(n25_adj_4466), .I1(\FRAME_MATCHER.state [24]), 
            .I2(n26_adj_4453), .I3(\FRAME_MATCHER.state [16]), .O(n36381));
    defparam i1_4_lut_adj_1309.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1310 (.I0(\data_out_frame[19] [2]), .I1(n29054), 
            .I2(n44476), .I3(n44459), .O(n44710));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1311 (.I0(\FRAME_MATCHER.state [5]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n36029));
    defparam i3_4_lut_adj_1311.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n29777));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n29776));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n29775));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n29774));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n29773));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n29772));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n29771));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n29770));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n29769));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n29768));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n29767));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16382_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n29909));
    defparam i16382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n29766));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n28078));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n29765));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1313 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44634));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h6666;
    SB_LUT4 i16383_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n29910));
    defparam i16383_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16384_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n29911));
    defparam i16384_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1314 (.I0(\data_out_frame[12] [3]), .I1(n44470), 
            .I2(n44309), .I3(\data_out_frame[12] [5]), .O(n1673));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44681));
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44687));
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1317 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(n44687), .I3(n44681), .O(n10_adj_4468));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i16385_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n29912));
    defparam i16385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1318 (.I0(\data_out_frame[10] [5]), .I1(n10_adj_4468), 
            .I2(n44262), .I3(GND_net), .O(n44319));   // verilog/coms.v(73[16:42])
    defparam i5_3_lut_adj_1318.LUT_INIT = 16'h9696;
    SB_LUT4 i16386_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n29913));
    defparam i16386_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1319 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n44230));
    defparam i2_3_lut_adj_1319.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1320 (.I0(n28041), .I1(n28045), .I2(\data_out_frame[4] [5]), 
            .I3(n6_adj_4469), .O(n44696));   // verilog/coms.v(71[16:62])
    defparam i4_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n28392));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'h6666;
    SB_LUT4 i16387_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n29914));
    defparam i16387_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(71[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44840));
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'h6666;
    SB_LUT4 i16388_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n29915));
    defparam i16388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44795));
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1324 (.I0(n44795), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[8] [7]), .I3(n44840), .O(n10_adj_4470));
    defparam i4_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i16389_3_lut_4_lut (.I0(n8), .I1(n44169), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n29916));
    defparam i16389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_287_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_287_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i5_3_lut_adj_1325 (.I0(\data_out_frame[7] [1]), .I1(n10_adj_4470), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n44259));
    defparam i5_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 equal_278_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4402));   // verilog/coms.v(154[7:23])
    defparam equal_278_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_3_lut_adj_1326 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n44387));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1327 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44843));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1327.LUT_INIT = 16'h6666;
    SB_LUT4 i17915_3_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n35517));
    defparam i17915_3_lut_3_lut.LUT_INIT = 16'hdada;
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27958), .I3(GND_net), .O(n27866));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35975 (.I0(byte_transmit_counter[1]), 
            .I1(n49705), .I2(n49706), .I3(byte_transmit_counter[2]), .O(n51405));
    defparam byte_transmit_counter_1__bdd_4_lut_35975.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44693));
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1329 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44420));
    defparam i1_2_lut_adj_1329.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_4_lut_adj_1330 (.I0(\data_out_frame[12] [3]), .I1(n1513), 
            .I2(n44271), .I3(\data_out_frame[14] [5]), .O(n8_adj_4467));   // verilog/coms.v(74[16:43])
    defparam i3_3_lut_4_lut_adj_1330.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1331 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n44615));
    defparam i2_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44405));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h6666;
    SB_LUT4 i22_4_lut_adj_1333 (.I0(\data_out_frame[9] [5]), .I1(n44405), 
            .I2(\data_out_frame[10] [1]), .I3(n29027), .O(n52_adj_4471));   // verilog/coms.v(85[17:63])
    defparam i22_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1334 (.I0(\data_out_frame[9] [3]), .I1(n44615), 
            .I2(n44678), .I3(n44268), .O(n50_adj_4472));   // verilog/coms.v(85[17:63])
    defparam i20_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1335 (.I0(n44221), .I1(n28045), .I2(\data_out_frame[4] [5]), 
            .I3(n28104), .O(n51));   // verilog/coms.v(85[17:63])
    defparam i21_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 n51405_bdd_4_lut (.I0(n51405), .I1(n17_adj_4256), .I2(n16_adj_4255), 
            .I3(byte_transmit_counter[2]), .O(n51408));
    defparam n51405_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19_4_lut_adj_1336 (.I0(\data_out_frame[7] [6]), .I1(n44259), 
            .I2(n44649), .I3(\data_out_frame[4] [2]), .O(n49_adj_4473));   // verilog/coms.v(85[17:63])
    defparam i19_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1337 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[4] [3]), 
            .I2(n44387), .I3(\data_out_frame[6] [4]), .O(n32_adj_4474));   // verilog/coms.v(85[17:63])
    defparam i2_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i16374_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n29901));
    defparam i16374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_1338 (.I0(\data_out_frame[11] [2]), .I1(n1191), 
            .I2(\data_out_frame[11] [1]), .I3(n44328), .O(n48));   // verilog/coms.v(85[17:63])
    defparam i18_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1339 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(n44668), .I3(n1673), .O(n47));   // verilog/coms.v(85[17:63])
    defparam i17_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n49_adj_4473), .I1(n51), .I2(n50_adj_4472), 
            .I3(n52_adj_4471), .O(n58_adj_4475));   // verilog/coms.v(85[17:63])
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1340 (.I0(\data_out_frame[10] [2]), .I1(n31_adj_4462), 
            .I2(\data_out_frame[10] [6]), .I3(n32_adj_4474), .O(n53_adj_4476));   // verilog/coms.v(85[17:63])
    defparam i23_4_lut_adj_1340.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n53_adj_4476), .I1(n58_adj_4475), .I2(n47), 
            .I3(n48), .O(n27574));   // verilog/coms.v(85[17:63])
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44556));
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h6666;
    SB_LUT4 i16375_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n29902));
    defparam i16375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(n27574), .I1(n44319), .I2(GND_net), 
            .I3(GND_net), .O(n41523));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\data_out_frame[14] [7]), .I1(n27574), 
            .I2(GND_net), .I3(GND_net), .O(n29039));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n29027));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1345 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[6] [1]), .I3(GND_net), .O(n44678));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44377));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h6666;
    SB_LUT4 i16376_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n29903));
    defparam i16376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1347 (.I0(n44377), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[5] [5]), .I3(n44678), .O(n10_adj_4477));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28531));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1349 (.I0(n29039), .I1(n41523), .I2(\data_out_frame[17] [1]), 
            .I3(n44556), .O(n10_adj_4455));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1350 (.I0(n36029), .I1(n36381), .I2(n36247), 
            .I3(GND_net), .O(n27958));   // verilog/coms.v(231[5:23])
    defparam i2_3_lut_adj_1350.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28713));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1352 (.I0(n44380), .I1(n44459), .I2(\data_out_frame[14] [3]), 
            .I3(GND_net), .O(n44725));
    defparam i2_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 i16377_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n29904));
    defparam i16377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1353 (.I0(\FRAME_MATCHER.state [2]), .I1(n27866), 
            .I2(GND_net), .I3(GND_net), .O(n103_adj_4478));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1353.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1354 (.I0(n4_adj_4479), .I1(\data_out_frame[20] [7]), 
            .I2(n41659), .I3(GND_net), .O(n27722));
    defparam i2_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1355 (.I0(n44710), .I1(\data_out_frame[23] [5]), 
            .I2(n44437), .I3(GND_net), .O(n41655));
    defparam i2_3_lut_adj_1355.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1356 (.I0(n1510), .I1(n27572), .I2(GND_net), 
            .I3(GND_net), .O(n44735));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1356.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35960 (.I0(byte_transmit_counter[1]), 
            .I1(n49708), .I2(n49709), .I3(byte_transmit_counter[2]), .O(n51399));
    defparam byte_transmit_counter_1__bdd_4_lut_35960.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1357 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44470));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1357.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1358 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n28104));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1358.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1359 (.I0(\data_out_frame[9] [4]), .I1(n28104), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[7] [2]), .O(n44265));
    defparam i3_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1360 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[12] [0]), 
            .I2(\data_out_frame[11] [7]), .I3(GND_net), .O(n44668));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1361 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n44738));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n28045));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h6666;
    SB_LUT4 i16378_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n29905));
    defparam i16378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16379_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n29906));
    defparam i16379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1363 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44358));
    defparam i1_2_lut_adj_1363.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1364 (.I0(n28388), .I1(n44473), .I2(\data_out_frame[7] [6]), 
            .I3(\data_out_frame[10] [0]), .O(n12_adj_4480));
    defparam i5_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1365 (.I0(\data_out_frame[11] [7]), .I1(n12_adj_4480), 
            .I2(n44738), .I3(\data_out_frame[5] [5]), .O(n27572));
    defparam i6_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i16380_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n29907));
    defparam i16380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1366 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(n44358), .I3(n44668), .O(n15_adj_4481));
    defparam i6_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1367 (.I0(n15_adj_4481), .I1(n44265), .I2(n14_adj_4456), 
            .I3(\data_out_frame[9] [6]), .O(n41545));
    defparam i8_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i16381_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44169), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n29908));
    defparam i16381_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1368 (.I0(n44470), .I1(n44735), .I2(\data_out_frame[14] [3]), 
            .I3(GND_net), .O(n41531));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1369 (.I0(\data_out_frame[16] [4]), .I1(n41531), 
            .I2(n41545), .I3(GND_net), .O(n44537));
    defparam i2_3_lut_adj_1369.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1370 (.I0(n41791), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[18] [6]), .I3(n28141), .O(n44559));
    defparam i1_2_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1371 (.I0(n41791), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[18] [6]), .I3(n45757), .O(n4_adj_4479));
    defparam i1_2_lut_4_lut_adj_1371.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_1372 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[10] [3]), .I3(\data_out_frame[6] [1]), .O(n12_adj_4482));   // verilog/coms.v(85[17:70])
    defparam i5_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1373 (.I0(\data_out_frame[8] [2]), .I1(n12_adj_4482), 
            .I2(n44322), .I3(\data_out_frame[4] [0]), .O(n1516));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1374 (.I0(n1516), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44628));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1374.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1375 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n44328));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1375.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1376 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n28805));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1376.LUT_INIT = 16'h6666;
    SB_LUT4 i16366_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n29893));
    defparam i16366_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1377 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[10] [0]), 
            .I2(n28805), .I3(\data_out_frame[10] [1]), .O(n12_adj_4483));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1378 (.I0(\data_out_frame[5] [6]), .I1(n12_adj_4483), 
            .I2(n44328), .I3(\data_out_frame[5] [2]), .O(n1510));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 i16367_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n29894));
    defparam i16367_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1379 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44476));
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1380 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n29054));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1380.LUT_INIT = 16'h9696;
    SB_LUT4 i16368_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n29895));
    defparam i16368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16369_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n29896));
    defparam i16369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16370_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n29897));
    defparam i16370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1381 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(n44537), .I3(\data_out_frame[16] [6]), .O(n14_adj_4484));
    defparam i6_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1382 (.I0(\data_out_frame[19] [0]), .I1(n14_adj_4484), 
            .I2(n10_adj_4485), .I3(n44628), .O(n41659));
    defparam i7_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i16371_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n29898));
    defparam i16371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16372_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n29899));
    defparam i16372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33396_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48833));
    defparam i33396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1383 (.I0(\data_out_frame[19] [1]), .I1(n41659), 
            .I2(n29054), .I3(n28874), .O(n12_adj_4486));
    defparam i5_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1384 (.I0(\data_out_frame[18] [7]), .I1(n12_adj_4486), 
            .I2(\data_out_frame[23] [3]), .I3(n44380), .O(n44762));
    defparam i6_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1385 (.I0(n44590), .I1(n44762), .I2(GND_net), 
            .I3(GND_net), .O(n41601));
    defparam i1_2_lut_adj_1385.LUT_INIT = 16'h6666;
    SB_LUT4 i33397_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48834));
    defparam i33397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16373_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44169), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n29900));
    defparam i16373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33448_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48885));
    defparam i33448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16358_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n29885));
    defparam i16358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16359_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n29886));
    defparam i16359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16360_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n29887));
    defparam i16360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i16361_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n29888));
    defparam i16361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16362_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n29889));
    defparam i16362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16363_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n29890));
    defparam i16363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16364_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n29891));
    defparam i16364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16365_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44169), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n29892));
    defparam i16365_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33447_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48884));
    defparam i33447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33399_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48836));
    defparam i33399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33400_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n48837));
    defparam i33400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1386 (.I0(n4_adj_4457), .I1(n4_adj_4479), 
            .I2(\data_out_frame[23] [2]), .I3(n44762), .O(n46263));
    defparam i2_3_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1387 (.I0(\FRAME_MATCHER.i_31__N_2626 ), .I1(\FRAME_MATCHER.i_31__N_2624 ), 
            .I2(n82), .I3(GND_net), .O(n2987));
    defparam i2_3_lut_adj_1387.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_1388 (.I0(n4_adj_4457), .I1(n4_adj_4479), 
            .I2(\data_out_frame[23] [0]), .I3(n44533), .O(n27588));
    defparam i2_3_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1389 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(\data_out_frame[20] [3]), .I3(\data_out_frame[20] [4]), 
            .O(n44390));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(n42403), .I3(GND_net), .O(n4_adj_4457));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i16350_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n29877));
    defparam i16350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16351_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n29878));
    defparam i16351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16352_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n29879));
    defparam i16352_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16353_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n29880));
    defparam i16353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16354_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n29881));
    defparam i16354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16355_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n29882));
    defparam i16355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16356_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n29883));
    defparam i16356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16357_3_lut_4_lut (.I0(n10_adj_4454), .I1(n44163), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n29884));
    defparam i16357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(\data_out_frame[11] [3]), .I1(n27665), 
            .I2(\data_out_frame[15] [4]), .I3(n44463), .O(n42360));
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i16342_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n29869));
    defparam i16342_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16343_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n29870));
    defparam i16343_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n51399_bdd_4_lut (.I0(n51399), .I1(n17_adj_4254), .I2(n16_adj_4253), 
            .I3(byte_transmit_counter[2]), .O(n51402));
    defparam n51399_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16344_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n29871));
    defparam i16344_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16345_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n29872));
    defparam i16345_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16346_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n29873));
    defparam i16346_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_adj_1392 (.I0(\FRAME_MATCHER.state_31__N_2724 [3]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.i_31__N_2621 ), .I3(n44186), .O(n43691));
    defparam i1_4_lut_adj_1392.LUT_INIT = 16'heca0;
    SB_LUT4 i29743_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n44134), .I2(n103_adj_4478), 
            .I3(n45036), .O(n45105));
    defparam i29743_4_lut.LUT_INIT = 16'ha8aa;
    SB_LUT4 i1_4_lut_adj_1393 (.I0(\FRAME_MATCHER.state [3]), .I1(n188), 
            .I2(n44062), .I3(n45105), .O(n43485));
    defparam i1_4_lut_adj_1393.LUT_INIT = 16'h88a8;
    SB_LUT4 i16347_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n29874));
    defparam i16347_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35955 (.I0(byte_transmit_counter[1]), 
            .I1(n49711), .I2(n49712), .I3(byte_transmit_counter[2]), .O(n51393));
    defparam byte_transmit_counter_1__bdd_4_lut_35955.LUT_INIT = 16'he4aa;
    SB_LUT4 i16348_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n29875));
    defparam i16348_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16349_3_lut_4_lut (.I0(n10_adj_4454), .I1(n45615), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n29876));
    defparam i16349_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16334_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n29861));
    defparam i16334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1394 (.I0(\FRAME_MATCHER.state [4]), .I1(n11_adj_4487), 
            .I2(GND_net), .I3(GND_net), .O(n43489));
    defparam i1_2_lut_adj_1394.LUT_INIT = 16'h8888;
    SB_LUT4 n51393_bdd_4_lut (.I0(n51393), .I1(n17_adj_4251), .I2(n16_adj_4249), 
            .I3(byte_transmit_counter[2]), .O(n51396));
    defparam n51393_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16335_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n29862));
    defparam i16335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35950 (.I0(byte_transmit_counter[1]), 
            .I1(n49717), .I2(n49718), .I3(byte_transmit_counter[2]), .O(n51387));
    defparam byte_transmit_counter_1__bdd_4_lut_35950.LUT_INIT = 16'he4aa;
    SB_LUT4 i16336_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n29863));
    defparam i16336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16337_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n29864));
    defparam i16337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16338_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n29865));
    defparam i16338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n51387_bdd_4_lut (.I0(n51387), .I1(n17_adj_4248), .I2(n16_adj_4247), 
            .I3(byte_transmit_counter[2]), .O(n51390));
    defparam n51387_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i16339_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n29866));
    defparam i16339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16340_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n29867));
    defparam i16340_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(\FRAME_MATCHER.state [8]), .I1(n11_adj_4487), 
            .I2(GND_net), .I3(GND_net), .O(n43509));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h8888;
    SB_LUT4 i29701_2_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n36247), 
            .I2(n36381), .I3(n36029), .O(n45062));
    defparam i29701_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35901_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n29452));
    defparam i35901_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i22272_2_lut_4_lut (.I0(n25324), .I1(n31_adj_4230), .I2(n31), 
            .I3(\FRAME_MATCHER.state [1]), .O(n1_c));
    defparam i22272_2_lut_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i16341_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44176), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n29868));
    defparam i16341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1396 (.I0(\FRAME_MATCHER.state [10]), .I1(n11_adj_4487), 
            .I2(GND_net), .I3(GND_net), .O(n43493));
    defparam i1_2_lut_adj_1396.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1397 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [0]), 
            .I2(n44602), .I3(\data_in_frame[0] [1]), .O(n44331));   // verilog/coms.v(70[16:62])
    defparam i1_2_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(\data_out_frame[25] [1]), .I1(n27588), 
            .I2(n42364), .I3(GND_net), .O(n44577));
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1399 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[9] [3]), .I3(n41577), .O(n44578));
    defparam i1_2_lut_3_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1400 (.I0(\data_out_frame[25] [1]), .I1(n27588), 
            .I2(\data_out_frame[25] [2]), .I3(n27652), .O(n45583));
    defparam i2_3_lut_4_lut_adj_1400.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1401 (.I0(n28289), .I1(\data_in_frame[8] [3]), 
            .I2(n44296), .I3(n44416), .O(n28349));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1402 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [3]), 
            .I2(n46780), .I3(n28849), .O(n44581));
    defparam i2_3_lut_4_lut_adj_1402.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1403 (.I0(\FRAME_MATCHER.state [11]), .I1(n11_adj_4487), 
            .I2(GND_net), .I3(GND_net), .O(n43505));
    defparam i1_2_lut_adj_1403.LUT_INIT = 16'h8888;
    SB_LUT4 i29680_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n27958), .I3(\FRAME_MATCHER.state [3]), .O(n45036));
    defparam i29680_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1404 (.I0(n28658), .I1(\data_out_frame[17] [6]), 
            .I2(n44242), .I3(n28201), .O(n44798));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1405 (.I0(n28658), .I1(\data_out_frame[17] [6]), 
            .I2(n42360), .I3(n44512), .O(n42428));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1406 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(\FRAME_MATCHER.state[0] ), .I2(n27958), .I3(\FRAME_MATCHER.state [1]), 
            .O(n7_adj_4241));
    defparam i1_2_lut_3_lut_4_lut_adj_1406.LUT_INIT = 16'hfffe;
    SB_LUT4 i16326_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n29853));
    defparam i16326_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16327_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n29854));
    defparam i16327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16328_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n29855));
    defparam i16328_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16329_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n29856));
    defparam i16329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29578_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n44134), .I2(n45036), 
            .I3(GND_net), .O(n44934));
    defparam i29578_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1_4_lut_adj_1407 (.I0(n31443), .I1(n44183), .I2(n44934), 
            .I3(n44062), .O(n11_adj_4487));
    defparam i1_4_lut_adj_1407.LUT_INIT = 16'hcdcc;
    SB_LUT4 i16330_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n29857));
    defparam i16330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1408 (.I0(\FRAME_MATCHER.state [12]), .I1(n11_adj_4487), 
            .I2(GND_net), .I3(GND_net), .O(n43513));
    defparam i1_2_lut_adj_1408.LUT_INIT = 16'h8888;
    SB_LUT4 i16331_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n29858));
    defparam i16331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1409 (.I0(\data_out_frame[19] [6]), .I1(n28776), 
            .I2(n28849), .I3(\data_out_frame[20] [3]), .O(n10_adj_4405));
    defparam i2_2_lut_3_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(n41659), .I1(n4_adj_4457), .I2(\data_out_frame[20] [7]), 
            .I3(GND_net), .O(n41571));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i16332_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n29859));
    defparam i16332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1410 (.I0(n2987), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_4451), 
            .O(n44176));
    defparam i1_2_lut_3_lut_4_lut_adj_1410.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1411 (.I0(n2987), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_4454), 
            .O(n44169));
    defparam i1_2_lut_3_lut_4_lut_adj_1411.LUT_INIT = 16'hfff7;
    SB_LUT4 i16333_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44176), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n29860));
    defparam i16333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16318_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n29845));
    defparam i16318_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1412 (.I0(n2987), .I1(n25063), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n7_adj_4241), .O(n44062));
    defparam i2_3_lut_4_lut_adj_1412.LUT_INIT = 16'h4404;
    SB_LUT4 i21673_2_lut_3_lut (.I0(n2987), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n35182));
    defparam i21673_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(n169), .I1(n103), .I2(n4_adj_4431), 
            .I3(GND_net), .O(n44186));
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1414 (.I0(\data_out_frame[11] [3]), .I1(n27665), 
            .I2(\data_out_frame[13] [5]), .I3(\data_out_frame[16] [1]), 
            .O(n10_adj_4448));
    defparam i2_2_lut_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i16319_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n29846));
    defparam i16319_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1415 (.I0(n44590), .I1(n44762), .I2(\data_out_frame[25] [5]), 
            .I3(\data_out_frame[25] [6]), .O(n46112));
    defparam i2_3_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i16320_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n29847));
    defparam i16320_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut_adj_1416 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n45062), .O(n29310));
    defparam i3_3_lut_4_lut_adj_1416.LUT_INIT = 16'h0010;
    SB_LUT4 i16321_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n29848));
    defparam i16321_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1417 (.I0(n44710), .I1(\data_out_frame[23] [5]), 
            .I2(n44437), .I3(n41940), .O(n44590));
    defparam i1_2_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i16322_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n29849));
    defparam i16322_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[14] [5]), .I3(GND_net), .O(n28874));
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[10] [2]), .I3(\data_out_frame[6] [0]), .O(n44322));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1420 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[7] [3]), .O(n28388));
    defparam i2_3_lut_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n27866), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2624 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'h0404;
    SB_LUT4 i2_3_lut_4_lut_adj_1422 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[9] [5]), .I3(\data_out_frame[5] [3]), .O(n44473));
    defparam i2_3_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1423 (.I0(n27722), .I1(n44725), .I2(n28713), 
            .I3(\data_out_frame[18] [7]), .O(n41940));
    defparam i1_2_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i16323_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n29850));
    defparam i16323_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16324_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n29851));
    defparam i16324_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1424 (.I0(\data_out_frame[8] [1]), .I1(n10_adj_4477), 
            .I2(\data_out_frame[10] [3]), .I3(\data_out_frame[10] [4]), 
            .O(n1519));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1425 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[8] [3]), .O(n44221));
    defparam i2_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1426 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[5] [3]), .O(n44649));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1427 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[9] [3]), .I3(\data_out_frame[6] [7]), .O(n6_adj_4469));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1428 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[8] [2]), .I3(n1191), .O(n44262));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1429 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n44309));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1430 (.I0(\data_out_frame[13] [0]), .I1(n27608), 
            .I2(\data_out_frame[14] [6]), .I3(n41523), .O(n6_adj_4465));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1431 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[10] [4]), .I3(GND_net), .O(n10_adj_4464));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_3_lut_adj_1431.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1432 (.I0(\data_out_frame[13] [7]), .I1(n1519), 
            .I2(n10_adj_4461), .I3(n1516), .O(n42433));
    defparam i1_2_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1433 (.I0(\data_out_frame[4] [0]), .I1(n1673), 
            .I2(\data_out_frame[8] [3]), .I3(\data_out_frame[4] [1]), .O(n14_adj_4460));
    defparam i5_3_lut_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1434 (.I0(n1510), .I1(\data_out_frame[12] [2]), 
            .I2(\data_out_frame[14] [4]), .I3(\data_out_frame[14] [5]), 
            .O(n10_adj_4485));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(n26043), .I3(GND_net), .O(n6_adj_4449));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i16325_3_lut_4_lut (.I0(n8), .I1(n44176), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n29852));
    defparam i16325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1436 (.I0(n44492), .I1(n44750), .I2(\data_out_frame[25] [3]), 
            .I3(n41636), .O(n45838));
    defparam i2_3_lut_4_lut_adj_1436.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1437 (.I0(n41331), .I1(n46780), .I2(n28776), 
            .I3(\data_out_frame[20] [4]), .O(n46040));
    defparam i2_3_lut_4_lut_adj_1437.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1438 (.I0(n44434), .I1(n44707), .I2(\data_out_frame[20] [0]), 
            .I3(n28588), .O(n41591));
    defparam i1_2_lut_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i6_2_lut_4_lut (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(\data_out_frame[19] [5]), 
            .O(n18_adj_4445));
    defparam i6_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1439 (.I0(n44434), .I1(n44707), .I2(\data_out_frame[20] [0]), 
            .I3(\data_out_frame[24] [3]), .O(n41584));
    defparam i1_2_lut_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1440 (.I0(n44312), .I1(n44643), .I2(n45973), 
            .I3(n44518), .O(n46120));
    defparam i2_3_lut_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1441 (.I0(n44312), .I1(n44643), .I2(\data_out_frame[20] [2]), 
            .I3(n28904), .O(n44434));
    defparam i2_3_lut_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1442 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[17] [3]), .I3(GND_net), .O(n14_adj_4441));
    defparam i1_2_lut_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1443 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[11] [0]), .O(n14_adj_4433));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i16310_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n29837));
    defparam i16310_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16311_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n29838));
    defparam i16311_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1444 (.I0(\data_out_frame[19] [6]), .I1(n28776), 
            .I2(n28849), .I3(GND_net), .O(n44509));
    defparam i1_2_lut_3_lut_adj_1444.LUT_INIT = 16'h9696;
    SB_LUT4 i16312_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n29839));
    defparam i16312_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16313_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n29840));
    defparam i16313_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1445 (.I0(n41659), .I1(n46085), .I2(n4_adj_4457), 
            .I3(GND_net), .O(n41331));
    defparam i2_2_lut_3_lut_adj_1445.LUT_INIT = 16'h6969;
    SB_LUT4 i16314_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n29841));
    defparam i16314_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1446 (.I0(n46263), .I1(n10_adj_4419), .I2(n41575), 
            .I3(n42364), .O(n28794));
    defparam i1_2_lut_4_lut_adj_1446.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1447 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[25] [6]), .I3(GND_net), .O(n8_adj_4418));   // verilog/coms.v(71[16:27])
    defparam i2_2_lut_3_lut_adj_1447.LUT_INIT = 16'h9696;
    SB_LUT4 i16315_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n29842));
    defparam i16315_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16316_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n29843));
    defparam i16316_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16317_3_lut_4_lut (.I0(n8_adj_4402), .I1(n44176), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n29844));
    defparam i16317_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16302_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n29829));
    defparam i16302_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16303_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n29830));
    defparam i16303_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1448 (.I0(n35205), .I1(n70), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n27874), .O(n45660));
    defparam i3_4_lut_adj_1448.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1449 (.I0(n46780), .I1(n28776), .I2(n28855), 
            .I3(\data_out_frame[20] [1]), .O(n6_adj_4411));
    defparam i1_2_lut_4_lut_adj_1449.LUT_INIT = 16'h9669;
    SB_LUT4 i16304_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n29831));
    defparam i16304_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16305_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n29832));
    defparam i16305_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16306_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n29833));
    defparam i16306_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16307_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n29834));
    defparam i16307_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16308_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n29835));
    defparam i16308_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16309_3_lut_4_lut (.I0(n8_adj_4421), .I1(n44176), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n29836));
    defparam i16309_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_622_Select_1_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4352));
    defparam select_622_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_2_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4350));
    defparam select_622_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[19] [5]), 
            .I2(\data_out_frame[20] [5]), .I3(n44390), .O(n44640));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'h6996;
    SB_LUT4 select_622_Select_3_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4348));
    defparam select_622_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_4_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4346));
    defparam select_622_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[20] [5]), 
            .I2(n44390), .I3(GND_net), .O(n28904));
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 select_622_Select_5_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4344));
    defparam select_622_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_6_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4342));
    defparam select_622_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_7_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4340));
    defparam select_622_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_8_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4338));
    defparam select_622_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_9_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4336));
    defparam select_622_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_10_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4334));
    defparam select_622_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_11_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4332));
    defparam select_622_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i2_3_lut_4_lut_adj_1452 (.I0(\data_out_frame[20] [5]), .I1(n44390), 
            .I2(n41638), .I3(n41584), .O(n45780));
    defparam i2_3_lut_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 select_622_Select_12_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4330));
    defparam select_622_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_13_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4328));
    defparam select_622_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_14_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4326));
    defparam select_622_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_15_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4325));
    defparam select_622_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_16_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4324));
    defparam select_622_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_17_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4323));
    defparam select_622_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_18_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4322));
    defparam select_622_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_19_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4321));
    defparam select_622_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_20_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4320));
    defparam select_622_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_21_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4319));
    defparam select_622_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_22_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4318));
    defparam select_622_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_23_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4317));
    defparam select_622_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_24_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4316));
    defparam select_622_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 mux_1817_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[19] [1]), .O(n6561));
    defparam mux_1817_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_622_Select_25_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4315));
    defparam select_622_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_26_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4314));
    defparam select_622_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_27_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4313));
    defparam select_622_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 mux_1817_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[19] [2]), .O(n6562));
    defparam mux_1817_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1817_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[19] [3]), .O(n6563));
    defparam mux_1817_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i29561_2_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n27958), .O(n44134));
    defparam i29561_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 select_622_Select_28_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4312));
    defparam select_622_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 mux_1817_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[19] [4]), .O(n6564));
    defparam mux_1817_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_622_Select_29_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4310));
    defparam select_622_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 mux_1817_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[19] [5]), .O(n6565));
    defparam mux_1817_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 select_622_Select_30_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4308));
    defparam select_622_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 mux_1817_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[19] [6]), .O(n6566));
    defparam mux_1817_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1453 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[18] [1]), .I3(\data_in_frame[10] [7]), .O(n6_adj_4395));
    defparam i1_2_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 select_622_Select_31_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4306));
    defparam select_622_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_622_Select_0_i3_2_lut_4_lut (.I0(n2987), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n7_adj_4241), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_622_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i3_3_lut_4_lut_adj_1454 (.I0(n46645), .I1(n42347), .I2(\data_in_frame[19] [7]), 
            .I3(\data_in_frame[19] [6]), .O(n12_adj_4394));   // verilog/coms.v(85[17:28])
    defparam i3_3_lut_4_lut_adj_1454.LUT_INIT = 16'h9669;
    SB_LUT4 i4_3_lut_4_lut (.I0(n44416), .I1(\data_in_frame[15] [1]), .I2(\data_in_frame[14] [7]), 
            .I3(n28264), .O(n14_adj_4375));
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1455 (.I0(n28289), .I1(\data_in_frame[8] [3]), 
            .I2(n44296), .I3(GND_net), .O(n28313));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1455.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1456 (.I0(\data_in_frame[4] [0]), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n44256));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1456.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n6_adj_4364));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1458 (.I0(n28289), .I1(\data_in_frame[8] [2]), 
            .I2(n28160), .I3(\data_in_frame[10] [4]), .O(n44416));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[19] [7]), .O(n6567));
    defparam mux_1817_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1459 (.I0(n28289), .I1(\data_in_frame[8] [2]), 
            .I2(n28160), .I3(GND_net), .O(n4_adj_4229));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1459.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1460 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[3] [5]), .I3(GND_net), .O(n44495));
    defparam i1_2_lut_3_lut_adj_1460.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1461 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [6]), .O(n44293));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1462 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n28843));
    defparam i1_2_lut_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1463 (.I0(n44725), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[19] [1]), .I3(\data_out_frame[18] [7]), 
            .O(n44373));
    defparam i2_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1464 (.I0(\data_in_frame[5] [0]), .I1(n4_c), 
            .I2(n29017), .I3(GND_net), .O(n44453));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1464.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1465 (.I0(n35182), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n44156));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1465.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_3_lut_4_lut_adj_1466 (.I0(n27608), .I1(\data_out_frame[14] [6]), 
            .I2(n27574), .I3(n44319), .O(n44807));
    defparam i2_3_lut_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1467 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [7]), 
            .I2(\data_in_frame[6] [6]), .I3(\data_in_frame[6] [1]), .O(n44831));
    defparam i2_3_lut_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1468 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [3]), 
            .I2(n10_adj_4353), .I3(\data_in_frame[5] [7]), .O(n28796));   // verilog/coms.v(74[16:27])
    defparam i5_3_lut_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[18] [0]), .O(n6568));
    defparam mux_1817_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1469 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[7] [7]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[5] [5]), .O(n44413));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n44744));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i16294_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n29821));
    defparam i16294_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16295_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n29822));
    defparam i16295_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1471 (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(n25063), 
            .I2(n3303), .I3(GND_net), .O(n4_adj_4431));
    defparam i1_3_lut_adj_1471.LUT_INIT = 16'h0808;
    SB_LUT4 i16296_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n29823));
    defparam i16296_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1472 (.I0(n771), .I1(n82), .I2(n25063), .I3(GND_net), 
            .O(n103));   // verilog/coms.v(115[11:12])
    defparam i1_3_lut_adj_1472.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1473 (.I0(n103), .I1(n4_adj_4431), .I2(GND_net), 
            .I3(GND_net), .O(n44183));
    defparam i1_2_lut_adj_1473.LUT_INIT = 16'heeee;
    SB_LUT4 i189_2_lut (.I0(n25063), .I1(n45880), .I2(GND_net), .I3(GND_net), 
            .O(n190));
    defparam i189_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1474 (.I0(\data_in_frame[8] [7]), .I1(\data_in_frame[6] [5]), 
            .I2(n44658), .I3(GND_net), .O(n28837));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_3_lut_adj_1474.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1817_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[18] [1]), .O(n6569));
    defparam mux_1817_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16297_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n29824));
    defparam i16297_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[18] [2]), .O(n6570));
    defparam mux_1817_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i187_3_lut (.I0(\FRAME_MATCHER.i_31__N_2626 ), .I1(n4452), .I2(n25063), 
            .I3(GND_net), .O(n188));   // verilog/coms.v(115[11:12])
    defparam i187_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i2_3_lut_4_lut_adj_1475 (.I0(n28736), .I1(\data_in_frame[12] [7]), 
            .I2(n28289), .I3(n44637), .O(n44343));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1476 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[7] [0]), .I3(n28624), .O(n44431));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1477 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[2] [6]), 
            .I2(n44384), .I3(GND_net), .O(n29057));
    defparam i1_2_lut_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1478 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(n29060), .I3(GND_net), .O(n28840));
    defparam i1_2_lut_3_lut_adj_1478.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1479 (.I0(n28445), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n44652));
    defparam i1_2_lut_3_lut_adj_1479.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1817_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[18] [3]), .O(n6571));
    defparam mux_1817_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_4_lut_adj_1480 (.I0(\data_in_frame[10] [7]), .I1(n28719), 
            .I2(\data_in_frame[15] [2]), .I3(\data_in_frame[11] [0]), .O(n44661));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[18] [4]), .O(n6572));
    defparam mux_1817_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16298_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n29825));
    defparam i16298_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16299_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n29826));
    defparam i16299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16300_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n29827));
    defparam i16300_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[18] [5]), .O(n6573));
    defparam mux_1817_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16301_3_lut_4_lut (.I0(n8_adj_4406), .I1(n44176), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n29828));
    defparam i16301_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(n28313), .I1(n44416), .I2(n28753), 
            .I3(\data_in_frame[12] [5]), .O(n28264));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1482 (.I0(Kp_23__N_1217), .I1(\data_in_frame[7] [0]), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[9] [1]), .O(n28655));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1483 (.I0(\data_in_frame[2] [6]), .I1(n44349), 
            .I2(Kp_23__N_981), .I3(n29060), .O(n28342));
    defparam i2_3_lut_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48781), .I3(n48779), .O(n7_adj_4360));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48823), .I3(n48821), .O(n7_adj_4359));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48817), .I3(n48815), .O(n7_adj_4304));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48808), .I3(n48806), .O(n7_adj_4303));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48802), .I3(n48800), .O(n7_adj_4302));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 mux_1817_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[18] [6]), .O(n6574));
    defparam mux_1817_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1817_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[18] [7]), .O(n6575));
    defparam mux_1817_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48796), .I3(n48794), .O(n7_adj_4301));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48784), .I3(n48782), .O(n7_adj_4299));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 mux_1817_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[17] [0]), .O(n6576));
    defparam mux_1817_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n48790), .I3(n48788), .O(n7_adj_4300));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i16286_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n29813));
    defparam i16286_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16287_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n29814));
    defparam i16287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1484 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n28342), .I3(n28347), .O(n27552));
    defparam i2_3_lut_4_lut_adj_1484.LUT_INIT = 16'h6996;
    SB_LUT4 i16288_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n29815));
    defparam i16288_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16289_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n29816));
    defparam i16289_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[17] [1]), .O(n6577));
    defparam mux_1817_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_1817_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[17] [2]), .O(n6578));
    defparam mux_1817_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16290_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n29817));
    defparam i16290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1485 (.I0(\data_in_frame[7] [6]), .I1(n28238), 
            .I2(n44834), .I3(GND_net), .O(n28347));
    defparam i1_2_lut_3_lut_adj_1485.LUT_INIT = 16'h9696;
    SB_LUT4 i16291_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n29818));
    defparam i16291_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16292_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n29819));
    defparam i16292_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16293_3_lut_4_lut (.I0(n10_adj_4451), .I1(n44163), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n29820));
    defparam i16293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16278_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n29805));
    defparam i16278_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16279_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n29806));
    defparam i16279_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_1817_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[17] [3]), .O(n6579));
    defparam mux_1817_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16280_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n29807));
    defparam i16280_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_1817_i21_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[17] [4]), .O(n6580));
    defparam mux_1817_i21_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_3_lut_4_lut_adj_1486 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_988), 
            .I2(n28445), .I3(Kp_23__N_981), .O(n8_adj_4279));
    defparam i3_3_lut_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1487 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [3]), 
            .I2(n41577), .I3(GND_net), .O(n41622));
    defparam i1_2_lut_3_lut_adj_1487.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1488 (.I0(n44671), .I1(n44367), .I2(n27552), 
            .I3(\data_in_frame[10] [0]), .O(n44524));
    defparam i1_2_lut_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1489 (.I0(\data_in_frame[7] [1]), .I1(Kp_23__N_1228), 
            .I2(n44578), .I3(GND_net), .O(n42356));
    defparam i1_2_lut_3_lut_adj_1489.LUT_INIT = 16'h9696;
    SB_LUT4 i16281_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n29808));
    defparam i16281_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[12] [0]), .I3(GND_net), .O(n18_adj_4276));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1490 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[14] [7]), 
            .I2(n28264), .I3(GND_net), .O(n44252));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1490.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1491 (.I0(n42341), .I1(n28753), .I2(\data_in_frame[12] [4]), 
            .I3(\data_in_frame[14] [6]), .O(n44540));
    defparam i1_2_lut_4_lut_adj_1491.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1492 (.I0(\data_in_frame[16] [6]), .I1(n28235), 
            .I2(n44505), .I3(GND_net), .O(n6_adj_4265));
    defparam i2_2_lut_3_lut_adj_1492.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1493 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n27866), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2623 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1493.LUT_INIT = 16'h0808;
    SB_LUT4 i16282_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n29809));
    defparam i16282_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_1817_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[17] [5]), .O(n6581));
    defparam mux_1817_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_3_lut_4_lut_adj_1494 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n6), .O(n8_adj_4234));
    defparam i3_3_lut_4_lut_adj_1494.LUT_INIT = 16'hff7f;
    SB_LUT4 i16283_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n29810));
    defparam i16283_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i29531_4_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n27958), .I3(n2_adj_4488), .O(n44882));
    defparam i29531_4_lut_4_lut.LUT_INIT = 16'hfdf8;
    SB_LUT4 i1_2_lut_3_lut_adj_1495 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n2_adj_4488));
    defparam i1_2_lut_3_lut_adj_1495.LUT_INIT = 16'ha8a8;
    SB_LUT4 i16284_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n29811));
    defparam i16284_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i16285_3_lut_4_lut (.I0(n10_adj_4451), .I1(n45615), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n29812));
    defparam i16285_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_1817_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[17] [6]), .O(n6582));
    defparam mux_1817_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1496 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[4] [1]), .I3(GND_net), .O(n44611));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1496.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1497 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n27958), .O(n36505));
    defparam i2_3_lut_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1498 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[6] [1]), .O(n44622));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1817_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[17] [7]), .O(n6583));
    defparam mux_1817_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16270_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n29797));
    defparam i16270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16271_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n29798));
    defparam i16271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1817_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n35205), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[19] [0]), .O(n6560));
    defparam mux_1817_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i16272_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n29799));
    defparam i16272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16273_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n29800));
    defparam i16273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16274_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n29801));
    defparam i16274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16275_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n29802));
    defparam i16275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16276_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n29803));
    defparam i16276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1499 (.I0(\data_in_frame[11] [1]), .I1(n44837), 
            .I2(\data_in_frame[10] [5]), .I3(n44343), .O(n44813));
    defparam i1_2_lut_3_lut_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i16277_3_lut_4_lut (.I0(n8_adj_4217), .I1(n44156), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n29804));
    defparam i16277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16262_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n29789));
    defparam i16262_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16263_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n29790));
    defparam i16263_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1500 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n6935));
    defparam i1_2_lut_3_lut_adj_1500.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_3_lut_adj_1501 (.I0(n63_adj_4224), .I1(n63_adj_4221), 
            .I2(n63), .I3(GND_net), .O(n25063));   // verilog/coms.v(136[7:86])
    defparam i1_2_lut_3_lut_adj_1501.LUT_INIT = 16'h8080;
    SB_LUT4 i16264_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n29791));
    defparam i16264_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35945 (.I0(byte_transmit_counter[1]), 
            .I1(n49720), .I2(n49721), .I3(byte_transmit_counter[2]), .O(n51381));
    defparam byte_transmit_counter_1__bdd_4_lut_35945.LUT_INIT = 16'he4aa;
    SB_LUT4 n51381_bdd_4_lut (.I0(n51381), .I1(n17_adj_4245), .I2(n16_adj_4244), 
            .I3(byte_transmit_counter[2]), .O(n51384));
    defparam n51381_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35940 (.I0(byte_transmit_counter[1]), 
            .I1(n49723), .I2(n49724), .I3(byte_transmit_counter[2]), .O(n51375));
    defparam byte_transmit_counter_1__bdd_4_lut_35940.LUT_INIT = 16'he4aa;
    SB_LUT4 n51375_bdd_4_lut (.I0(n51375), .I1(n17_adj_4242), .I2(n16_adj_4240), 
            .I3(byte_transmit_counter[2]), .O(n51378));
    defparam n51375_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35935 (.I0(byte_transmit_counter[1]), 
            .I1(n49726), .I2(n49727), .I3(byte_transmit_counter[2]), .O(n51369));
    defparam byte_transmit_counter_1__bdd_4_lut_35935.LUT_INIT = 16'he4aa;
    SB_LUT4 n51369_bdd_4_lut (.I0(n51369), .I1(n17_adj_4238), .I2(n16_adj_4237), 
            .I3(byte_transmit_counter[2]), .O(n51372));
    defparam n51369_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_35930 (.I0(byte_transmit_counter[1]), 
            .I1(n49729), .I2(n49730), .I3(byte_transmit_counter[2]), .O(n51363));
    defparam byte_transmit_counter_1__bdd_4_lut_35930.LUT_INIT = 16'he4aa;
    SB_LUT4 n51363_bdd_4_lut (.I0(n51363), .I1(n17_adj_4236), .I2(n16_adj_4235), 
            .I3(byte_transmit_counter[2]), .O(n51366));
    defparam n51363_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_650_Select_1_i1_3_lut_4_lut (.I0(n123), .I1(n82), .I2(n63), 
            .I3(n771), .O(n1));
    defparam select_650_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'h3323;
    SB_LUT4 i1_3_lut_adj_1502 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n18_adj_4490));
    defparam i1_3_lut_adj_1502.LUT_INIT = 16'h8484;
    SB_LUT4 i4_4_lut_adj_1503 (.I0(Kp_23__N_981), .I1(Kp_23__N_974), .I2(\data_in_frame[2] [6]), 
            .I3(\data_in_frame[1] [0]), .O(n21_adj_4491));
    defparam i4_4_lut_adj_1503.LUT_INIT = 16'h2184;
    SB_LUT4 i1_3_lut_4_lut_adj_1504 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n27981), .I3(\FRAME_MATCHER.i [1]), .O(n5));
    defparam i1_3_lut_4_lut_adj_1504.LUT_INIT = 16'hfefc;
    SB_LUT4 i16265_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n29792));
    defparam i16265_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1505 (.I0(n29017), .I1(n44599), .I2(n44602), 
            .I3(\data_in_frame[0] [5]), .O(n20_adj_4492));
    defparam i3_4_lut_adj_1505.LUT_INIT = 16'h4114;
    SB_LUT4 i13_4_lut_adj_1506 (.I0(n48504), .I1(\data_in_frame[2] [0]), 
            .I2(n18_adj_4490), .I3(n44331), .O(n30_adj_4493));
    defparam i13_4_lut_adj_1506.LUT_INIT = 16'h4010;
    SB_LUT4 i11_4_lut_adj_1507 (.I0(n21_adj_4491), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [4]), .I3(n44331), .O(n28_adj_4494));
    defparam i11_4_lut_adj_1507.LUT_INIT = 16'h2080;
    SB_LUT4 i12_4_lut_adj_1508 (.I0(\data_in_frame[1] [3]), .I1(n25324), 
            .I2(\data_in_frame[1] [6]), .I3(n28445), .O(n29_adj_4495));
    defparam i12_4_lut_adj_1508.LUT_INIT = 16'h0020;
    SB_LUT4 i10_4_lut_adj_1509 (.I0(\data_in_frame[1] [2]), .I1(n20_adj_4492), 
            .I2(Kp_23__N_977), .I3(\data_in_frame[2] [2]), .O(n27_adj_4496));
    defparam i10_4_lut_adj_1509.LUT_INIT = 16'h8008;
    SB_LUT4 i16_4_lut_adj_1510 (.I0(n27_adj_4496), .I1(n29_adj_4495), .I2(n28_adj_4494), 
            .I3(n30_adj_4493), .O(\FRAME_MATCHER.state_31__N_2724 [3]));
    defparam i16_4_lut_adj_1510.LUT_INIT = 16'h8000;
    SB_LUT4 i35908_4_lut (.I0(n45066), .I1(\FRAME_MATCHER.state [3]), .I2(n35343), 
            .I3(n29452), .O(n46485));
    defparam i35908_4_lut.LUT_INIT = 16'h0501;
    SB_LUT4 i16266_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n29793));
    defparam i16266_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1511 (.I0(n1_c), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state_31__N_2724 [3]), 
            .O(n15_adj_4497));
    defparam i1_4_lut_adj_1511.LUT_INIT = 16'ha0ac;
    SB_LUT4 i1_4_lut_adj_1512 (.I0(n44882), .I1(n15_adj_4497), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(n36505), .O(n4_adj_4498));
    defparam i1_4_lut_adj_1512.LUT_INIT = 16'haeaa;
    SB_LUT4 i35310_4_lut (.I0(n29452), .I1(n4_adj_4498), .I2(n36505), 
            .I3(\FRAME_MATCHER.state [3]), .O(n46541));
    defparam i35310_4_lut.LUT_INIT = 16'h2223;
    SB_LUT4 i1_2_lut_3_lut_adj_1513 (.I0(n63_adj_4224), .I1(n63_adj_4221), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n123));   // verilog/coms.v(136[7:86])
    defparam i1_2_lut_3_lut_adj_1513.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_adj_1514 (.I0(n36247), .I1(n36381), .I2(n36029), 
            .I3(GND_net), .O(n45024));
    defparam i2_3_lut_adj_1514.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_280_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4458));
    defparam equal_280_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i16267_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n29794));
    defparam i16267_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16268_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n29795));
    defparam i16268_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24_4_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n13));
    defparam i24_4_lut_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i29705_2_lut (.I0(n44882), .I1(n45062), .I2(GND_net), .I3(GND_net), 
            .O(n45066));
    defparam i29705_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_281_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4217));
    defparam equal_281_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i35905_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n45066), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(\FRAME_MATCHER.state [1]), .O(n46530));
    defparam i35905_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut_adj_1515 (.I0(\FRAME_MATCHER.state[0] ), .I1(n45024), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n45517));
    defparam i2_3_lut_adj_1515.LUT_INIT = 16'h1010;
    SB_LUT4 i35911_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n44882), .I3(n45517), .O(n46735));
    defparam i35911_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i35301_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n88));
    defparam i35301_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i16269_3_lut_4_lut (.I0(n8_adj_4458), .I1(n44156), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n29796));
    defparam i16269_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1516 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n35182), .O(n45615));
    defparam i2_3_lut_4_lut_adj_1516.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_adj_1517 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[6] [3]), .I3(GND_net), .O(n44596));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1517.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1518 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[6] [5]), 
            .I2(n44399), .I3(Kp_23__N_1096), .O(n28719));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1518.LUT_INIT = 16'h6996;
    uart_tx tx (.CLK_c(CLK_c), .n29234(n29234), .\r_SM_Main_2__N_3613[1] (\r_SM_Main_2__N_3613[1] ), 
            .r_SM_Main({r_SM_Main}), .GND_net(GND_net), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .tx_o(tx_o), .tx_data({tx_data}), .n44068(n44068), .n29667(n29667), 
            .n29662(n29662), .tx_active(tx_active), .n51668(n51668), .VCC_net(VCC_net), 
            .\r_SM_Main_2__N_3616[0] (r_SM_Main_2__N_3616[0]), .n20400(n20400), 
            .n4(n4_adj_6), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.CLK_c(CLK_c), .n29246(n29246), .r_Rx_Data(r_Rx_Data), 
            .r_SM_Main({r_SM_Main_adj_14}), .GND_net(GND_net), .RX_N_10(RX_N_10), 
            .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_10 ), .n44059(n44059), 
            .\r_SM_Main_2__N_3542[2] (\r_SM_Main_2__N_3542[2] ), .n27976(n27976), 
            .n4(n4_adj_11), .n29679(n29679), .rx_data({rx_data}), .n29672(n29672), 
            .n43733(n43733), .rx_data_ready(rx_data_ready), .n29650(n29650), 
            .n29649(n29649), .n29648(n29648), .n29647(n29647), .n29646(n29646), 
            .n29645(n29645), .n29644(n29644), .n44138(n44138), .VCC_net(VCC_net), 
            .n4_adj_4(n4_adj_12), .n4_adj_5(n4_adj_13), .n27971(n27971), 
            .n35414(n35414)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (CLK_c, n29234, \r_SM_Main_2__N_3613[1] , r_SM_Main, 
            GND_net, \r_Bit_Index[0] , tx_o, tx_data, n44068, n29667, 
            n29662, tx_active, n51668, VCC_net, \r_SM_Main_2__N_3616[0] , 
            n20400, n4, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output n29234;
    output \r_SM_Main_2__N_3613[1] ;
    output [2:0]r_SM_Main;
    input GND_net;
    output \r_Bit_Index[0] ;
    output tx_o;
    input [7:0]tx_data;
    output n44068;
    input n29667;
    input n29662;
    output tx_active;
    input n51668;
    input VCC_net;
    input \r_SM_Main_2__N_3616[0] ;
    output n20400;
    output n4;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]n41;
    
    wire n6852;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n29528;
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n29492, n21286, n21287, o_Tx_Serial_N_3644, n3;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n48839, n48840, n25095, n48846, n48845, n3_adj_4210;
    wire [2:0]r_SM_Main_2__N_3610;
    
    wire n51471, n40523, n40522, n40521, n40520, n40519, n40518, 
        n40517, n40516, n46462, n10;
    
    SB_DFFESR r_Clock_Count_2065__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n6852), 
            .D(n41[8]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n6852), 
            .D(n41[7]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n6852), 
            .D(n41[6]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n6852), 
            .D(n41[5]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n6852), 
            .D(n41[4]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n6852), 
            .D(n41[3]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n6852), 
            .D(n41[2]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n6852), 
            .D(n41[1]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2065__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n6852), 
            .D(n41[0]), .R(n29528));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n29234), 
            .D(n307[1]), .R(n29492));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n29234), 
            .D(n307[2]), .R(n29492));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i7900_3_lut (.I0(n21286), .I1(\r_SM_Main_2__N_3613[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21287));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7900_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3644), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i33402_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48839));
    defparam i33402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33403_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48840));
    defparam i33403_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n6852), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n25095), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n21287), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i33409_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48846));
    defparam i33409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33408_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n48845));
    defparam i33408_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4210), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n25095), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n25095), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2200_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2200_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n44068));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n25095), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n25095), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n25095), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n25095), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n25095), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i22580_2_lut (.I0(n44068), .I1(\r_SM_Main_2__N_3613[1] ), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3610[0]));
    defparam i22580_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2193_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2193_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n48845), 
            .I2(n48846), .I3(r_Bit_Index[2]), .O(n51471));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51471_bdd_4_lut (.I0(n51471), .I1(n48840), .I2(n48839), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_3644));
    defparam n51471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i11355_2_lut_3_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4210));
    defparam i11355_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n29667));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n29662));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n51668));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_2065_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n40523), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2065_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n40522), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_9 (.CI(n40522), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n40523));
    SB_LUT4 r_Clock_Count_2065_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n40521), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_8 (.CI(n40521), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n40522));
    SB_LUT4 r_Clock_Count_2065_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n40520), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_7 (.CI(n40520), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n40521));
    SB_LUT4 r_Clock_Count_2065_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n40519), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_6 (.CI(n40519), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n40520));
    SB_LUT4 r_Clock_Count_2065_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n40518), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_5 (.CI(n40518), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n40519));
    SB_LUT4 r_Clock_Count_2065_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n40517), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_4 (.CI(n40517), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n40518));
    SB_LUT4 r_Clock_Count_2065_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n40516), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_3 (.CI(n40516), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n40517));
    SB_LUT4 r_Clock_Count_2065_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2065_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2065_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n40516));
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n46462));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7018_2_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n20400));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7018_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n46462), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3613[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i35194_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3613[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n29528));
    defparam i35194_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3616[0] ), 
            .I3(r_SM_Main[1]), .O(n25095));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3610[0]), .O(n29492));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_869 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3613[1] ), .O(n29234));
    defparam i1_3_lut_4_lut_adj_869.LUT_INIT = 16'h1101;
    SB_LUT4 i1985_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n6852));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1985_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i7899_3_lut_4_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(n44068), 
            .I2(\r_SM_Main_2__N_3613[1] ), .I3(r_SM_Main[1]), .O(n21286));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7899_3_lut_4_lut.LUT_INIT = 16'hc0aa;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (CLK_c, n29246, r_Rx_Data, r_SM_Main, GND_net, RX_N_10, 
            \r_Bit_Index[0] , n44059, \r_SM_Main_2__N_3542[2] , n27976, 
            n4, n29679, rx_data, n29672, n43733, rx_data_ready, 
            n29650, n29649, n29648, n29647, n29646, n29645, n29644, 
            n44138, VCC_net, n4_adj_4, n4_adj_5, n27971, n35414) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output n29246;
    output r_Rx_Data;
    output [2:0]r_SM_Main;
    input GND_net;
    input RX_N_10;
    output \r_Bit_Index[0] ;
    output n44059;
    output \r_SM_Main_2__N_3542[2] ;
    output n27976;
    output n4;
    input n29679;
    output [7:0]rx_data;
    input n29672;
    input n43733;
    output rx_data_ready;
    input n29650;
    input n29649;
    input n29648;
    input n29647;
    input n29646;
    input n29645;
    input n29644;
    input n44138;
    input VCC_net;
    output n4_adj_4;
    output n4_adj_5;
    output n27971;
    output n35414;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n37;
    
    wire n29315;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n29526;
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n29494;
    wire [2:0]r_SM_Main_2__N_3548;
    
    wire n1, n36093, n3, r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_3545;
    
    wire n36195, n9, n27831, n6, n49716, n49714, n6_adj_4207, 
        n27846, n40515, n40514, n40513, n40512, n40511, n40510, 
        n40509, n49667;
    
    SB_DFFESR r_Clock_Count_2063__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n29315), 
            .D(n37[7]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n29315), 
            .D(n37[6]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n29315), 
            .D(n37[5]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n29315), 
            .D(n37[4]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n29315), 
            .D(n37[3]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n29315), 
            .D(n37[2]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n29315), 
            .D(n37[1]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2063__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n29315), 
            .D(n37[0]), .R(n29526));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n29246), 
            .D(n326[1]), .R(n29494));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n29246), 
            .D(n326[2]), .R(n29494));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n36093), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i2178_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2178_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n44059));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i22582_2_lut (.I0(n44059), .I1(\r_SM_Main_2__N_3542[2] ), .I2(GND_net), 
            .I3(GND_net), .O(r_SM_Main_2__N_3545[0]));
    defparam i22582_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2171_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2171_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n36195), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i4_4_lut (.I0(n9), .I1(n27831), .I2(r_Clock_Count[3]), .I3(r_Clock_Count[1]), 
            .O(r_SM_Main_2__N_3548[0]));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22565_4_lut (.I0(r_Clock_Count[0]), .I1(n27831), .I2(n6), 
            .I3(r_Clock_Count[1]), .O(\r_SM_Main_2__N_3542[2] ));
    defparam i22565_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i3_2_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(GND_net), .O(n9));
    defparam i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[5]), .O(n27831));   // verilog/uart_rx.v(118[17:47])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34386_4_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[1]), .I2(n27831), 
            .I3(r_Clock_Count[3]), .O(n49716));
    defparam i34386_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i34477_3_lut (.I0(n49716), .I1(r_SM_Main[0]), .I2(n9), .I3(GND_net), 
            .O(n49714));
    defparam i34477_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n49714), .I2(\r_SM_Main_2__N_3542[2] ), 
            .I3(r_SM_Main[1]), .O(n29526));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_2_lut_adj_865 (.I0(r_SM_Main_2__N_3548[0]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4207));
    defparam i2_2_lut_adj_865.LUT_INIT = 16'h4444;
    SB_LUT4 i35191_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4207), 
            .I3(r_Rx_Data), .O(n29315));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i35191_4_lut.LUT_INIT = 16'h4555;
    SB_LUT4 i3_4_lut_adj_866 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3542[2] ), .O(n27846));
    defparam i3_4_lut_adj_866.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(n27846), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27976));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_312_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_312_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n29679));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n29672));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n43733));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n29650));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n29649));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n29648));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n29647));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n29646));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n29645));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n29644));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n44138));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_2063_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n40515), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2063_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n40514), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_8 (.CI(n40514), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n40515));
    SB_LUT4 r_Clock_Count_2063_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n40513), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_7 (.CI(n40513), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n40514));
    SB_LUT4 r_Clock_Count_2063_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n40512), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_6 (.CI(n40512), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n40513));
    SB_LUT4 r_Clock_Count_2063_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n40511), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_5 (.CI(n40511), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n40512));
    SB_LUT4 r_Clock_Count_2063_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n40510), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_4 (.CI(n40510), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n40511));
    SB_LUT4 r_Clock_Count_2063_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n40509), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_3 (.CI(n40509), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n40510));
    SB_LUT4 r_Clock_Count_2063_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2063_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2063_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n40509));
    SB_LUT4 equal_310_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_310_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_308_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5));   // verilog/uart_rx.v(97[17:39])
    defparam equal_308_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_867 (.I0(n27846), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n27971));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_867.LUT_INIT = 16'hbbbb;
    SB_LUT4 i21904_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35414));
    defparam i21904_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3545[0]), .O(n29494));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_868 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3542[2] ), .O(n29246));
    defparam i1_3_lut_4_lut_adj_868.LUT_INIT = 16'h1101;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_3_lut (.I0(n44059), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n36093));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i34446_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n49667));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34446_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n49667), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n36195));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, enable_slow_N_4190, \state[1] , CLK_c, \state[0] , 
            \state[3] , \state[0]_adj_2 , read, n5740, \state[2] , 
            n29661, rw, n43841, data_ready, n6387, sda_enable, \state_7__N_4087[0] , 
            \saved_addr[0] , \state_7__N_4103[3] , n6935, scl_enable, 
            n10, n35178, n35422, n8, VCC_net, n29675, data, n4, 
            n4_adj_3, scl, sda_out, n30212, n29664, n29663, n29631, 
            n29630, n29629, n29628, n29627, n49702, n27984, n28004) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    output enable_slow_N_4190;
    output \state[1] ;
    input CLK_c;
    output \state[0] ;
    output \state[3] ;
    output \state[0]_adj_2 ;
    input read;
    output [0:0]n5740;
    output \state[2] ;
    input n29661;
    output rw;
    input n43841;
    output data_ready;
    output n6387;
    output sda_enable;
    output \state_7__N_4087[0] ;
    output \saved_addr[0] ;
    input \state_7__N_4103[3] ;
    input n6935;
    output scl_enable;
    output n10;
    output n35178;
    output n35422;
    input n8;
    input VCC_net;
    input n29675;
    output [7:0]data;
    output n4;
    output n4_adj_3;
    output scl;
    output sda_out;
    input n30212;
    input n29664;
    input n29663;
    input n29631;
    input n29630;
    input n29629;
    input n29628;
    input n29627;
    output n49702;
    output n27984;
    output n28004;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3989;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    wire [15:0]n4132;
    
    wire n39234, n41199, n15, n49698, n29288, n29509, n7, n27844, 
        n46909, n13, n43709, enable;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n43707, n28, n26, n27, n25, n39248, n39247, n39246, 
        n39245, n39244, n39243, n39242, n39241, n39240, n39239, 
        n39238, n39237, n39236, n39235;
    
    SB_LUT4 add_908_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4132[14]), 
            .I3(GND_net), .O(delay_counter_15__N_3989[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4132[14]), 
            .CO(n39234));
    SB_LUT4 i34385_4_lut (.I0(n41199), .I1(enable_slow_N_4190), .I2(\state[1] ), 
            .I3(n15), .O(n49698));   // verilog/eeprom.v(23[11:16])
    defparam i34385_4_lut.LUT_INIT = 16'hfaee;
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[1]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[2]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[3]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[4]), .S(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[5]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[6]), .S(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[7]), .S(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[8]), .S(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[9]), .S(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[10]), .S(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[11]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[12]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[13]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[14]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[15]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 state_7__I_0_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/eeprom.v(51[5:9])
    defparam state_7__I_0_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut (.I0(n7), .I1(\state[3] ), .I2(\state[0]_adj_2 ), 
            .I3(n27844), .O(n41199));   // verilog/eeprom.v(42[12:28])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(n15), .I1(n46909), .I2(enable_slow_N_4190), 
            .I3(n13), .O(n43709));   // verilog/coms.v(145[4] 299[11])
    defparam i1_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 mux_1366_Mux_0_i1_4_lut (.I0(read), .I1(n27844), .I2(\state[0] ), 
            .I3(enable_slow_N_4190), .O(n5740[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_1366_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n5740[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n29288), 
            .D(delay_counter_15__N_3989[0]), .R(n29509));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i15995_2_lut (.I0(n29288), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n29509));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15995_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n29288));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n43709));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n43707));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n29661));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n43841));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_908_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4132[14]), 
            .I3(n39248), .O(delay_counter_15__N_3989[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_908_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4132[14]), 
            .I3(n39247), .O(delay_counter_15__N_3989[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_16 (.CI(n39247), .I0(delay_counter[14]), .I1(n4132[14]), 
            .CO(n39248));
    SB_LUT4 add_908_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4132[14]), 
            .I3(n39246), .O(delay_counter_15__N_3989[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_15 (.CI(n39246), .I0(delay_counter[13]), .I1(n4132[14]), 
            .CO(n39247));
    SB_LUT4 add_908_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4132[14]), 
            .I3(n39245), .O(delay_counter_15__N_3989[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_14 (.CI(n39245), .I0(delay_counter[12]), .I1(n4132[14]), 
            .CO(n39246));
    SB_LUT4 add_908_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4132[14]), 
            .I3(n39244), .O(delay_counter_15__N_3989[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_13 (.CI(n39244), .I0(delay_counter[11]), .I1(n4132[14]), 
            .CO(n39245));
    SB_LUT4 add_908_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4132[14]), 
            .I3(n39243), .O(delay_counter_15__N_3989[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_12 (.CI(n39243), .I0(delay_counter[10]), .I1(n4132[14]), 
            .CO(n39244));
    SB_LUT4 add_908_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4132[14]), 
            .I3(n39242), .O(delay_counter_15__N_3989[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_11 (.CI(n39242), .I0(delay_counter[9]), .I1(n4132[14]), 
            .CO(n39243));
    SB_LUT4 add_908_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4132[14]), 
            .I3(n39241), .O(delay_counter_15__N_3989[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_10 (.CI(n39241), .I0(delay_counter[8]), .I1(n4132[14]), 
            .CO(n39242));
    SB_LUT4 add_908_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4132[14]), 
            .I3(n39240), .O(delay_counter_15__N_3989[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_9 (.CI(n39240), .I0(delay_counter[7]), .I1(n4132[14]), 
            .CO(n39241));
    SB_LUT4 add_908_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4132[14]), 
            .I3(n39239), .O(delay_counter_15__N_3989[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_8 (.CI(n39239), .I0(delay_counter[6]), .I1(n4132[14]), 
            .CO(n39240));
    SB_LUT4 add_908_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4132[14]), 
            .I3(n39238), .O(delay_counter_15__N_3989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_7 (.CI(n39238), .I0(delay_counter[5]), .I1(n4132[14]), 
            .CO(n39239));
    SB_LUT4 add_908_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4132[14]), 
            .I3(n39237), .O(delay_counter_15__N_3989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_6 (.CI(n39237), .I0(delay_counter[4]), .I1(n4132[14]), 
            .CO(n39238));
    SB_LUT4 add_908_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4132[14]), 
            .I3(n39236), .O(delay_counter_15__N_3989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_5 (.CI(n39236), .I0(delay_counter[3]), .I1(n4132[14]), 
            .CO(n39237));
    SB_LUT4 add_908_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4132[14]), 
            .I3(n39235), .O(delay_counter_15__N_3989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_4 (.CI(n39235), .I0(delay_counter[2]), .I1(n4132[14]), 
            .CO(n39236));
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n27844));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35229_2_lut (.I0(n27844), .I1(enable_slow_N_4190), .I2(GND_net), 
            .I3(GND_net), .O(n4132[14]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i35229_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_908_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4132[14]), 
            .I3(n39234), .O(delay_counter_15__N_3989[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_908_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_908_3 (.CI(n39234), .I0(delay_counter[1]), .I1(n4132[14]), 
            .CO(n39235));
    SB_LUT4 i24_4_lut_4_lut (.I0(\state[1] ), .I1(read), .I2(\state[0] ), 
            .I3(n49698), .O(n43707));   // verilog/eeprom.v(23[11:16])
    defparam i24_4_lut_4_lut.LUT_INIT = 16'hf404;
    SB_LUT4 i2_4_lut_4_lut (.I0(n41199), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n46909));   // verilog/coms.v(145[4] 299[11])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[1] ), .I1(enable_slow_N_4190), .I2(read), 
            .I3(\state[0] ), .O(n13));   // verilog/coms.v(145[4] 299[11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'haa8a;
    i2c_controller i2c (.CLK_c(CLK_c), .n6387(n6387), .\state[1] (state[1]), 
            .\state[2] (\state[2] ), .\state[3] (\state[3] ), .sda_enable(sda_enable), 
            .\state_7__N_4087[0] (\state_7__N_4087[0] ), .enable_slow_N_4190(enable_slow_N_4190), 
            .GND_net(GND_net), .\saved_addr[0] (\saved_addr[0] ), .\state[0] (\state[0]_adj_2 ), 
            .\state_7__N_4103[3] (\state_7__N_4103[3] ), .n6935(n6935), 
            .scl_enable(scl_enable), .enable(enable), .n10(n10), .n35178(n35178), 
            .n35422(n35422), .n8(n8), .VCC_net(VCC_net), .n29675(n29675), 
            .data({data}), .n4(n4), .n4_adj_1(n4_adj_3), .scl(scl), 
            .sda_out(sda_out), .n30212(n30212), .n29664(n29664), .n29663(n29663), 
            .n29631(n29631), .n29630(n29630), .n29629(n29629), .n29628(n29628), 
            .n29627(n29627), .n49702(n49702), .n27984(n27984), .n28004(n28004)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (CLK_c, n6387, \state[1] , \state[2] , \state[3] , 
            sda_enable, \state_7__N_4087[0] , enable_slow_N_4190, GND_net, 
            \saved_addr[0] , \state[0] , \state_7__N_4103[3] , n6935, 
            scl_enable, enable, n10, n35178, n35422, n8, VCC_net, 
            n29675, data, n4, n4_adj_1, scl, sda_out, n30212, 
            n29664, n29663, n29631, n29630, n29629, n29628, n29627, 
            n49702, n27984, n28004) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    output n6387;
    output \state[1] ;
    output \state[2] ;
    output \state[3] ;
    output sda_enable;
    output \state_7__N_4087[0] ;
    output enable_slow_N_4190;
    input GND_net;
    output \saved_addr[0] ;
    output \state[0] ;
    input \state_7__N_4103[3] ;
    input n6935;
    output scl_enable;
    input enable;
    output n10;
    output n35178;
    output n35422;
    input n8;
    input VCC_net;
    input n29675;
    output [7:0]data;
    output n4;
    output n4_adj_1;
    output scl;
    output sda_out;
    input n30212;
    input n29664;
    input n29663;
    input n29631;
    input n29630;
    input n29629;
    input n29628;
    input n29627;
    output n49702;
    output n27984;
    output n28004;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n29529, n5, n36107, n35511, n36105, n43891, n46742, n20075, 
        n6809, n29486, enable_slow_N_4189, i2c_clk_N_4176;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n49675, n49630, n6058;
    wire [0:0]n6094;
    
    wire n15, n44967, n6380, n37, n29358;
    wire [7:0]n119;
    
    wire n29571, n43781, sda_out_adj_4194, scl_enable_N_4177, n33, 
        n34, n39, n29238, n7, n10_c, n10_adj_4195, n49731, n11, 
        n12, n9, state_7__N_4086, n11_adj_4197, n11_adj_4198, n10_adj_4199, 
        n39424, n39423, n39422, n39421, n39420, n39419, n39418, 
        n11_adj_4203, n40559, n40558, n40557, n40556, n40555;
    
    SB_DFFSR counter2_2067_2068__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n29529));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6387), .D(n5), 
            .S(n36107));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6387), .D(n35511), 
            .S(n36105));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6387), .D(n43891), 
            .S(n46742));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n6809), 
            .D(n20075), .S(n29486));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_LUT4 i35212_2_lut (.I0(\state_7__N_4087[0] ), .I1(enable_slow_N_4190), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4189));   // verilog/i2c_controller.v(62[6:32])
    defparam i35212_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n29529), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4176));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34339_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n49675));   // verilog/i2c_controller.v(198[28:35])
    defparam i34339_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i34380_4_lut (.I0(n49675), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n49630));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i34380_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 mux_1503_i1_4_lut (.I0(n49630), .I1(\state[0] ), .I2(n6058), 
            .I3(\state[2] ), .O(n6094[0]));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam mux_1503_i1_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i29611_2_lut (.I0(\state_7__N_4103[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n44967));
    defparam i29611_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n6380), .I1(n44967), .I2(n6935), .I3(n37), 
            .O(n29358));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n29358), .D(n119[6]), 
            .R(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n29358), .D(n119[5]), 
            .R(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4194), .C(i2c_clk), .E(n43781), 
            .D(n6094[0]));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n29358), .D(n119[0]), 
            .S(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n29358), .D(n119[4]), 
            .R(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4176));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4177));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n29486));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_860 (.I0(n34), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i1_2_lut_adj_860.LUT_INIT = 16'heeee;
    SB_LUT4 i35240_4_lut (.I0(n6058), .I1(n39), .I2(\state[2] ), .I3(\state[1] ), 
            .O(n6809));
    defparam i35240_4_lut.LUT_INIT = 16'hc8cc;
    SB_LUT4 i35205_2_lut (.I0(\state[0] ), .I1(n6058), .I2(GND_net), .I3(GND_net), 
            .O(n20075));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i35205_2_lut.LUT_INIT = 16'h4444;
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4087[0] ), .C(CLK_c), .E(n29238), 
            .D(enable_slow_N_4189));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n29358), .D(n119[3]), 
            .R(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_adj_861 (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_861.LUT_INIT = 16'h4444;
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n29358), .D(n119[2]), 
            .S(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i34433_4_lut (.I0(n10_c), .I1(n10_adj_4195), .I2(\state_7__N_4103[3] ), 
            .I3(enable), .O(n49731));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i34433_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n7), .I2(n49731), .I3(\state[0] ), 
            .O(n43891));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i35304_2_lut (.I0(\state_7__N_4103[3] ), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n35511));
    defparam i35304_2_lut.LUT_INIT = 16'h1111;
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n29358), .D(n119[1]), 
            .S(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4195));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6380));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i35200_4_lut (.I0(state_7__N_4086), .I1(n6380), .I2(n11_adj_4197), 
            .I3(n35178), .O(n6387));
    defparam i35200_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut_adj_862 (.I0(n11_adj_4198), .I1(n11), .I2(\state_7__N_4103[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_862.LUT_INIT = 16'h5755;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4199));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4199), .I2(counter2[0]), 
            .I3(GND_net), .O(n29529));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i21912_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35422));
    defparam i21912_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n29675));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_316_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_316_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_318_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_318_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i21769_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i21769_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2367_2_lut (.I0(sda_out_adj_4194), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_259_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_c));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_259_i10_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n30212));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n39424), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n39423), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n39423), .I0(counter[6]), .I1(VCC_net), 
            .CO(n39424));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n39422), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n39422), .I0(counter[5]), .I1(VCC_net), 
            .CO(n39423));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n39421), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n39421), .I0(counter[4]), .I1(VCC_net), 
            .CO(n39422));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n39420), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n39420), .I0(counter[3]), .I1(VCC_net), 
            .CO(n39421));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n39419), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n39419), .I0(counter[2]), .I1(VCC_net), 
            .CO(n39420));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n39418), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n39418), .I0(counter[1]), .I1(VCC_net), 
            .CO(n39419));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n39418));
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n29664));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n29663));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n29631));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n29630));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n29629));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n29628));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n29627));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2067_2068__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n29529));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n29529));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n29529));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n29529));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2067_2068__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n29529));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i34381_3_lut_4_lut (.I0(n11_adj_4197), .I1(n11_adj_4203), .I2(enable_slow_N_4190), 
            .I3(\state_7__N_4087[0] ), .O(n49702));
    defparam i34381_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 counter2_2067_2068_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n40559), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2067_2068_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n40558), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_6 (.CI(n40558), .I0(GND_net), .I1(counter2[4]), 
            .CO(n40559));
    SB_LUT4 counter2_2067_2068_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n40557), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_5 (.CI(n40557), .I0(GND_net), .I1(counter2[3]), 
            .CO(n40558));
    SB_LUT4 counter2_2067_2068_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n40556), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_4 (.CI(n40556), .I0(GND_net), .I1(counter2[2]), 
            .CO(n40557));
    SB_LUT4 counter2_2067_2068_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n40555), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_3 (.CI(n40555), .I0(GND_net), .I1(counter2[1]), 
            .CO(n40556));
    SB_LUT4 counter2_2067_2068_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2067_2068_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2067_2068_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n40555));
    SB_LUT4 i35252_3_lut_4_lut (.I0(n11_adj_4197), .I1(n11_adj_4203), .I2(n15), 
            .I3(n6387), .O(n36107));
    defparam i35252_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4203));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n29358), .D(n119[7]), 
            .R(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i22507_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_4086));
    defparam i22507_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i35250_3_lut_4_lut (.I0(n9), .I1(n10_adj_4195), .I2(n11_adj_4203), 
            .I3(n6387), .O(n36105));   // verilog/i2c_controller.v(151[5:14])
    defparam i35250_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10_adj_4195), .I2(counter[0]), 
            .I3(GND_net), .O(n27984));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_863 (.I0(n9), .I1(n10_adj_4195), .I2(counter[0]), 
            .I3(GND_net), .O(n28004));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_863.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 i22527_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4177));
    defparam i22527_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(\state[2] ), .O(n6058));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h001c;
    SB_LUT4 equal_2051_i19_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4190));
    defparam equal_2051_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4198));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 equal_259_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_259_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4197));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i22479_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n35178));
    defparam i22479_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i35248_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6387), .O(n46742));
    defparam i35248_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 i29560_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n44967), .O(n29571));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i29560_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_3_lut_adj_864 (.I0(enable), .I1(\state_7__N_4087[0] ), 
            .I2(enable_slow_N_4190), .I3(GND_net), .O(n29238));
    defparam i1_2_lut_3_lut_adj_864.LUT_INIT = 16'heaea;
    SB_LUT4 i35238_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n43781));
    defparam i35238_4_lut_4_lut.LUT_INIT = 16'h0156;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (\a_new[1] , b_prev, GND_net, ENCODER1_B_N_keep, 
            n1653, ENCODER1_A_N_keep, direction_N_3907, encoder1_position, 
            n29674, n1658, VCC_net) /* synthesis lattice_noprune=1 */ ;
    output \a_new[1] ;
    output b_prev;
    input GND_net;
    input ENCODER1_B_N_keep;
    input n1653;
    input ENCODER1_A_N_keep;
    output direction_N_3907;
    output [31:0]encoder1_position;
    input n29674;
    output n1658;
    input VCC_net;
    
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire a_prev_N_3913, direction_N_3906, debounce_cnt, n29688;
    wire [31:0]n133;
    
    wire direction_N_3910, a_prev, n29673, n40508, n40507, n40506, 
        n40505, n40504, n40503, n40502, n40501, n40500, n40499, 
        n40498, n40497, n40496, n40495, n40494, n40493, n40492, 
        n40491, n40490, n40489, n40488, n40487, n40486, n40485, 
        n40484, n40483, n40482, n40481, n40480, n40479, n40478;
    
    SB_LUT4 i35222_4_lut (.I0(a_new[0]), .I1(b_new[0]), .I2(\a_new[1] ), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i35222_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(\a_new[1] ), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1653), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new[0]), .C(n1653), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1653), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(\a_new[1] ), .C(n1653), .D(a_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1653), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1653), .D(n29688));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2061__i0 (.Q(encoder1_position[0]), .C(n1653), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(\a_new[1] ), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_DFF direction_57 (.Q(n1658), .C(n1653), .D(n29674));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1653), .D(n29673));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2061__i1 (.Q(encoder1_position[1]), .C(n1653), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i2 (.Q(encoder1_position[2]), .C(n1653), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i3 (.Q(encoder1_position[3]), .C(n1653), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i4 (.Q(encoder1_position[4]), .C(n1653), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i5 (.Q(encoder1_position[5]), .C(n1653), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i6 (.Q(encoder1_position[6]), .C(n1653), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i7 (.Q(encoder1_position[7]), .C(n1653), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i8 (.Q(encoder1_position[8]), .C(n1653), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i9 (.Q(encoder1_position[9]), .C(n1653), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i10 (.Q(encoder1_position[10]), .C(n1653), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i11 (.Q(encoder1_position[11]), .C(n1653), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i12 (.Q(encoder1_position[12]), .C(n1653), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i13 (.Q(encoder1_position[13]), .C(n1653), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i14 (.Q(encoder1_position[14]), .C(n1653), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i15 (.Q(encoder1_position[15]), .C(n1653), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i16 (.Q(encoder1_position[16]), .C(n1653), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i17 (.Q(encoder1_position[17]), .C(n1653), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i18 (.Q(encoder1_position[18]), .C(n1653), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i19 (.Q(encoder1_position[19]), .C(n1653), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i20 (.Q(encoder1_position[20]), .C(n1653), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i21 (.Q(encoder1_position[21]), .C(n1653), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i22 (.Q(encoder1_position[22]), .C(n1653), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i23 (.Q(encoder1_position[23]), .C(n1653), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i24 (.Q(encoder1_position[24]), .C(n1653), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i25 (.Q(encoder1_position[25]), .C(n1653), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i26 (.Q(encoder1_position[26]), .C(n1653), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i27 (.Q(encoder1_position[27]), .C(n1653), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i28 (.Q(encoder1_position[28]), .C(n1653), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i29 (.Q(encoder1_position[29]), .C(n1653), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i30 (.Q(encoder1_position[30]), .C(n1653), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2061__i31 (.Q(encoder1_position[31]), .C(n1653), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 i16161_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n29688));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16161_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 position_2061_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[31]), .I3(n40508), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2061_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[30]), .I3(n40507), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_32 (.CI(n40507), .I0(direction_N_3906), 
            .I1(encoder1_position[30]), .CO(n40508));
    SB_LUT4 position_2061_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[29]), .I3(n40506), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_31 (.CI(n40506), .I0(direction_N_3906), 
            .I1(encoder1_position[29]), .CO(n40507));
    SB_LUT4 position_2061_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[28]), .I3(n40505), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_30 (.CI(n40505), .I0(direction_N_3906), 
            .I1(encoder1_position[28]), .CO(n40506));
    SB_LUT4 position_2061_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[27]), .I3(n40504), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_29 (.CI(n40504), .I0(direction_N_3906), 
            .I1(encoder1_position[27]), .CO(n40505));
    SB_LUT4 position_2061_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[26]), .I3(n40503), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_28 (.CI(n40503), .I0(direction_N_3906), 
            .I1(encoder1_position[26]), .CO(n40504));
    SB_LUT4 position_2061_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[25]), .I3(n40502), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_27 (.CI(n40502), .I0(direction_N_3906), 
            .I1(encoder1_position[25]), .CO(n40503));
    SB_LUT4 position_2061_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[24]), .I3(n40501), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_26 (.CI(n40501), .I0(direction_N_3906), 
            .I1(encoder1_position[24]), .CO(n40502));
    SB_LUT4 position_2061_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[23]), .I3(n40500), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_25 (.CI(n40500), .I0(direction_N_3906), 
            .I1(encoder1_position[23]), .CO(n40501));
    SB_LUT4 position_2061_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[22]), .I3(n40499), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_24 (.CI(n40499), .I0(direction_N_3906), 
            .I1(encoder1_position[22]), .CO(n40500));
    SB_LUT4 position_2061_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[21]), .I3(n40498), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16146_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(\a_new[1] ), 
            .I3(a_prev), .O(n29673));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i16146_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY position_2061_add_4_23 (.CI(n40498), .I0(direction_N_3906), 
            .I1(encoder1_position[21]), .CO(n40499));
    SB_LUT4 position_2061_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[20]), .I3(n40497), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_22 (.CI(n40497), .I0(direction_N_3906), 
            .I1(encoder1_position[20]), .CO(n40498));
    SB_LUT4 position_2061_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[19]), .I3(n40496), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_21 (.CI(n40496), .I0(direction_N_3906), 
            .I1(encoder1_position[19]), .CO(n40497));
    SB_LUT4 position_2061_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[18]), .I3(n40495), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_20 (.CI(n40495), .I0(direction_N_3906), 
            .I1(encoder1_position[18]), .CO(n40496));
    SB_LUT4 position_2061_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[17]), .I3(n40494), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_19 (.CI(n40494), .I0(direction_N_3906), 
            .I1(encoder1_position[17]), .CO(n40495));
    SB_LUT4 position_2061_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[16]), .I3(n40493), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_18 (.CI(n40493), .I0(direction_N_3906), 
            .I1(encoder1_position[16]), .CO(n40494));
    SB_LUT4 position_2061_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[15]), .I3(n40492), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_17 (.CI(n40492), .I0(direction_N_3906), 
            .I1(encoder1_position[15]), .CO(n40493));
    SB_LUT4 position_2061_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[14]), .I3(n40491), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_16 (.CI(n40491), .I0(direction_N_3906), 
            .I1(encoder1_position[14]), .CO(n40492));
    SB_LUT4 position_2061_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[13]), .I3(n40490), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_15 (.CI(n40490), .I0(direction_N_3906), 
            .I1(encoder1_position[13]), .CO(n40491));
    SB_LUT4 position_2061_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[12]), .I3(n40489), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_14 (.CI(n40489), .I0(direction_N_3906), 
            .I1(encoder1_position[12]), .CO(n40490));
    SB_LUT4 position_2061_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[11]), .I3(n40488), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_13 (.CI(n40488), .I0(direction_N_3906), 
            .I1(encoder1_position[11]), .CO(n40489));
    SB_LUT4 position_2061_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[10]), .I3(n40487), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_12 (.CI(n40487), .I0(direction_N_3906), 
            .I1(encoder1_position[10]), .CO(n40488));
    SB_LUT4 position_2061_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[9]), .I3(n40486), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_11 (.CI(n40486), .I0(direction_N_3906), 
            .I1(encoder1_position[9]), .CO(n40487));
    SB_LUT4 position_2061_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[8]), .I3(n40485), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_10 (.CI(n40485), .I0(direction_N_3906), 
            .I1(encoder1_position[8]), .CO(n40486));
    SB_LUT4 position_2061_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[7]), .I3(n40484), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_9 (.CI(n40484), .I0(direction_N_3906), 
            .I1(encoder1_position[7]), .CO(n40485));
    SB_LUT4 position_2061_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[6]), .I3(n40483), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_8 (.CI(n40483), .I0(direction_N_3906), 
            .I1(encoder1_position[6]), .CO(n40484));
    SB_LUT4 position_2061_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[5]), .I3(n40482), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_7 (.CI(n40482), .I0(direction_N_3906), 
            .I1(encoder1_position[5]), .CO(n40483));
    SB_LUT4 position_2061_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[4]), .I3(n40481), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_6 (.CI(n40481), .I0(direction_N_3906), 
            .I1(encoder1_position[4]), .CO(n40482));
    SB_LUT4 position_2061_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[3]), .I3(n40480), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_5 (.CI(n40480), .I0(direction_N_3906), 
            .I1(encoder1_position[3]), .CO(n40481));
    SB_LUT4 position_2061_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[2]), .I3(n40479), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_4 (.CI(n40479), .I0(direction_N_3906), 
            .I1(encoder1_position[2]), .CO(n40480));
    SB_LUT4 position_2061_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[1]), .I3(n40478), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_3 (.CI(n40478), .I0(direction_N_3906), 
            .I1(encoder1_position[1]), .CO(n40479));
    SB_LUT4 position_2061_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2061_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2061_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n40478));
    
endmodule
//
// Verilog Description of module \grp_debouncer(3,1000) 
//

module \grp_debouncer(3,1000)  (reg_B, CLK_c, n29693, data_o, n29692, 
            data_i, n46952, n29624, GND_net, VCC_net);
    output [2:0]reg_B;
    input CLK_c;
    input n29693;
    output [2:0]data_o;
    input n29692;
    input [2:0]data_i;
    output n46952;
    input n29624;
    input GND_net;
    input VCC_net;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [9:0]n45;
    wire [9:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_9__N_812, n6, n40477, n40476, n40475, n40474, 
        n40473, n40472, n40471, n40470, n40469, n16, n17;
    
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(CLK_c), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(CLK_c), .D(n29693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i2 (.Q(data_o[2]), .C(CLK_c), .D(n29692));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_2060__i0 (.Q(cnt_reg[0]), .C(CLK_c), .D(n45[0]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i2 (.Q(reg_B[2]), .C(CLK_c), .D(reg_A[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(CLK_c), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(CLK_c), .D(data_i[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(CLK_c), .D(data_i[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(reg_B[1]), .I2(reg_A[0]), .I3(reg_A[1]), 
            .O(n6));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(n46952), .I1(n6), .I2(reg_B[2]), .I3(reg_A[2]), 
            .O(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i3_4_lut.LUT_INIT = 16'hdffd;
    SB_DFFSR cnt_reg_2060__i1 (.Q(cnt_reg[1]), .C(CLK_c), .D(n45[1]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i2 (.Q(cnt_reg[2]), .C(CLK_c), .D(n45[2]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i3 (.Q(cnt_reg[3]), .C(CLK_c), .D(n45[3]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i4 (.Q(cnt_reg[4]), .C(CLK_c), .D(n45[4]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i5 (.Q(cnt_reg[5]), .C(CLK_c), .D(n45[5]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i6 (.Q(cnt_reg[6]), .C(CLK_c), .D(n45[6]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i7 (.Q(cnt_reg[7]), .C(CLK_c), .D(n45[7]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i8 (.Q(cnt_reg[8]), .C(CLK_c), .D(n45[8]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2060__i9 (.Q(cnt_reg[9]), .C(CLK_c), .D(n45[9]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(CLK_c), .D(n29624));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i2 (.Q(reg_A[2]), .C(CLK_c), .D(data_i[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_2060_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[9]), 
            .I3(n40477), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_2060_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[8]), 
            .I3(n40476), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_10 (.CI(n40476), .I0(GND_net), .I1(cnt_reg[8]), 
            .CO(n40477));
    SB_LUT4 cnt_reg_2060_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[7]), 
            .I3(n40475), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_9 (.CI(n40475), .I0(GND_net), .I1(cnt_reg[7]), 
            .CO(n40476));
    SB_LUT4 cnt_reg_2060_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n40474), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_8 (.CI(n40474), .I0(GND_net), .I1(cnt_reg[6]), 
            .CO(n40475));
    SB_LUT4 cnt_reg_2060_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n40473), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_7 (.CI(n40473), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n40474));
    SB_LUT4 cnt_reg_2060_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n40472), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_6 (.CI(n40472), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n40473));
    SB_LUT4 cnt_reg_2060_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n40471), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_5 (.CI(n40471), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n40472));
    SB_LUT4 cnt_reg_2060_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n40470), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_4 (.CI(n40470), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n40471));
    SB_LUT4 cnt_reg_2060_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n40469), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_3 (.CI(n40469), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n40470));
    SB_LUT4 cnt_reg_2060_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2060_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2060_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n40469));
    SB_LUT4 i6_4_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[7]), 
            .I3(cnt_reg[2]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut (.I0(cnt_reg[4]), .I1(cnt_reg[9]), .I2(cnt_reg[8]), 
            .I3(cnt_reg[5]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(cnt_reg[6]), .I2(n16), .I3(cnt_reg[3]), 
            .O(n46952));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (GND_net, pwm_out, clk32MHz, VCC_net, pwm_setpoint) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output pwm_out;
    input clk32MHz;
    input VCC_net;
    input [23:0]pwm_setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n40448;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n40449, pwm_out_N_797;
    wire [23:0]n101;
    
    wire n40447, n40446, pwm_counter_23__N_795, n46515, n22, n15, 
        n20, n24, n19, n41, n39, n45, n43, n37, n29, n31, 
        n23, n25, n35, n33, n11, n13, n15_adj_4191, n27, n9, 
        n17, n19_adj_4192, n21, n49877, n49826, n12, n30, n49888, 
        n50160, n50156, n50505, n50325, n50541, n6, n50405, n50406, 
        n16, n24_adj_4193, n49797, n8, n49790, n50411, n50115, 
        n4, n50489, n50490, n49815, n10, n49812, n50556, n50408, 
        n50602, n50603, n50583, n49800, n50495, n40, n50497, n40468, 
        n40467, n40466, n40465, n40464, n40463, n40462, n40461, 
        n40460, n40459, n40458, n40457, n40456, n40455, n40454, 
        n40453, n40452, n40451, n40450;
    
    SB_CARRY pwm_counter_2059_add_4_5 (.CI(n40448), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n40449));
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_797));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_2059_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n40447), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_4 (.CI(n40447), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n40448));
    SB_LUT4 pwm_counter_2059_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n40446), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_3 (.CI(n40446), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n40447));
    SB_LUT4 pwm_counter_2059_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n40446));
    SB_DFFSR pwm_counter_2059__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n46515));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i9_4_lut (.I0(pwm_counter[18]), .I1(pwm_counter[20]), .I2(pwm_counter[15]), 
            .I3(pwm_counter[16]), .O(n22));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n46515), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n15));
    defparam i2_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[17]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15), .I1(n22), .I2(pwm_counter[12]), .I3(pwm_counter[22]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[19]), .I1(pwm_counter[14]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i35913_4_lut (.I0(pwm_counter[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(pwm_counter_23__N_795));   // verilog/pwm.v(18[8:40])
    defparam i35913_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4191));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4192));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34440_4_lut (.I0(n21), .I1(n19_adj_4192), .I2(n17), .I3(n9), 
            .O(n49877));
    defparam i34440_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34389_4_lut (.I0(n27), .I1(n15_adj_4191), .I2(n13), .I3(n11), 
            .O(n49826));
    defparam i34389_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34723_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n49888), 
            .O(n50160));
    defparam i34723_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34719_4_lut (.I0(n19_adj_4192), .I1(n17), .I2(n15_adj_4191), 
            .I3(n50160), .O(n50156));
    defparam i34719_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35067_4_lut (.I0(n25), .I1(n23), .I2(n21), .I3(n50156), 
            .O(n50505));
    defparam i35067_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34887_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n50505), 
            .O(n50325));
    defparam i34887_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35103_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n50325), 
            .O(n50541));
    defparam i35103_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34967_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21), .I3(GND_net), 
            .O(n50405));   // verilog/pwm.v(21[8:24])
    defparam i34967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34968_3_lut (.I0(n50405), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n50406));   // verilog/pwm.v(21[8:24])
    defparam i34968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4193));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34360_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n49877), 
            .O(n49797));
    defparam i34360_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34973_4_lut (.I0(n24_adj_4193), .I1(n8), .I2(n45), .I3(n49790), 
            .O(n50411));   // verilog/pwm.v(21[8:24])
    defparam i34973_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34678_3_lut (.I0(n50406), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n50115));   // verilog/pwm.v(21[8:24])
    defparam i34678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i35051_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n50489));   // verilog/pwm.v(21[8:24])
    defparam i35051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35052_3_lut (.I0(n50489), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n50490));   // verilog/pwm.v(21[8:24])
    defparam i35052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34378_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n49826), 
            .O(n49815));
    defparam i34378_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35118_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n49812), 
            .O(n50556));   // verilog/pwm.v(21[8:24])
    defparam i35118_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34970_3_lut (.I0(n50490), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n50408));   // verilog/pwm.v(21[8:24])
    defparam i34970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35164_4_lut (.I0(n50408), .I1(n50556), .I2(n35), .I3(n49815), 
            .O(n50602));   // verilog/pwm.v(21[8:24])
    defparam i35164_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35165_3_lut (.I0(n50602), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n50603));   // verilog/pwm.v(21[8:24])
    defparam i35165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35145_3_lut (.I0(n50603), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n50583));   // verilog/pwm.v(21[8:24])
    defparam i35145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34363_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n50541), 
            .O(n49800));
    defparam i34363_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35057_4_lut (.I0(n50115), .I1(n50411), .I2(n45), .I3(n49797), 
            .O(n50495));   // verilog/pwm.v(21[8:24])
    defparam i35057_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35135_3_lut (.I0(n50583), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n40));   // verilog/pwm.v(21[8:24])
    defparam i35135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35059_4_lut (.I0(n40), .I1(n50495), .I2(n45), .I3(n49800), 
            .O(n50497));   // verilog/pwm.v(21[8:24])
    defparam i35059_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35060_3_lut (.I0(n50497), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_797));   // verilog/pwm.v(21[8:24])
    defparam i35060_3_lut.LUT_INIT = 16'h8e8e;
    SB_DFFSR pwm_counter_2059__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2059__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_2059_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n40468), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2059_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n40467), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_24 (.CI(n40467), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n40468));
    SB_LUT4 pwm_counter_2059_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n40466), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_23 (.CI(n40466), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n40467));
    SB_LUT4 pwm_counter_2059_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n40465), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_22 (.CI(n40465), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n40466));
    SB_LUT4 pwm_counter_2059_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n40464), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_21 (.CI(n40464), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n40465));
    SB_LUT4 pwm_counter_2059_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n40463), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_20 (.CI(n40463), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n40464));
    SB_LUT4 pwm_counter_2059_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n40462), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_19 (.CI(n40462), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n40463));
    SB_LUT4 pwm_counter_2059_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n40461), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_18 (.CI(n40461), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n40462));
    SB_LUT4 pwm_counter_2059_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n40460), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_17 (.CI(n40460), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n40461));
    SB_LUT4 pwm_counter_2059_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n40459), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_16 (.CI(n40459), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n40460));
    SB_LUT4 pwm_counter_2059_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n40458), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_15 (.CI(n40458), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n40459));
    SB_LUT4 pwm_counter_2059_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n40457), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_14 (.CI(n40457), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n40458));
    SB_LUT4 pwm_counter_2059_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n40456), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_13 (.CI(n40456), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n40457));
    SB_LUT4 pwm_counter_2059_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n40455), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_12 (.CI(n40455), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n40456));
    SB_LUT4 pwm_counter_2059_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n40454), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_11 (.CI(n40454), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n40455));
    SB_LUT4 pwm_counter_2059_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n40453), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_10 (.CI(n40453), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n40454));
    SB_LUT4 pwm_counter_2059_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n40452), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_9 (.CI(n40452), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n40453));
    SB_LUT4 pwm_counter_2059_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n40451), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_8 (.CI(n40451), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n40452));
    SB_LUT4 pwm_counter_2059_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n40450), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_7 (.CI(n40450), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n40451));
    SB_LUT4 pwm_counter_2059_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n40449), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2059_add_4_6 (.CI(n40449), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n40450));
    SB_LUT4 pwm_counter_2059_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n40448), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2059_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34451_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n49888));   // verilog/pwm.v(21[8:24])
    defparam i34451_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34353_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n49790));
    defparam i34353_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34375_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n49812));
    defparam i34375_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
