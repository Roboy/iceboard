-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 12 2017 08:26:01

-- File Generated:     Jan 29 2020 18:32:34

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TinyFPGA_B" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TinyFPGA_B
entity TinyFPGA_B is
port (
    USBPU : out std_logic;
    TX : out std_logic;
    SDA : inout std_logic;
    SCL : inout std_logic;
    RX : in std_logic;
    NEOPXL : out std_logic;
    LED : out std_logic;
    INLC : out std_logic;
    INLB : out std_logic;
    INLA : out std_logic;
    INHC : out std_logic;
    INHB : out std_logic;
    INHA : out std_logic;
    HALL3 : in std_logic;
    HALL2 : in std_logic;
    HALL1 : in std_logic;
    FAULT_N : in std_logic;
    ENCODER1_B : in std_logic;
    ENCODER1_A : in std_logic;
    ENCODER0_B : in std_logic;
    ENCODER0_A : in std_logic;
    DE : out std_logic;
    CS_MISO : in std_logic;
    CS_CLK : out std_logic;
    CS : out std_logic;
    CLK : in std_logic);
end TinyFPGA_B;

-- Architecture of TinyFPGA_B
-- View name is \INTERFACE\
architecture \INTERFACE\ of TinyFPGA_B is

signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30136\ : std_logic;
signal \N__30129\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30127\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30102\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30091\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30073\ : std_logic;
signal \N__30066\ : std_logic;
signal \N__30065\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30056\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30047\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30037\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30028\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30011\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30002\ : std_logic;
signal \N__30001\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29980\ : std_logic;
signal \N__29977\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29945\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29926\ : std_logic;
signal \N__29923\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29915\ : std_logic;
signal \N__29912\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29897\ : std_logic;
signal \N__29896\ : std_logic;
signal \N__29893\ : std_logic;
signal \N__29890\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29878\ : std_logic;
signal \N__29875\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29867\ : std_logic;
signal \N__29866\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29821\ : std_logic;
signal \N__29818\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29813\ : std_logic;
signal \N__29810\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29798\ : std_logic;
signal \N__29797\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29756\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29750\ : std_logic;
signal \N__29747\ : std_logic;
signal \N__29744\ : std_logic;
signal \N__29741\ : std_logic;
signal \N__29738\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29695\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29687\ : std_logic;
signal \N__29684\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29657\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29633\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29603\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29578\ : std_logic;
signal \N__29575\ : std_logic;
signal \N__29572\ : std_logic;
signal \N__29569\ : std_logic;
signal \N__29566\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29507\ : std_logic;
signal \N__29504\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29500\ : std_logic;
signal \N__29497\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29491\ : std_logic;
signal \N__29488\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29458\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29419\ : std_logic;
signal \N__29414\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29395\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29287\ : std_logic;
signal \N__29284\ : std_logic;
signal \N__29281\ : std_logic;
signal \N__29276\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29269\ : std_logic;
signal \N__29266\ : std_logic;
signal \N__29263\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29252\ : std_logic;
signal \N__29251\ : std_logic;
signal \N__29248\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29211\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29208\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29205\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29198\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29185\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29181\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29176\ : std_logic;
signal \N__29175\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29173\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29171\ : std_logic;
signal \N__29170\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29165\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29144\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29112\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29098\ : std_logic;
signal \N__29097\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29094\ : std_logic;
signal \N__29091\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29084\ : std_logic;
signal \N__29081\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29044\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29025\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29001\ : std_logic;
signal \N__28998\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28971\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28928\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28925\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28921\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28915\ : std_logic;
signal \N__28912\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28901\ : std_logic;
signal \N__28898\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28896\ : std_logic;
signal \N__28893\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28885\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28882\ : std_logic;
signal \N__28879\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28824\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28778\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28771\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28766\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28763\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28717\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28714\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28690\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28651\ : std_logic;
signal \N__28648\ : std_logic;
signal \N__28645\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28625\ : std_logic;
signal \N__28616\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28576\ : std_logic;
signal \N__28573\ : std_logic;
signal \N__28570\ : std_logic;
signal \N__28567\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28561\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28557\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28544\ : std_logic;
signal \N__28543\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28538\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28480\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28460\ : std_logic;
signal \N__28451\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28441\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28433\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28412\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28379\ : std_logic;
signal \N__28376\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28306\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28298\ : std_logic;
signal \N__28295\ : std_logic;
signal \N__28292\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28289\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28247\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28204\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28153\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28129\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28063\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28033\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__28003\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27988\ : std_logic;
signal \N__27985\ : std_logic;
signal \N__27970\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27957\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27899\ : std_logic;
signal \N__27896\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27843\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27793\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27749\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27741\ : std_logic;
signal \N__27738\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27713\ : std_logic;
signal \N__27710\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27656\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27648\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27614\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27607\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27594\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27515\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27503\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27494\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27485\ : std_logic;
signal \N__27482\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27443\ : std_logic;
signal \N__27440\ : std_logic;
signal \N__27437\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27419\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27401\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27326\ : std_logic;
signal \N__27311\ : std_logic;
signal \N__27308\ : std_logic;
signal \N__27305\ : std_logic;
signal \N__27302\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27298\ : std_logic;
signal \N__27295\ : std_logic;
signal \N__27290\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27269\ : std_logic;
signal \N__27268\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27242\ : std_logic;
signal \N__27239\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27233\ : std_logic;
signal \N__27230\ : std_logic;
signal \N__27227\ : std_logic;
signal \N__27224\ : std_logic;
signal \N__27221\ : std_logic;
signal \N__27218\ : std_logic;
signal \N__27215\ : std_logic;
signal \N__27212\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27191\ : std_logic;
signal \N__27188\ : std_logic;
signal \N__27185\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27179\ : std_logic;
signal \N__27176\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27171\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27152\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27129\ : std_logic;
signal \N__27126\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27112\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__26993\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26987\ : std_logic;
signal \N__26986\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26979\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26968\ : std_logic;
signal \N__26965\ : std_logic;
signal \N__26962\ : std_logic;
signal \N__26951\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26897\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26886\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26877\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26828\ : std_logic;
signal \N__26825\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26819\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26816\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26807\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26785\ : std_logic;
signal \N__26782\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26752\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26744\ : std_logic;
signal \N__26743\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26713\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26663\ : std_logic;
signal \N__26660\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26626\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26620\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26614\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26608\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26576\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26560\ : std_logic;
signal \N__26557\ : std_logic;
signal \N__26554\ : std_logic;
signal \N__26551\ : std_logic;
signal \N__26550\ : std_logic;
signal \N__26547\ : std_logic;
signal \N__26544\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26520\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26516\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26513\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26478\ : std_logic;
signal \N__26475\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26369\ : std_logic;
signal \N__26366\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26356\ : std_logic;
signal \N__26353\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26315\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26300\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26279\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26270\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26261\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26015\ : std_logic;
signal \N__26012\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25997\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25988\ : std_logic;
signal \N__25985\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25979\ : std_logic;
signal \N__25976\ : std_logic;
signal \N__25973\ : std_logic;
signal \N__25970\ : std_logic;
signal \N__25967\ : std_logic;
signal \N__25964\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25943\ : std_logic;
signal \N__25940\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25907\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25871\ : std_logic;
signal \N__25868\ : std_logic;
signal \N__25865\ : std_logic;
signal \N__25862\ : std_logic;
signal \N__25859\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25761\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25680\ : std_logic;
signal \N__25677\ : std_logic;
signal \N__25674\ : std_logic;
signal \N__25667\ : std_logic;
signal \N__25664\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25649\ : std_logic;
signal \N__25646\ : std_logic;
signal \N__25643\ : std_logic;
signal \N__25640\ : std_logic;
signal \N__25637\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25601\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25571\ : std_logic;
signal \N__25568\ : std_logic;
signal \N__25565\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25547\ : std_logic;
signal \N__25544\ : std_logic;
signal \N__25541\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25499\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25472\ : std_logic;
signal \N__25469\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25445\ : std_logic;
signal \N__25442\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25438\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25411\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25403\ : std_logic;
signal \N__25400\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25391\ : std_logic;
signal \N__25388\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25345\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25158\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25152\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25134\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25062\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25049\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25022\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24979\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24915\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24827\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24805\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24709\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24689\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24676\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24664\ : std_logic;
signal \N__24659\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24650\ : std_logic;
signal \N__24647\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24607\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24581\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24575\ : std_logic;
signal \N__24572\ : std_logic;
signal \N__24569\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24487\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24428\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24418\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24398\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24386\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24331\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24250\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24071\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24026\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23980\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23924\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23826\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23789\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23675\ : std_logic;
signal \N__23672\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23645\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23633\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23476\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23407\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23396\ : std_logic;
signal \N__23393\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23314\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23186\ : std_logic;
signal \N__23183\ : std_logic;
signal \N__23180\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23054\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23050\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22950\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22754\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22730\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22666\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22364\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22139\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22042\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21734\ : std_logic;
signal \N__21731\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21445\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21425\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21419\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21404\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21316\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21204\ : std_logic;
signal \N__21201\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20786\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20624\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20474\ : std_logic;
signal \N__20471\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20438\ : std_logic;
signal \N__20435\ : std_logic;
signal \N__20432\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20393\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19931\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19787\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19754\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19379\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19289\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18917\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18866\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18857\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18841\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18677\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18530\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18518\ : std_logic;
signal \N__18515\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18377\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18350\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18332\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18125\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17984\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17942\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17327\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16793\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15932\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \CLK_pad_gb_input\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \LED_c\ : std_logic;
signal n26 : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal n25 : std_logic;
signal n3906 : std_logic;
signal n24 : std_logic;
signal n3907 : std_logic;
signal n23 : std_logic;
signal n3908 : std_logic;
signal n22 : std_logic;
signal n3909 : std_logic;
signal n21 : std_logic;
signal n3910 : std_logic;
signal n20 : std_logic;
signal n3911 : std_logic;
signal n19 : std_logic;
signal n3912 : std_logic;
signal n3913 : std_logic;
signal n18 : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal n17 : std_logic;
signal n3914 : std_logic;
signal n16 : std_logic;
signal n3915 : std_logic;
signal n15 : std_logic;
signal n3916 : std_logic;
signal n14 : std_logic;
signal n3917 : std_logic;
signal n13 : std_logic;
signal n3918 : std_logic;
signal n12 : std_logic;
signal n3919 : std_logic;
signal n11_adj_364 : std_logic;
signal n3920 : std_logic;
signal n3921 : std_logic;
signal n10_adj_363 : std_logic;
signal \bfn_17_19_0_\ : std_logic;
signal n9 : std_logic;
signal n3922 : std_logic;
signal n8_adj_362 : std_logic;
signal n3923 : std_logic;
signal n7 : std_logic;
signal n3924 : std_logic;
signal n6 : std_logic;
signal n3925 : std_logic;
signal n3926 : std_logic;
signal n3927 : std_logic;
signal n3928 : std_logic;
signal n3929 : std_logic;
signal \bfn_17_20_0_\ : std_logic;
signal n3930 : std_logic;
signal blink_counter_25 : std_logic;
signal \bfn_17_21_0_\ : std_logic;
signal \eeprom.n4183\ : std_logic;
signal \eeprom.n4184\ : std_logic;
signal \eeprom.n4185\ : std_logic;
signal \eeprom.n4186\ : std_logic;
signal \eeprom.n4187\ : std_logic;
signal \eeprom.n4188\ : std_logic;
signal \eeprom.n4189\ : std_logic;
signal \eeprom.n4190\ : std_logic;
signal \bfn_17_22_0_\ : std_logic;
signal \eeprom.n4191\ : std_logic;
signal \eeprom.n4192\ : std_logic;
signal \eeprom.n4193\ : std_logic;
signal \eeprom.n4194\ : std_logic;
signal \eeprom.n4195\ : std_logic;
signal \eeprom.n4196\ : std_logic;
signal \eeprom.n4197\ : std_logic;
signal \eeprom.n4198\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \eeprom.n4199\ : std_logic;
signal \eeprom.n4200\ : std_logic;
signal \eeprom.n4201\ : std_logic;
signal \eeprom.n4202\ : std_logic;
signal \eeprom.n4203\ : std_logic;
signal \eeprom.n4204\ : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal \eeprom.n4162\ : std_logic;
signal \eeprom.n4163\ : std_logic;
signal \eeprom.n4164\ : std_logic;
signal \eeprom.n4165\ : std_logic;
signal \eeprom.n4166\ : std_logic;
signal \eeprom.n4167\ : std_logic;
signal \eeprom.n4168\ : std_logic;
signal \eeprom.n4169\ : std_logic;
signal \bfn_17_25_0_\ : std_logic;
signal \eeprom.n4170\ : std_logic;
signal \eeprom.n4171\ : std_logic;
signal \eeprom.n4172\ : std_logic;
signal \eeprom.n4173\ : std_logic;
signal \eeprom.n4174\ : std_logic;
signal \eeprom.n3372\ : std_logic;
signal \eeprom.n4175\ : std_logic;
signal \eeprom.n4176\ : std_logic;
signal \eeprom.n4177\ : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal \eeprom.n4178\ : std_logic;
signal \eeprom.n4179\ : std_logic;
signal \eeprom.n4180\ : std_logic;
signal \eeprom.n4181\ : std_logic;
signal \eeprom.n4182\ : std_logic;
signal \bfn_17_27_0_\ : std_logic;
signal \eeprom.n4142\ : std_logic;
signal \eeprom.n4143\ : std_logic;
signal \eeprom.n4144\ : std_logic;
signal \eeprom.n4145\ : std_logic;
signal \eeprom.n4146\ : std_logic;
signal \eeprom.n4147\ : std_logic;
signal \eeprom.n4148\ : std_logic;
signal \eeprom.n4149\ : std_logic;
signal \bfn_17_28_0_\ : std_logic;
signal \eeprom.n3277\ : std_logic;
signal \eeprom.n4150\ : std_logic;
signal \eeprom.n4151\ : std_logic;
signal \eeprom.n4152\ : std_logic;
signal \eeprom.n4153\ : std_logic;
signal \eeprom.n4154\ : std_logic;
signal \eeprom.n4155\ : std_logic;
signal \eeprom.n4156\ : std_logic;
signal \eeprom.n4157\ : std_logic;
signal \bfn_17_29_0_\ : std_logic;
signal \eeprom.n4158\ : std_logic;
signal \eeprom.n4159\ : std_logic;
signal \eeprom.n4160\ : std_logic;
signal \eeprom.n4161\ : std_logic;
signal \bfn_18_17_0_\ : std_logic;
signal \eeprom.n3966\ : std_logic;
signal \eeprom.n3967\ : std_logic;
signal \eeprom.n3968\ : std_logic;
signal \eeprom.n3969\ : std_logic;
signal \eeprom.n3970\ : std_logic;
signal \eeprom.n3971\ : std_logic;
signal \eeprom.n3972\ : std_logic;
signal n5421 : std_logic;
signal blink_counter_24 : std_logic;
signal blink_counter_22 : std_logic;
signal blink_counter_23 : std_logic;
signal blink_counter_21 : std_logic;
signal n5420 : std_logic;
signal \eeprom.n1203\ : std_logic;
signal \eeprom.n3713_cascade_\ : std_logic;
signal \eeprom.n3618_cascade_\ : std_logic;
signal \eeprom.n3615_cascade_\ : std_logic;
signal \eeprom.n5221_cascade_\ : std_logic;
signal \eeprom.n5225\ : std_logic;
signal \eeprom.n3614\ : std_logic;
signal \eeprom.n3605\ : std_logic;
signal \eeprom.n3471\ : std_logic;
signal \eeprom.n32_cascade_\ : std_logic;
signal \eeprom.n3529_cascade_\ : std_logic;
signal \eeprom.n3481\ : std_logic;
signal \eeprom.n3513_cascade_\ : std_logic;
signal \eeprom.n3473\ : std_logic;
signal \eeprom.n3505_cascade_\ : std_logic;
signal \eeprom.n30_adj_273\ : std_logic;
signal \eeprom.n3478\ : std_logic;
signal \eeprom.n3472\ : std_logic;
signal \eeprom.n3484\ : std_logic;
signal \eeprom.n3475\ : std_logic;
signal \eeprom.n3507_cascade_\ : std_logic;
signal \eeprom.n31\ : std_logic;
signal \eeprom.n3482\ : std_logic;
signal \eeprom.n3514_cascade_\ : std_logic;
signal \eeprom.n5323_cascade_\ : std_logic;
signal \eeprom.n5321\ : std_logic;
signal \eeprom.n4753\ : std_logic;
signal \eeprom.n3376\ : std_logic;
signal \eeprom.n3380\ : std_logic;
signal \eeprom.n3412\ : std_logic;
signal \eeprom.n3412_cascade_\ : std_logic;
signal \eeprom.n3479\ : std_logic;
signal \eeprom.n3375\ : std_logic;
signal \eeprom.n3378\ : std_logic;
signal \eeprom.n3410\ : std_logic;
signal \eeprom.n3477\ : std_logic;
signal \eeprom.n3410_cascade_\ : std_logic;
signal \eeprom.n3465\ : std_logic;
signal \eeprom.n3367\ : std_logic;
signal \eeprom.n3267\ : std_logic;
signal \eeprom.n3299_cascade_\ : std_logic;
signal \eeprom.n3298\ : std_logic;
signal \eeprom.n3379\ : std_logic;
signal \eeprom.n3299\ : std_logic;
signal \eeprom.n3366\ : std_logic;
signal \eeprom.n3269\ : std_logic;
signal \eeprom.n3301\ : std_logic;
signal \eeprom.n3301_cascade_\ : std_logic;
signal \eeprom.n3368\ : std_logic;
signal \eeprom.n3374\ : std_logic;
signal \eeprom.n3406\ : std_logic;
signal \eeprom.n3370\ : std_logic;
signal \eeprom.n3268\ : std_logic;
signal \eeprom.n3300\ : std_logic;
signal \eeprom.n3200\ : std_logic;
signal \eeprom.n3200_cascade_\ : std_logic;
signal \eeprom.n3286\ : std_logic;
signal \eeprom.n3280\ : std_logic;
signal \eeprom.n3275\ : std_logic;
signal \eeprom.n3276\ : std_logic;
signal \eeprom.n3279\ : std_logic;
signal \eeprom.n3204_cascade_\ : std_logic;
signal \eeprom.n3273\ : std_logic;
signal \eeprom.n3206_cascade_\ : std_logic;
signal \eeprom.n3108_cascade_\ : std_logic;
signal \eeprom.n3202\ : std_logic;
signal \eeprom.n3201\ : std_logic;
signal \eeprom.n3203\ : std_logic;
signal \eeprom.n3270\ : std_logic;
signal \eeprom.n3203_cascade_\ : std_logic;
signal \eeprom.n3113_cascade_\ : std_logic;
signal \eeprom.n5305_cascade_\ : std_logic;
signal \eeprom.n3034_cascade_\ : std_logic;
signal \bfn_18_29_0_\ : std_logic;
signal \eeprom.n3085\ : std_logic;
signal \eeprom.n4105\ : std_logic;
signal \eeprom.n3084\ : std_logic;
signal \eeprom.n4106\ : std_logic;
signal \eeprom.n3083\ : std_logic;
signal \eeprom.n4107\ : std_logic;
signal \eeprom.n4108\ : std_logic;
signal \eeprom.n3081\ : std_logic;
signal \eeprom.n4109\ : std_logic;
signal \eeprom.n4110\ : std_logic;
signal \eeprom.n3079\ : std_logic;
signal \eeprom.n4111\ : std_logic;
signal \eeprom.n4112\ : std_logic;
signal \bfn_18_30_0_\ : std_logic;
signal \eeprom.n3077\ : std_logic;
signal \eeprom.n4113\ : std_logic;
signal \eeprom.n3076\ : std_logic;
signal \eeprom.n4114\ : std_logic;
signal \eeprom.n3075\ : std_logic;
signal \eeprom.n4115\ : std_logic;
signal \eeprom.n4116\ : std_logic;
signal \eeprom.n4117\ : std_logic;
signal \eeprom.n4118\ : std_logic;
signal \eeprom.n4119\ : std_logic;
signal \eeprom.n4120\ : std_logic;
signal \eeprom.n3070\ : std_logic;
signal \bfn_18_31_0_\ : std_logic;
signal \eeprom.n3069\ : std_logic;
signal \eeprom.n4121\ : std_logic;
signal \eeprom.n4122\ : std_logic;
signal \eeprom.n3071\ : std_logic;
signal \eeprom.n3004\ : std_logic;
signal \eeprom.n3613\ : std_logic;
signal \eeprom.n1202\ : std_logic;
signal \eeprom.n3712_cascade_\ : std_logic;
signal \eeprom.n1207\ : std_logic;
signal \eeprom.n3618\ : std_logic;
signal \eeprom.n3717_cascade_\ : std_logic;
signal \eeprom.n1208\ : std_logic;
signal \eeprom.n5362_cascade_\ : std_logic;
signal \eeprom.n1206\ : std_logic;
signal \eeprom.n1205\ : std_logic;
signal \eeprom.n3616\ : std_logic;
signal \eeprom.n3715_cascade_\ : std_logic;
signal \eeprom.n5017\ : std_logic;
signal \eeprom.n5019_cascade_\ : std_logic;
signal \eeprom.n28_adj_342_cascade_\ : std_logic;
signal \eeprom.n3615\ : std_logic;
signal \eeprom.n3628_cascade_\ : std_logic;
signal \eeprom.n1204\ : std_logic;
signal \eeprom.n3714_cascade_\ : std_logic;
signal \eeprom.n1201\ : std_logic;
signal \eeprom.n3628\ : std_logic;
signal \eeprom.n5025_cascade_\ : std_logic;
signal \eeprom.n5027_cascade_\ : std_logic;
signal \eeprom.n5029_cascade_\ : std_logic;
signal \eeprom.n5031_cascade_\ : std_logic;
signal \eeprom.n5161\ : std_logic;
signal \eeprom.n29_adj_274\ : std_logic;
signal \eeprom.n3612\ : std_logic;
signal \eeprom.n3617\ : std_logic;
signal \eeprom.n3596\ : std_logic;
signal \eeprom.n3609_cascade_\ : std_logic;
signal \eeprom.n5021_cascade_\ : std_logic;
signal \eeprom.n5023\ : std_logic;
signal \eeprom.n3474\ : std_logic;
signal \eeprom.n3407\ : std_logic;
signal \eeprom.n3486\ : std_logic;
signal \eeprom.n3468\ : std_logic;
signal \eeprom.n3608_cascade_\ : std_logic;
signal \eeprom.n3480\ : std_logic;
signal \eeprom.n3512_cascade_\ : std_logic;
signal \eeprom.n5175\ : std_logic;
signal \eeprom.n5177_cascade_\ : std_logic;
signal \eeprom.n31_adj_341\ : std_logic;
signal \eeprom.n3598\ : std_logic;
signal \eeprom.n3483\ : std_logic;
signal \eeprom.n3485\ : std_logic;
signal \eeprom.n3398\ : std_logic;
signal \eeprom.n3397\ : std_logic;
signal \eeprom.n3408\ : std_logic;
signal \eeprom.n3411\ : std_logic;
signal \eeprom.n18_cascade_\ : std_logic;
signal \eeprom.n29\ : std_logic;
signal \eeprom.n30_cascade_\ : std_logic;
signal \eeprom.n3430_cascade_\ : std_logic;
signal \eeprom.n3467\ : std_logic;
signal \eeprom.n3466\ : std_logic;
signal \eeprom.n3498_cascade_\ : std_logic;
signal \eeprom.n28_adj_267\ : std_logic;
signal \eeprom.n3476\ : std_logic;
signal \eeprom.n3373\ : std_logic;
signal \eeprom.n3369\ : std_logic;
signal \eeprom.n3401\ : std_logic;
signal \eeprom.n3400\ : std_logic;
signal \eeprom.n3399\ : std_logic;
signal \eeprom.n3401_cascade_\ : std_logic;
signal \eeprom.n27_adj_263\ : std_logic;
signal \eeprom.n3402\ : std_logic;
signal \eeprom.n3469\ : std_logic;
signal \eeprom.n3307\ : std_logic;
signal \eeprom.n3311\ : std_logic;
signal \eeprom.n3312\ : std_logic;
signal \eeprom.n3309\ : std_logic;
signal \eeprom.n28_cascade_\ : std_logic;
signal \eeprom.n25\ : std_logic;
signal \eeprom.n3385\ : std_logic;
signal \eeprom.n3331_cascade_\ : std_logic;
signal \eeprom.n3281\ : std_logic;
signal \eeprom.n3206\ : std_logic;
signal \eeprom.n20_adj_301_cascade_\ : std_logic;
signal \eeprom.n16_adj_303\ : std_logic;
signal \eeprom.n3212\ : std_logic;
signal \eeprom.n28_adj_305_cascade_\ : std_logic;
signal \eeprom.n24_adj_304\ : std_logic;
signal \eeprom.n3232_cascade_\ : std_logic;
signal \eeprom.n3274\ : std_logic;
signal \eeprom.n3306\ : std_logic;
signal \eeprom.n3305\ : std_logic;
signal \eeprom.n3306_cascade_\ : std_logic;
signal \eeprom.n3308\ : std_logic;
signal \eeprom.n27\ : std_logic;
signal \eeprom.n5309\ : std_logic;
signal \eeprom.n18_adj_260_cascade_\ : std_logic;
signal \eeprom.n24\ : std_logic;
signal \eeprom.n22\ : std_logic;
signal \eeprom.n26_adj_262_cascade_\ : std_logic;
signal \eeprom.n3133_cascade_\ : std_logic;
signal \eeprom.n3205\ : std_logic;
signal \eeprom.n3272\ : std_logic;
signal \eeprom.n3205_cascade_\ : std_logic;
signal \eeprom.n3204\ : std_logic;
signal \eeprom.n3271\ : std_logic;
signal \eeprom.n3207\ : std_logic;
signal \eeprom.n3017\ : std_logic;
signal \eeprom.n3017_cascade_\ : std_logic;
signal \eeprom.n5147_cascade_\ : std_logic;
signal \eeprom.n3009\ : std_logic;
signal \eeprom.n3002\ : std_logic;
signal \eeprom.n3002_cascade_\ : std_logic;
signal \eeprom.n20_adj_337\ : std_logic;
signal \eeprom.n3078\ : std_logic;
signal \eeprom.n3016\ : std_logic;
signal \eeprom.n3018\ : std_logic;
signal \eeprom.n2914_cascade_\ : std_logic;
signal \eeprom.n3073\ : std_logic;
signal \eeprom.n3014\ : std_logic;
signal \eeprom.n3007\ : std_logic;
signal \eeprom.n3074\ : std_logic;
signal \eeprom.n3007_cascade_\ : std_logic;
signal \eeprom.n3006\ : std_logic;
signal \eeprom.n21_adj_336\ : std_logic;
signal \eeprom.n3006_cascade_\ : std_logic;
signal \eeprom.n18_adj_335\ : std_logic;
signal \eeprom.n24_adj_340\ : std_logic;
signal \eeprom.n3008\ : std_logic;
signal \eeprom.n3005\ : std_logic;
signal \eeprom.n3005_cascade_\ : std_logic;
signal \eeprom.n3072\ : std_logic;
signal \eeprom.n3082\ : std_logic;
signal \eeprom.n3010\ : std_logic;
signal \eeprom.n3012\ : std_logic;
signal \eeprom.n3003\ : std_logic;
signal \eeprom.n3086\ : std_logic;
signal \eeprom.n3186\ : std_logic;
signal \bfn_19_30_0_\ : std_logic;
signal \eeprom.n4123\ : std_logic;
signal \eeprom.n3117\ : std_logic;
signal \eeprom.n3184\ : std_logic;
signal \eeprom.n4124\ : std_logic;
signal \eeprom.n4125\ : std_logic;
signal \eeprom.n4126\ : std_logic;
signal \eeprom.n4127\ : std_logic;
signal \eeprom.n3113\ : std_logic;
signal \eeprom.n3180\ : std_logic;
signal \eeprom.n4128\ : std_logic;
signal \eeprom.n3179\ : std_logic;
signal \eeprom.n4129\ : std_logic;
signal \eeprom.n4130\ : std_logic;
signal \eeprom.n3111\ : std_logic;
signal \eeprom.n3178\ : std_logic;
signal \bfn_19_31_0_\ : std_logic;
signal \eeprom.n4131\ : std_logic;
signal \eeprom.n4132\ : std_logic;
signal \eeprom.n3108\ : std_logic;
signal \eeprom.n3175\ : std_logic;
signal \eeprom.n4133\ : std_logic;
signal \eeprom.n3107\ : std_logic;
signal \eeprom.n3174\ : std_logic;
signal \eeprom.n4134\ : std_logic;
signal \eeprom.n3106\ : std_logic;
signal \eeprom.n3173\ : std_logic;
signal \eeprom.n4135\ : std_logic;
signal \eeprom.n3105\ : std_logic;
signal \eeprom.n3172\ : std_logic;
signal \eeprom.n4136\ : std_logic;
signal \eeprom.n3104\ : std_logic;
signal \eeprom.n3171\ : std_logic;
signal \eeprom.n4137\ : std_logic;
signal \eeprom.n4138\ : std_logic;
signal \eeprom.n3103\ : std_logic;
signal \eeprom.n3170\ : std_logic;
signal \bfn_19_32_0_\ : std_logic;
signal \eeprom.n3102\ : std_logic;
signal \eeprom.n3169\ : std_logic;
signal \eeprom.n4139\ : std_logic;
signal \eeprom.n3101\ : std_logic;
signal \eeprom.n3168\ : std_logic;
signal \eeprom.n4140\ : std_logic;
signal \eeprom.n3100\ : std_logic;
signal \eeprom.n4141\ : std_logic;
signal \eeprom.n3199\ : std_logic;
signal \bfn_20_17_0_\ : std_logic;
signal \eeprom.n4228\ : std_logic;
signal \eeprom.n4229\ : std_logic;
signal \eeprom.n4230\ : std_logic;
signal \eeprom.n4231\ : std_logic;
signal \eeprom.n4232\ : std_logic;
signal \eeprom.n4233\ : std_logic;
signal \eeprom.n5547\ : std_logic;
signal \eeprom.n5362\ : std_logic;
signal \eeprom.n4234\ : std_logic;
signal \eeprom.n4235\ : std_logic;
signal \eeprom.n5550\ : std_logic;
signal \eeprom.n3717\ : std_logic;
signal \bfn_20_18_0_\ : std_logic;
signal \eeprom.n4236\ : std_logic;
signal \eeprom.n5556\ : std_logic;
signal \eeprom.n3715\ : std_logic;
signal \eeprom.n4237\ : std_logic;
signal \eeprom.n5559\ : std_logic;
signal \eeprom.n3714\ : std_logic;
signal \eeprom.n4238\ : std_logic;
signal \eeprom.n5562\ : std_logic;
signal \eeprom.n3713\ : std_logic;
signal \eeprom.n4239\ : std_logic;
signal \eeprom.n5565\ : std_logic;
signal \eeprom.n3712\ : std_logic;
signal \eeprom.n4240\ : std_logic;
signal \eeprom.n3711\ : std_logic;
signal \eeprom.n5568\ : std_logic;
signal \eeprom.n4241\ : std_logic;
signal \eeprom.n3716\ : std_logic;
signal \eeprom.n5553\ : std_logic;
signal \eeprom.n3586\ : std_logic;
signal \bfn_20_19_0_\ : std_logic;
signal \eeprom.n3518\ : std_logic;
signal \eeprom.n3585_adj_296\ : std_logic;
signal \eeprom.n4205\ : std_logic;
signal \eeprom.n3517\ : std_logic;
signal \eeprom.n3584\ : std_logic;
signal \eeprom.n4206\ : std_logic;
signal \eeprom.n3516\ : std_logic;
signal \eeprom.n3583\ : std_logic;
signal \eeprom.n4207\ : std_logic;
signal \eeprom.n3515\ : std_logic;
signal \eeprom.n3582\ : std_logic;
signal \eeprom.n4208\ : std_logic;
signal \eeprom.n3514\ : std_logic;
signal \eeprom.n3581_adj_292\ : std_logic;
signal \eeprom.n4209\ : std_logic;
signal \eeprom.n3513\ : std_logic;
signal \eeprom.n3580\ : std_logic;
signal \eeprom.n4210\ : std_logic;
signal \eeprom.n3512\ : std_logic;
signal \eeprom.n3579\ : std_logic;
signal \eeprom.n4211\ : std_logic;
signal \eeprom.n4212\ : std_logic;
signal \eeprom.n3511\ : std_logic;
signal \eeprom.n3578\ : std_logic;
signal \bfn_20_20_0_\ : std_logic;
signal \eeprom.n3510\ : std_logic;
signal \eeprom.n3577\ : std_logic;
signal \eeprom.n4213\ : std_logic;
signal \eeprom.n3509\ : std_logic;
signal \eeprom.n3576\ : std_logic;
signal \eeprom.n4214\ : std_logic;
signal \eeprom.n3508\ : std_logic;
signal \eeprom.n3575\ : std_logic;
signal \eeprom.n4215\ : std_logic;
signal \eeprom.n3507\ : std_logic;
signal \eeprom.n3574\ : std_logic;
signal \eeprom.n4216\ : std_logic;
signal \eeprom.n3506\ : std_logic;
signal \eeprom.n3573\ : std_logic;
signal \eeprom.n4217\ : std_logic;
signal \eeprom.n3505\ : std_logic;
signal \eeprom.n3572\ : std_logic;
signal \eeprom.n4218\ : std_logic;
signal \eeprom.n3504\ : std_logic;
signal \eeprom.n3571\ : std_logic;
signal \eeprom.n4219\ : std_logic;
signal \eeprom.n4220\ : std_logic;
signal \eeprom.n3503\ : std_logic;
signal \eeprom.n3570\ : std_logic;
signal \bfn_20_21_0_\ : std_logic;
signal \eeprom.n3569\ : std_logic;
signal \eeprom.n4221\ : std_logic;
signal \eeprom.n3501\ : std_logic;
signal \eeprom.n3568\ : std_logic;
signal \eeprom.n4222\ : std_logic;
signal \eeprom.n3500\ : std_logic;
signal \eeprom.n3567\ : std_logic;
signal \eeprom.n4223\ : std_logic;
signal \eeprom.n3499\ : std_logic;
signal \eeprom.n3566\ : std_logic;
signal \eeprom.n4224\ : std_logic;
signal \eeprom.n3498\ : std_logic;
signal \eeprom.n3565\ : std_logic;
signal \eeprom.n4225\ : std_logic;
signal \eeprom.n3497\ : std_logic;
signal \eeprom.n3564\ : std_logic;
signal \eeprom.n4226\ : std_logic;
signal \eeprom.n3496\ : std_logic;
signal \eeprom.n3529\ : std_logic;
signal \eeprom.n4227\ : std_logic;
signal \eeprom.n5355\ : std_logic;
signal \eeprom.n3382\ : std_logic;
signal \eeprom.n3414\ : std_logic;
signal \eeprom.n3417\ : std_logic;
signal \eeprom.n3414_cascade_\ : std_logic;
signal \eeprom.n5291_cascade_\ : std_logic;
signal \eeprom.n3405\ : std_logic;
signal \eeprom.n4824_cascade_\ : std_logic;
signal \eeprom.n3404\ : std_logic;
signal \eeprom.n28_adj_261\ : std_logic;
signal \eeprom.n3386\ : std_logic;
signal \eeprom.n3418\ : std_logic;
signal \eeprom.n3384\ : std_logic;
signal \eeprom.n3416\ : std_logic;
signal \eeprom.n3383\ : std_logic;
signal \eeprom.n3313\ : std_logic;
signal \eeprom.n3371\ : std_logic;
signal \eeprom.n3282\ : std_logic;
signal \eeprom.n3381\ : std_logic;
signal \eeprom.n3314_cascade_\ : std_logic;
signal \eeprom.n3413\ : std_logic;
signal \eeprom.n3413_cascade_\ : std_logic;
signal \eeprom.n3415\ : std_logic;
signal \eeprom.n5289\ : std_logic;
signal \eeprom.n3278\ : std_logic;
signal \eeprom.n3310\ : std_logic;
signal \eeprom.n3331\ : std_logic;
signal \eeprom.n3310_cascade_\ : std_logic;
signal \eeprom.n3377\ : std_logic;
signal \eeprom.n3409\ : std_logic;
signal \eeprom.n3284\ : std_logic;
signal \eeprom.n3218\ : std_logic;
signal \eeprom.n3285\ : std_logic;
signal \eeprom.n3317\ : std_logic;
signal \eeprom.n3314\ : std_logic;
signal \eeprom.n3317_cascade_\ : std_logic;
signal \eeprom.n3316\ : std_logic;
signal \eeprom.n3318\ : std_logic;
signal \eeprom.n5315_cascade_\ : std_logic;
signal \eeprom.n5313\ : std_logic;
signal \eeprom.n3303\ : std_logic;
signal \eeprom.n3304\ : std_logic;
signal \eeprom.n4820_cascade_\ : std_logic;
signal \eeprom.n3302\ : std_logic;
signal \eeprom.n26\ : std_logic;
signal \eeprom.n3283\ : std_logic;
signal \eeprom.n3232\ : std_logic;
signal \eeprom.n3315\ : std_logic;
signal \eeprom.n3114\ : std_logic;
signal \eeprom.n3181\ : std_logic;
signal \eeprom.n3213\ : std_logic;
signal \eeprom.n3213_cascade_\ : std_logic;
signal \eeprom.n3182\ : std_logic;
signal \eeprom.n3115\ : std_logic;
signal \eeprom.n3214\ : std_logic;
signal \eeprom.n3216\ : std_logic;
signal \eeprom.n3214_cascade_\ : std_logic;
signal \eeprom.n5205\ : std_logic;
signal \eeprom.n5209\ : std_logic;
signal \eeprom.n3116\ : std_logic;
signal \eeprom.n3183\ : std_logic;
signal \eeprom.n3215\ : std_logic;
signal \eeprom.n3185\ : std_logic;
signal \eeprom.n3118\ : std_logic;
signal \eeprom.n3217\ : std_logic;
signal \eeprom.n3109\ : std_logic;
signal \eeprom.n3176\ : std_logic;
signal \eeprom.n3208\ : std_logic;
signal \eeprom.n3211\ : std_logic;
signal \eeprom.n3208_cascade_\ : std_logic;
signal \eeprom.n3210\ : std_logic;
signal \eeprom.n26_adj_302\ : std_logic;
signal \eeprom.n3080\ : std_logic;
signal \eeprom.n3013_cascade_\ : std_logic;
signal \eeprom.n3034\ : std_logic;
signal \eeprom.n3112\ : std_logic;
signal \eeprom.n3011\ : std_logic;
signal \eeprom.n5301\ : std_logic;
signal \eeprom.n3110\ : std_logic;
signal \eeprom.n3133\ : std_logic;
signal \eeprom.n3177\ : std_logic;
signal \eeprom.n3209\ : std_logic;
signal \eeprom.n2910_cascade_\ : std_logic;
signal \eeprom.n15_adj_300\ : std_logic;
signal \eeprom.n22_adj_331_cascade_\ : std_logic;
signal \eeprom.n18_adj_330\ : std_logic;
signal \eeprom.n2935_cascade_\ : std_logic;
signal \eeprom.n3015\ : std_logic;
signal \eeprom.n3013\ : std_logic;
signal \eeprom.n3015_cascade_\ : std_logic;
signal \eeprom.n5143\ : std_logic;
signal \eeprom.n18_adj_290_cascade_\ : std_logic;
signal \eeprom.n20_adj_291_cascade_\ : std_logic;
signal \eeprom.n2836_cascade_\ : std_logic;
signal \eeprom.n2913_cascade_\ : std_logic;
signal \eeprom.n5297\ : std_logic;
signal \eeprom.n2986\ : std_logic;
signal \bfn_20_29_0_\ : std_logic;
signal \eeprom.n2985\ : std_logic;
signal \eeprom.n4088\ : std_logic;
signal \eeprom.n2917\ : std_logic;
signal \eeprom.n2984\ : std_logic;
signal \eeprom.n4089\ : std_logic;
signal \eeprom.n2916\ : std_logic;
signal \eeprom.n2983\ : std_logic;
signal \eeprom.n4090\ : std_logic;
signal \eeprom.n2915\ : std_logic;
signal \eeprom.n2982\ : std_logic;
signal \eeprom.n4091\ : std_logic;
signal \eeprom.n2914\ : std_logic;
signal \eeprom.n2981\ : std_logic;
signal \eeprom.n4092\ : std_logic;
signal \eeprom.n2913\ : std_logic;
signal \eeprom.n2980\ : std_logic;
signal \eeprom.n4093\ : std_logic;
signal \eeprom.n2979\ : std_logic;
signal \eeprom.n4094\ : std_logic;
signal \eeprom.n4095\ : std_logic;
signal \eeprom.n2978\ : std_logic;
signal \bfn_20_30_0_\ : std_logic;
signal \eeprom.n2910\ : std_logic;
signal \eeprom.n2977\ : std_logic;
signal \eeprom.n4096\ : std_logic;
signal \eeprom.n2909\ : std_logic;
signal \eeprom.n2976\ : std_logic;
signal \eeprom.n4097\ : std_logic;
signal \eeprom.n2908\ : std_logic;
signal \eeprom.n2975\ : std_logic;
signal \eeprom.n4098\ : std_logic;
signal \eeprom.n2974\ : std_logic;
signal \eeprom.n4099\ : std_logic;
signal \eeprom.n2906\ : std_logic;
signal \eeprom.n2973\ : std_logic;
signal \eeprom.n4100\ : std_logic;
signal \eeprom.n2972\ : std_logic;
signal \eeprom.n4101\ : std_logic;
signal \eeprom.n2971\ : std_logic;
signal \eeprom.n4102\ : std_logic;
signal \eeprom.n4103\ : std_logic;
signal \eeprom.n2970\ : std_logic;
signal \bfn_20_31_0_\ : std_logic;
signal \eeprom.n2935\ : std_logic;
signal \eeprom.n4104\ : std_logic;
signal \eeprom.n3001\ : std_logic;
signal \eeprom.enable_N_60_0\ : std_logic;
signal \eeprom.enable_N_60_1\ : std_logic;
signal \eeprom.enable_N_60_2\ : std_logic;
signal \eeprom.enable_N_60_3\ : std_logic;
signal \eeprom.enable_N_60_4\ : std_logic;
signal \eeprom.n4847_cascade_\ : std_logic;
signal \eeprom.enable_N_60_5\ : std_logic;
signal \eeprom.enable_N_60_7\ : std_logic;
signal \eeprom.enable_N_60_6\ : std_logic;
signal \eeprom.n4853_cascade_\ : std_logic;
signal \eeprom.enable_N_60_8\ : std_logic;
signal \eeprom.enable_N_60_10\ : std_logic;
signal \eeprom.enable_N_60_9\ : std_logic;
signal \eeprom.n4859_cascade_\ : std_logic;
signal \eeprom.enable_N_60_11\ : std_logic;
signal \eeprom.n4865_cascade_\ : std_logic;
signal \eeprom.enable_N_59_cascade_\ : std_logic;
signal \eeprom.enable_N_60_12\ : std_logic;
signal \eeprom.enable_N_60_14\ : std_logic;
signal \eeprom.enable_N_60_13\ : std_logic;
signal \eeprom.n4865\ : std_logic;
signal \eeprom.n2211_cascade_\ : std_logic;
signal \eeprom.n2214_cascade_\ : std_logic;
signal \eeprom.n3720\ : std_logic;
signal \bfn_21_20_0_\ : std_logic;
signal \eeprom.n4007\ : std_logic;
signal \eeprom.n4008\ : std_logic;
signal \eeprom.n4009\ : std_logic;
signal \eeprom.n4010\ : std_logic;
signal \eeprom.n4011\ : std_logic;
signal \eeprom.n4012\ : std_logic;
signal \eeprom.n4013\ : std_logic;
signal \eeprom.n4014\ : std_logic;
signal \bfn_21_21_0_\ : std_logic;
signal \eeprom.n4015\ : std_logic;
signal \eeprom.n4016\ : std_logic;
signal \eeprom.n4017\ : std_logic;
signal \eeprom.n3403\ : std_logic;
signal \eeprom.n3470\ : std_logic;
signal \eeprom.n3430\ : std_logic;
signal \eeprom.n3502\ : std_logic;
signal \eeprom.n2511_cascade_\ : std_logic;
signal \eeprom.n2618_cascade_\ : std_logic;
signal \bfn_21_23_0_\ : std_logic;
signal \eeprom.n2685\ : std_logic;
signal \eeprom.n4043\ : std_logic;
signal \eeprom.n4044\ : std_logic;
signal \eeprom.n4045\ : std_logic;
signal \eeprom.n4046\ : std_logic;
signal \eeprom.n4047\ : std_logic;
signal \eeprom.n4048\ : std_logic;
signal \eeprom.n4049\ : std_logic;
signal \eeprom.n4050\ : std_logic;
signal \bfn_21_24_0_\ : std_logic;
signal \eeprom.n4051\ : std_logic;
signal \eeprom.n4052\ : std_logic;
signal \eeprom.n4053\ : std_logic;
signal \eeprom.n4054\ : std_logic;
signal \eeprom.n4055\ : std_logic;
signal \eeprom.n4056\ : std_logic;
signal \eeprom.n2677\ : std_logic;
signal \eeprom.n2678\ : std_logic;
signal \eeprom.n2710_cascade_\ : std_logic;
signal \eeprom.n2686\ : std_logic;
signal \eeprom.n2912\ : std_logic;
signal \eeprom.n5157_cascade_\ : std_logic;
signal \eeprom.n16\ : std_logic;
signal \eeprom.n5153\ : std_logic;
signal \eeprom.n2918\ : std_logic;
signal \eeprom.n2911\ : std_logic;
signal \eeprom.n2886\ : std_logic;
signal \bfn_21_27_0_\ : std_logic;
signal \eeprom.n2885\ : std_logic;
signal \eeprom.n4072\ : std_logic;
signal \eeprom.n2884\ : std_logic;
signal \eeprom.n4073\ : std_logic;
signal \eeprom.n2883\ : std_logic;
signal \eeprom.n4074\ : std_logic;
signal \eeprom.n2882\ : std_logic;
signal \eeprom.n4075\ : std_logic;
signal \eeprom.n2881\ : std_logic;
signal \eeprom.n4076\ : std_logic;
signal \eeprom.n2880\ : std_logic;
signal \eeprom.n4077\ : std_logic;
signal \eeprom.n2879\ : std_logic;
signal \eeprom.n4078\ : std_logic;
signal \eeprom.n4079\ : std_logic;
signal \eeprom.n2878\ : std_logic;
signal \bfn_21_28_0_\ : std_logic;
signal \eeprom.n2877\ : std_logic;
signal \eeprom.n4080\ : std_logic;
signal \eeprom.n2876\ : std_logic;
signal \eeprom.n4081\ : std_logic;
signal \eeprom.n4082\ : std_logic;
signal \eeprom.n2874\ : std_logic;
signal \eeprom.n4083\ : std_logic;
signal \eeprom.n4084\ : std_logic;
signal \eeprom.n4085\ : std_logic;
signal \eeprom.n4086\ : std_logic;
signal \eeprom.n4087\ : std_logic;
signal \bfn_21_29_0_\ : std_logic;
signal \eeprom.n2902\ : std_logic;
signal \eeprom.n2902_cascade_\ : std_logic;
signal \eeprom.n19_adj_327\ : std_logic;
signal \eeprom.n2872\ : std_logic;
signal \eeprom.n2904\ : std_logic;
signal \eeprom.n2873\ : std_logic;
signal \eeprom.n2905\ : std_logic;
signal \eeprom.n2871\ : std_logic;
signal \eeprom.n2903\ : std_logic;
signal \eeprom.n2875\ : std_logic;
signal \eeprom.n2836\ : std_logic;
signal \eeprom.n2907\ : std_logic;
signal \bfn_22_17_0_\ : std_logic;
signal \eeprom.n2285\ : std_logic;
signal \eeprom.n3997\ : std_logic;
signal \eeprom.n3998\ : std_logic;
signal \eeprom.n2283\ : std_logic;
signal \eeprom.n3999\ : std_logic;
signal \eeprom.n2215\ : std_logic;
signal \eeprom.n4000\ : std_logic;
signal \eeprom.n2214\ : std_logic;
signal \eeprom.n2281\ : std_logic;
signal \eeprom.n4001\ : std_logic;
signal \eeprom.n4002\ : std_logic;
signal \eeprom.n4003\ : std_logic;
signal \eeprom.n4004\ : std_logic;
signal \eeprom.n2278\ : std_logic;
signal \bfn_22_18_0_\ : std_logic;
signal \eeprom.n4005\ : std_logic;
signal \eeprom.n4006\ : std_logic;
signal \eeprom.n2216\ : std_logic;
signal \eeprom.n2143_cascade_\ : std_logic;
signal \eeprom.n2286\ : std_logic;
signal \eeprom.n2218\ : std_logic;
signal \eeprom.n5045\ : std_logic;
signal \eeprom.n2211\ : std_logic;
signal \eeprom.n4797_cascade_\ : std_logic;
signal \eeprom.n2242_cascade_\ : std_logic;
signal \eeprom.n2282\ : std_logic;
signal \eeprom.n5400_cascade_\ : std_logic;
signal \eeprom.n2217\ : std_logic;
signal \eeprom.n2284\ : std_logic;
signal \eeprom.n2280\ : std_logic;
signal \eeprom.n2213\ : std_logic;
signal \eeprom.n5405\ : std_logic;
signal \eeprom.n2316\ : std_logic;
signal \eeprom.n2317\ : std_logic;
signal \eeprom.n2314\ : std_logic;
signal \eeprom.n2318\ : std_logic;
signal \eeprom.n5085_cascade_\ : std_logic;
signal \eeprom.n2310\ : std_logic;
signal \eeprom.n2315\ : std_logic;
signal \eeprom.n2313\ : std_logic;
signal \eeprom.n5081\ : std_logic;
signal \eeprom.n2277\ : std_logic;
signal \eeprom.n2309\ : std_logic;
signal \eeprom.n2309_cascade_\ : std_logic;
signal \eeprom.n2308\ : std_logic;
signal \eeprom.n2312\ : std_logic;
signal \eeprom.n8_adj_322_cascade_\ : std_logic;
signal \eeprom.n7_adj_323\ : std_logic;
signal \eeprom.n2341\ : std_logic;
signal \eeprom.n2341_cascade_\ : std_logic;
signal \eeprom.n5576\ : std_logic;
signal \eeprom.n2279\ : std_logic;
signal \eeprom.n2311\ : std_logic;
signal \eeprom.n5073_cascade_\ : std_logic;
signal \eeprom.n4782_cascade_\ : std_logic;
signal \eeprom.n12_cascade_\ : std_logic;
signal \eeprom.n2440_cascade_\ : std_logic;
signal \eeprom.n5071\ : std_logic;
signal \bfn_22_22_0_\ : std_logic;
signal \eeprom.n4018\ : std_logic;
signal \eeprom.n4019\ : std_logic;
signal \eeprom.n4020\ : std_logic;
signal \eeprom.n4021\ : std_logic;
signal \eeprom.n2414\ : std_logic;
signal \eeprom.n2481\ : std_logic;
signal \eeprom.n4022\ : std_logic;
signal \eeprom.n2413\ : std_logic;
signal \eeprom.n2480\ : std_logic;
signal \eeprom.n4023\ : std_logic;
signal \eeprom.n2412\ : std_logic;
signal \eeprom.n2479\ : std_logic;
signal \eeprom.n4024\ : std_logic;
signal \eeprom.n4025\ : std_logic;
signal \bfn_22_23_0_\ : std_logic;
signal \eeprom.n4026\ : std_logic;
signal \eeprom.n2409\ : std_logic;
signal \eeprom.n2476\ : std_logic;
signal \eeprom.n4027\ : std_logic;
signal \eeprom.n4028\ : std_logic;
signal \eeprom.n2407\ : std_logic;
signal \eeprom.n4029\ : std_logic;
signal \eeprom.n2638_cascade_\ : std_logic;
signal \eeprom.n2684\ : std_logic;
signal \eeprom.n2716_cascade_\ : std_logic;
signal \eeprom.n2680\ : std_logic;
signal \eeprom.n2679\ : std_logic;
signal \eeprom.n2676\ : std_logic;
signal \eeprom.n2675\ : std_logic;
signal \eeprom.n2673\ : std_logic;
signal \eeprom.n2705_cascade_\ : std_logic;
signal \eeprom.n17_adj_339\ : std_logic;
signal \eeprom.n16_adj_338_cascade_\ : std_logic;
signal \eeprom.n2737_cascade_\ : std_logic;
signal \eeprom.n2818\ : std_logic;
signal \bfn_22_25_0_\ : std_logic;
signal \eeprom.n2817\ : std_logic;
signal \eeprom.n4057\ : std_logic;
signal \eeprom.n2717\ : std_logic;
signal \eeprom.n2816\ : std_logic;
signal \eeprom.n4058\ : std_logic;
signal \eeprom.n2716\ : std_logic;
signal \eeprom.n2815\ : std_logic;
signal \eeprom.n4059\ : std_logic;
signal \eeprom.n2814\ : std_logic;
signal \eeprom.n4060\ : std_logic;
signal \eeprom.n2813\ : std_logic;
signal \eeprom.n4061\ : std_logic;
signal \eeprom.n5575\ : std_logic;
signal \eeprom.n2812\ : std_logic;
signal \eeprom.n4062\ : std_logic;
signal \eeprom.n2712\ : std_logic;
signal \eeprom.n2811\ : std_logic;
signal \eeprom.n4063\ : std_logic;
signal \eeprom.n4064\ : std_logic;
signal \eeprom.n2711\ : std_logic;
signal \eeprom.n2810\ : std_logic;
signal \bfn_22_26_0_\ : std_logic;
signal \eeprom.n2710\ : std_logic;
signal \eeprom.n2809\ : std_logic;
signal \eeprom.n4065\ : std_logic;
signal \eeprom.n2709\ : std_logic;
signal \eeprom.n2808\ : std_logic;
signal \eeprom.n4066\ : std_logic;
signal \eeprom.n2708\ : std_logic;
signal \eeprom.n2807\ : std_logic;
signal \eeprom.n4067\ : std_logic;
signal \eeprom.n2707\ : std_logic;
signal \eeprom.n2806\ : std_logic;
signal \eeprom.n4068\ : std_logic;
signal \eeprom.n2805\ : std_logic;
signal \eeprom.n4069\ : std_logic;
signal \eeprom.n2705\ : std_logic;
signal \eeprom.n2804\ : std_logic;
signal \eeprom.n4070\ : std_logic;
signal \eeprom.n2704\ : std_logic;
signal \eeprom.n2737\ : std_logic;
signal \eeprom.n4071\ : std_logic;
signal \eeprom.n2803\ : std_logic;
signal \eeprom.n5005_cascade_\ : std_logic;
signal \eeprom.n5009_cascade_\ : std_logic;
signal \eeprom.n2044_cascade_\ : std_logic;
signal \eeprom.n2116_cascade_\ : std_logic;
signal \bfn_23_18_0_\ : std_logic;
signal \eeprom.n2085\ : std_logic;
signal \eeprom.n3980\ : std_logic;
signal \eeprom.n2084\ : std_logic;
signal \eeprom.n3981\ : std_logic;
signal \eeprom.n3982\ : std_logic;
signal \eeprom.n2082\ : std_logic;
signal \eeprom.n3983\ : std_logic;
signal \eeprom.n3984\ : std_logic;
signal \eeprom.n2080\ : std_logic;
signal \eeprom.n3985\ : std_logic;
signal \eeprom.n3986\ : std_logic;
signal \eeprom.n3987\ : std_logic;
signal \bfn_23_19_0_\ : std_logic;
signal \eeprom.n2242\ : std_logic;
signal \eeprom.n5501\ : std_logic;
signal \eeprom.n2081\ : std_logic;
signal \eeprom.n2086\ : std_logic;
signal \eeprom.n5061\ : std_logic;
signal \eeprom.n2118_cascade_\ : std_logic;
signal \eeprom.n4788\ : std_logic;
signal \eeprom.n2212\ : std_logic;
signal \eeprom.n2019\ : std_logic;
signal \eeprom.n3721\ : std_logic;
signal \eeprom.n3619\ : std_logic;
signal \eeprom.n2219\ : std_logic;
signal \eeprom.n3723\ : std_logic;
signal \eeprom.n2210\ : std_logic;
signal \eeprom.n6_adj_321\ : std_logic;
signal \eeprom.n2483\ : std_logic;
signal \eeprom.n2416\ : std_logic;
signal \eeprom.n2485\ : std_logic;
signal \eeprom.n2418\ : std_logic;
signal \eeprom.n2477\ : std_logic;
signal \eeprom.n2410\ : std_logic;
signal \eeprom.n2408\ : std_logic;
signal \eeprom.n2475\ : std_logic;
signal \eeprom.n2486\ : std_logic;
signal \eeprom.n2484\ : std_logic;
signal \eeprom.n2417\ : std_logic;
signal \eeprom.n2482\ : std_logic;
signal \eeprom.n2415\ : std_logic;
signal \eeprom.n13_adj_329_cascade_\ : std_logic;
signal \eeprom.n2539_cascade_\ : std_logic;
signal \eeprom.n2683\ : std_logic;
signal \eeprom.n2681\ : std_logic;
signal \eeprom.n2713\ : std_logic;
signal \eeprom.n2713_cascade_\ : std_logic;
signal \eeprom.n2715\ : std_logic;
signal \eeprom.n2612\ : std_logic;
signal \eeprom.n2611\ : std_logic;
signal \eeprom.n2612_cascade_\ : std_logic;
signal \eeprom.n2610\ : std_logic;
signal \eeprom.n16_adj_334\ : std_logic;
signal \eeprom.n2618\ : std_logic;
signal \eeprom.n12_adj_333\ : std_logic;
signal \eeprom.n2606\ : std_logic;
signal \eeprom.n2606_cascade_\ : std_logic;
signal \eeprom.n10_adj_332\ : std_logic;
signal \eeprom.n2718\ : std_logic;
signal \eeprom.n5213\ : std_logic;
signal \eeprom.n5215\ : std_logic;
signal \eeprom.n4830\ : std_logic;
signal \eeprom.n2682\ : std_logic;
signal \eeprom.n2714\ : std_logic;
signal \eeprom.n2609\ : std_logic;
signal \eeprom.n3319\ : std_logic;
signal \eeprom.n2608\ : std_logic;
signal \eeprom.n2607\ : std_logic;
signal \eeprom.n2674\ : std_logic;
signal \eeprom.n2607_cascade_\ : std_logic;
signal \eeprom.n2638\ : std_logic;
signal \eeprom.n2706\ : std_logic;
signal \eeprom.n2719\ : std_logic;
signal \eeprom.n2919\ : std_logic;
signal \eeprom.n2419\ : std_logic;
signal \eeprom.n3119\ : std_logic;
signal \eeprom.n2186\ : std_logic;
signal \bfn_24_17_0_\ : std_logic;
signal \eeprom.n2118\ : std_logic;
signal \eeprom.n2185\ : std_logic;
signal \eeprom.n3988\ : std_logic;
signal \eeprom.n2117\ : std_logic;
signal \eeprom.n2184\ : std_logic;
signal \eeprom.n3989\ : std_logic;
signal \eeprom.n2116\ : std_logic;
signal \eeprom.n2183\ : std_logic;
signal \eeprom.n3990\ : std_logic;
signal \eeprom.n2182\ : std_logic;
signal \eeprom.n3991\ : std_logic;
signal \eeprom.n2114\ : std_logic;
signal \eeprom.n2181\ : std_logic;
signal \eeprom.n3992\ : std_logic;
signal \eeprom.n2180\ : std_logic;
signal \eeprom.n3993\ : std_logic;
signal \eeprom.n2112\ : std_logic;
signal \eeprom.n2179\ : std_logic;
signal \eeprom.n3994\ : std_logic;
signal \eeprom.n3995\ : std_logic;
signal \eeprom.n2178\ : std_logic;
signal \bfn_24_18_0_\ : std_logic;
signal \eeprom.n2110\ : std_logic;
signal \eeprom.n2143\ : std_logic;
signal \eeprom.n3996\ : std_logic;
signal \eeprom.n2209\ : std_logic;
signal \eeprom.n3724\ : std_logic;
signal \eeprom.n2015\ : std_logic;
signal \eeprom.n2079\ : std_logic;
signal \eeprom.n2111\ : std_logic;
signal \eeprom.n2018\ : std_logic;
signal \eeprom.n1945_cascade_\ : std_logic;
signal \eeprom.n2017\ : std_logic;
signal \eeprom.n2014\ : std_logic;
signal \eeprom.n2016\ : std_logic;
signal \eeprom.n2083\ : std_logic;
signal \eeprom.n2016_cascade_\ : std_logic;
signal \eeprom.n2044\ : std_logic;
signal \eeprom.n2115\ : std_logic;
signal \eeprom.n2115_cascade_\ : std_logic;
signal \eeprom.n2113\ : std_logic;
signal \eeprom.n5059\ : std_logic;
signal \eeprom.n2013\ : std_logic;
signal \eeprom.n2012\ : std_logic;
signal \eeprom.n1986\ : std_logic;
signal \bfn_24_20_0_\ : std_logic;
signal \eeprom.n1985\ : std_logic;
signal \eeprom.n3973\ : std_logic;
signal \eeprom.n1984\ : std_logic;
signal \eeprom.n3974\ : std_logic;
signal \eeprom.n1983\ : std_logic;
signal \eeprom.n3975\ : std_logic;
signal \eeprom.n1982\ : std_logic;
signal \eeprom.n3976\ : std_logic;
signal \eeprom.n1981\ : std_logic;
signal \eeprom.n3977\ : std_logic;
signal \eeprom.n1980\ : std_logic;
signal \eeprom.n3978\ : std_logic;
signal \eeprom.n1945\ : std_logic;
signal \eeprom.n3979\ : std_logic;
signal \eeprom.n2011\ : std_logic;
signal \eeprom.n2411\ : std_logic;
signal \eeprom.n2478\ : std_logic;
signal \eeprom.n2440\ : std_logic;
signal \eeprom.n3419\ : std_logic;
signal \eeprom.n5169_cascade_\ : std_logic;
signal \eeprom.n5173_cascade_\ : std_logic;
signal \eeprom.n11_adj_328\ : std_logic;
signal \eeprom.n2615\ : std_logic;
signal \eeprom.n2615_cascade_\ : std_logic;
signal \eeprom.n2613\ : std_logic;
signal \eeprom.n2617\ : std_logic;
signal \eeprom.n2614\ : std_logic;
signal \eeprom.n5101_cascade_\ : std_logic;
signal \eeprom.n2616\ : std_logic;
signal \eeprom.n5105\ : std_logic;
signal \eeprom.n2586\ : std_logic;
signal \bfn_24_23_0_\ : std_logic;
signal \eeprom.n2518\ : std_logic;
signal \eeprom.n2585\ : std_logic;
signal \eeprom.n4030\ : std_logic;
signal \eeprom.n2517\ : std_logic;
signal \eeprom.n2584\ : std_logic;
signal \eeprom.n4031\ : std_logic;
signal \eeprom.n2516\ : std_logic;
signal \eeprom.n2583\ : std_logic;
signal \eeprom.n4032\ : std_logic;
signal \eeprom.n2515\ : std_logic;
signal \eeprom.n2582\ : std_logic;
signal \eeprom.n4033\ : std_logic;
signal \eeprom.n2514\ : std_logic;
signal \eeprom.n2581\ : std_logic;
signal \eeprom.n4034\ : std_logic;
signal \eeprom.n2513\ : std_logic;
signal \eeprom.n2580\ : std_logic;
signal \eeprom.n4035\ : std_logic;
signal \eeprom.n2512\ : std_logic;
signal \eeprom.n2579\ : std_logic;
signal \eeprom.n4036\ : std_logic;
signal \eeprom.n4037\ : std_logic;
signal \eeprom.n2511\ : std_logic;
signal \eeprom.n2578\ : std_logic;
signal \bfn_24_24_0_\ : std_logic;
signal \eeprom.n2510\ : std_logic;
signal \eeprom.n2577\ : std_logic;
signal \eeprom.n4038\ : std_logic;
signal \eeprom.n2509\ : std_logic;
signal \eeprom.n2576\ : std_logic;
signal \eeprom.n4039\ : std_logic;
signal \eeprom.n2508\ : std_logic;
signal \eeprom.n2575\ : std_logic;
signal \eeprom.n4040\ : std_logic;
signal \eeprom.n2507\ : std_logic;
signal \eeprom.n2574\ : std_logic;
signal \eeprom.n4041\ : std_logic;
signal \eeprom.n2539\ : std_logic;
signal \eeprom.n2506\ : std_logic;
signal \eeprom.n4042\ : std_logic;
signal \eeprom.n2605\ : std_logic;
signal \eeprom.n2519\ : std_logic;
signal \eeprom.n2619\ : std_logic;
signal \eeprom.n2819\ : std_logic;
signal \eeprom.n3219\ : std_logic;
signal \eeprom.n3019\ : std_logic;
signal \n1805_cascade_\ : std_logic;
signal n170 : std_logic;
signal \n1800_cascade_\ : std_logic;
signal n164 : std_logic;
signal n4_adj_361 : std_logic;
signal \n4_adj_361_cascade_\ : std_logic;
signal n162 : std_logic;
signal \n5361_cascade_\ : std_logic;
signal n172 : std_logic;
signal \n22_adj_367_cascade_\ : std_logic;
signal \n4_adj_369_cascade_\ : std_logic;
signal \n4_cascade_\ : std_logic;
signal n166 : std_logic;
signal n4 : std_logic;
signal n168 : std_logic;
signal n1805 : std_logic;
signal n158 : std_logic;
signal n8 : std_logic;
signal \n5461_cascade_\ : std_logic;
signal n1800 : std_logic;
signal n3585 : std_logic;
signal n160 : std_logic;
signal \eeprom.n2119\ : std_logic;
signal \eeprom.n2319\ : std_logic;
signal \bfn_26_21_0_\ : std_logic;
signal \eeprom.n3931\ : std_logic;
signal \eeprom.eeprom_counter_2\ : std_logic;
signal \eeprom.n3932\ : std_logic;
signal \eeprom.n3933\ : std_logic;
signal \eeprom.eeprom_counter_4\ : std_logic;
signal \eeprom.n3934\ : std_logic;
signal \eeprom.n3935\ : std_logic;
signal \eeprom.n3936\ : std_logic;
signal \eeprom.n3937\ : std_logic;
signal \eeprom.n3938\ : std_logic;
signal \bfn_26_22_0_\ : std_logic;
signal \eeprom.n3939\ : std_logic;
signal \eeprom.n3940\ : std_logic;
signal \eeprom.n3941\ : std_logic;
signal \eeprom.n3942\ : std_logic;
signal \eeprom.eeprom_counter_13\ : std_logic;
signal \eeprom.n3943\ : std_logic;
signal \eeprom.n3944\ : std_logic;
signal \eeprom.n3945\ : std_logic;
signal \eeprom.n3946\ : std_logic;
signal \bfn_26_23_0_\ : std_logic;
signal \eeprom.n3947\ : std_logic;
signal \eeprom.n3948\ : std_logic;
signal \eeprom.n3949\ : std_logic;
signal \eeprom.eeprom_counter_20\ : std_logic;
signal \eeprom.n3950\ : std_logic;
signal \eeprom.n3951\ : std_logic;
signal \eeprom.n3952\ : std_logic;
signal \eeprom.n3953\ : std_logic;
signal \eeprom.n3954\ : std_logic;
signal \bfn_26_24_0_\ : std_logic;
signal \eeprom.n3955\ : std_logic;
signal \eeprom.n3956\ : std_logic;
signal \eeprom.n3957\ : std_logic;
signal \eeprom.n3958\ : std_logic;
signal \eeprom.n3959\ : std_logic;
signal \eeprom.n3960\ : std_logic;
signal \eeprom.n3961\ : std_logic;
signal \eeprom.eeprom_counter_23\ : std_logic;
signal \eeprom.eeprom_counter_16\ : std_logic;
signal \eeprom.n1919\ : std_logic;
signal \eeprom.eeprom_counter_24\ : std_logic;
signal \eeprom.eeprom_counter_18\ : std_logic;
signal \eeprom.eeprom_counter_17\ : std_logic;
signal \eeprom.eeprom_counter_22\ : std_logic;
signal \eeprom.eeprom_counter_21\ : std_logic;
signal \bfn_27_17_0_\ : std_logic;
signal \eeprom.i2c.n3899\ : std_logic;
signal \eeprom.i2c.n3900\ : std_logic;
signal \eeprom.i2c.n3901\ : std_logic;
signal \eeprom.i2c.n3902\ : std_logic;
signal \eeprom.i2c.n3903\ : std_logic;
signal \eeprom.i2c.n3904\ : std_logic;
signal \eeprom.i2c.n3905\ : std_logic;
signal n11 : std_logic;
signal n10_adj_360 : std_logic;
signal n4733 : std_logic;
signal \eeprom.i2c.n1913\ : std_logic;
signal \eeprom.i2c.n534\ : std_logic;
signal \eeprom.i2c.n1829\ : std_logic;
signal \eeprom.i2c.n9\ : std_logic;
signal \eeprom.i2c.n9_cascade_\ : std_logic;
signal n1814 : std_logic;
signal \n1814_cascade_\ : std_logic;
signal \eeprom.i2c.n37\ : std_logic;
signal \eeprom.i2c.n37_cascade_\ : std_logic;
signal \eeprom.i2c.n33\ : std_logic;
signal \eeprom.i2c.n39_cascade_\ : std_logic;
signal \eeprom.i2c.n39\ : std_logic;
signal \eeprom.i2c.n407_cascade_\ : std_logic;
signal \eeprom.n917\ : std_logic;
signal \eeprom.eeprom_counter_5\ : std_logic;
signal \eeprom.n3722\ : std_logic;
signal \eeprom.eeprom_counter_30\ : std_logic;
signal \eeprom.n1256_cascade_\ : std_logic;
signal \eeprom.n1913\ : std_logic;
signal \eeprom.i2c.n13\ : std_logic;
signal \eeprom.eeprom_counter_7\ : std_logic;
signal \INVeeprom.i2c.i2c_scl_enable_124C_net\ : std_logic;
signal \eeprom.n1918\ : std_logic;
signal \eeprom.eeprom_counter_0\ : std_logic;
signal \eeprom.n1912\ : std_logic;
signal \eeprom.eeprom_counter_27\ : std_logic;
signal \eeprom.n1139_cascade_\ : std_logic;
signal \eeprom.eeprom_counter_3\ : std_logic;
signal \eeprom.n1916\ : std_logic;
signal \eeprom.n5035_cascade_\ : std_logic;
signal \eeprom.n5039\ : std_logic;
signal \eeprom.eeprom_counter_12\ : std_logic;
signal \eeprom.eeprom_counter_1\ : std_logic;
signal \eeprom.n892_cascade_\ : std_logic;
signal \eeprom.eeprom_counter_10\ : std_logic;
signal \eeprom.eeprom_counter_28\ : std_logic;
signal \eeprom.n1138_cascade_\ : std_logic;
signal \eeprom.n33_adj_289\ : std_logic;
signal \eeprom.n33\ : std_logic;
signal \bfn_27_23_0_\ : std_logic;
signal \eeprom.n32_adj_288\ : std_logic;
signal \eeprom.n32_adj_287\ : std_logic;
signal \eeprom.n4242\ : std_logic;
signal \eeprom.n31_adj_286\ : std_logic;
signal \eeprom.n31_adj_285\ : std_logic;
signal \eeprom.n4243\ : std_logic;
signal \eeprom.n30_adj_277\ : std_logic;
signal \eeprom.n30_adj_284\ : std_logic;
signal \eeprom.n4244\ : std_logic;
signal \eeprom.n29_adj_278\ : std_logic;
signal \eeprom.n29_adj_283\ : std_logic;
signal \eeprom.n4245\ : std_logic;
signal \eeprom.n28_adj_279\ : std_logic;
signal \eeprom.n28_adj_282\ : std_logic;
signal \eeprom.n4246\ : std_logic;
signal \eeprom.n27_adj_280\ : std_logic;
signal \eeprom.n4247\ : std_logic;
signal \eeprom.n26_adj_276\ : std_logic;
signal \eeprom.n26_adj_275\ : std_logic;
signal \eeprom.n4248\ : std_logic;
signal \eeprom.n4249\ : std_logic;
signal \bfn_27_24_0_\ : std_logic;
signal \eeprom.n24_adj_269\ : std_logic;
signal \eeprom.n4250\ : std_logic;
signal \eeprom.n23_adj_268\ : std_logic;
signal \eeprom.n23\ : std_logic;
signal \eeprom.n4251\ : std_logic;
signal \eeprom.n22_adj_265\ : std_logic;
signal \eeprom.n4252\ : std_logic;
signal \eeprom.n21_adj_264\ : std_logic;
signal \eeprom.n21\ : std_logic;
signal \eeprom.n4253\ : std_logic;
signal \eeprom.n20_adj_259\ : std_logic;
signal \eeprom.n20\ : std_logic;
signal \eeprom.n4254\ : std_logic;
signal \eeprom.n19_adj_320\ : std_logic;
signal \eeprom.n4255\ : std_logic;
signal \eeprom.n18_adj_326\ : std_logic;
signal \eeprom.n4256\ : std_logic;
signal \eeprom.n4257\ : std_logic;
signal \eeprom.n17\ : std_logic;
signal \eeprom.n17_adj_324\ : std_logic;
signal \bfn_27_25_0_\ : std_logic;
signal \eeprom.n16_adj_294\ : std_logic;
signal \eeprom.n16_adj_325\ : std_logic;
signal \eeprom.n4258\ : std_logic;
signal \eeprom.n15_adj_295\ : std_logic;
signal \eeprom.n15\ : std_logic;
signal \eeprom.n4259\ : std_logic;
signal \eeprom.n14\ : std_logic;
signal \eeprom.n4260\ : std_logic;
signal \eeprom.n13\ : std_logic;
signal \eeprom.n13_adj_318\ : std_logic;
signal \eeprom.n4261\ : std_logic;
signal \eeprom.n12_adj_298\ : std_logic;
signal \eeprom.n12_adj_319\ : std_logic;
signal \eeprom.n4262\ : std_logic;
signal \eeprom.n11_adj_299\ : std_logic;
signal \eeprom.n11\ : std_logic;
signal \eeprom.n4263\ : std_logic;
signal \eeprom.n10\ : std_logic;
signal \eeprom.n10_adj_343\ : std_logic;
signal \eeprom.n4264\ : std_logic;
signal \eeprom.n4265\ : std_logic;
signal \eeprom.n9\ : std_logic;
signal \eeprom.n9_adj_308\ : std_logic;
signal \bfn_27_26_0_\ : std_logic;
signal \eeprom.n8_adj_311\ : std_logic;
signal \eeprom.n4266\ : std_logic;
signal \eeprom.n7\ : std_logic;
signal \eeprom.n4267\ : std_logic;
signal \eeprom.n6\ : std_logic;
signal \eeprom.n6_adj_306\ : std_logic;
signal \eeprom.n4268\ : std_logic;
signal \eeprom.n5\ : std_logic;
signal \eeprom.n5_adj_317\ : std_logic;
signal \eeprom.n4269\ : std_logic;
signal \eeprom.n4\ : std_logic;
signal \eeprom.n4270\ : std_logic;
signal \eeprom.n3\ : std_logic;
signal \eeprom.n3_adj_312\ : std_logic;
signal \eeprom.n4271\ : std_logic;
signal \eeprom.n2\ : std_logic;
signal \eeprom.n4272\ : std_logic;
signal \eeprom.i2c.counter_3\ : std_logic;
signal \eeprom.i2c.counter_5\ : std_logic;
signal \eeprom.i2c.counter_4\ : std_logic;
signal \eeprom.i2c.counter_7\ : std_logic;
signal \eeprom.i2c.counter_6\ : std_logic;
signal \eeprom.i2c.n12_cascade_\ : std_logic;
signal \eeprom.i2c.n464\ : std_logic;
signal n4_adj_358 : std_logic;
signal \n10_cascade_\ : std_logic;
signal \state_7_N_162_3\ : std_logic;
signal \eeprom.i2c.n4579\ : std_logic;
signal n11_adj_359 : std_logic;
signal n5458 : std_logic;
signal \n6_adj_365_cascade_\ : std_logic;
signal n471 : std_logic;
signal state_3 : std_logic;
signal n3587 : std_logic;
signal \n3587_cascade_\ : std_logic;
signal n10 : std_logic;
signal n5454 : std_logic;
signal \eeprom.i2c.counter_1\ : std_logic;
signal \eeprom.i2c.counter_2\ : std_logic;
signal \eeprom.i2c.counter_0\ : std_logic;
signal \eeprom.i2c.n5464_cascade_\ : std_logic;
signal \eeprom.i2c.n5451_cascade_\ : std_logic;
signal \eeprom.i2c.sda_out\ : std_logic;
signal \INVeeprom.i2c.sda_out_133C_net\ : std_logic;
signal \eeprom.i2c.n4513\ : std_logic;
signal state_2 : std_logic;
signal n3595 : std_logic;
signal state_1 : std_logic;
signal n3581 : std_logic;
signal \eeprom.i2c.n407\ : std_logic;
signal state_0 : std_logic;
signal sda_enable : std_logic;
signal \INVeeprom.i2c.write_enable_132C_net\ : std_logic;
signal \eeprom.i2c.n524\ : std_logic;
signal \eeprom.i2c.n1901\ : std_logic;
signal \eeprom.n892\ : std_logic;
signal \eeprom.n1198\ : std_logic;
signal \bfn_28_21_0_\ : std_logic;
signal \eeprom.n4273\ : std_logic;
signal \eeprom.n1139\ : std_logic;
signal \eeprom.n1196\ : std_logic;
signal \eeprom.n4274\ : std_logic;
signal \eeprom.n4275\ : std_logic;
signal \eeprom.n4276\ : std_logic;
signal \eeprom.n5327\ : std_logic;
signal \eeprom.n5328\ : std_logic;
signal \eeprom.n4277\ : std_logic;
signal \eeprom.n4278\ : std_logic;
signal \eeprom.n1192\ : std_logic;
signal \eeprom.n1256\ : std_logic;
signal \eeprom.n1843_cascade_\ : std_logic;
signal \eeprom.n1195\ : std_logic;
signal \eeprom.n1915\ : std_logic;
signal \eeprom.eeprom_counter_29\ : std_logic;
signal \eeprom.n4_adj_310\ : std_logic;
signal \eeprom.n1138\ : std_logic;
signal \eeprom.n1137_cascade_\ : std_logic;
signal \eeprom.n4977\ : std_logic;
signal \eeprom.n4983\ : std_logic;
signal \eeprom.n1197\ : std_logic;
signal \eeprom.n1917\ : std_logic;
signal \eeprom.n1194\ : std_logic;
signal \eeprom.n1137\ : std_logic;
signal \eeprom.n1843\ : std_logic;
signal \eeprom.n1914\ : std_logic;
signal \eeprom.eeprom_counter_14\ : std_logic;
signal \eeprom.n19\ : std_logic;
signal \eeprom.n25_adj_271\ : std_logic;
signal \eeprom.n3519\ : std_logic;
signal \eeprom.n27_adj_281\ : std_logic;
signal \eeprom.eeprom_counter_6\ : std_logic;
signal \eeprom.n3719\ : std_logic;
signal \eeprom.eeprom_counter_19\ : std_logic;
signal \eeprom.n14_adj_297\ : std_logic;
signal \eeprom.eeprom_counter_26\ : std_logic;
signal \eeprom.n7_adj_309\ : std_logic;
signal \eeprom.n1140\ : std_logic;
signal \eeprom.eeprom_counter_8\ : std_logic;
signal \eeprom.n25_adj_272\ : std_logic;
signal \eeprom.eeprom_counter_31\ : std_logic;
signal \eeprom.n2_adj_307\ : std_logic;
signal \eeprom.n1135\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n174 : std_logic;
signal rw : std_logic;
signal saved_addr_0 : std_logic;
signal \state_7_N_146_0\ : std_logic;
signal \eeprom.enable\ : std_logic;
signal \eeprom.i2c.n1832\ : std_logic;
signal \eeprom.i2c.n6_adj_255_cascade_\ : std_logic;
signal \eeprom.eeprom_counter_9\ : std_logic;
signal \eeprom.n24_adj_270\ : std_logic;
signal \eeprom.i2c.i2c_clk\ : std_logic;
signal scl_enable : std_logic;
signal scl_c : std_logic;
signal \eeprom.eeprom_counter_11\ : std_logic;
signal \eeprom.n22_adj_266\ : std_logic;
signal \eeprom.eeprom_counter_25\ : std_logic;
signal \eeprom.n8\ : std_logic;
signal \eeprom.eeprom_counter_15\ : std_logic;
signal \eeprom.n18_adj_293\ : std_logic;
signal \eeprom.i2c.counter2_0\ : std_logic;
signal \bfn_30_20_0_\ : std_logic;
signal \eeprom.i2c.counter2_1\ : std_logic;
signal \eeprom.i2c.n3962\ : std_logic;
signal \eeprom.i2c.counter2_2\ : std_logic;
signal \eeprom.i2c.n3963\ : std_logic;
signal \eeprom.i2c.counter2_3\ : std_logic;
signal \eeprom.i2c.n3964\ : std_logic;
signal \eeprom.i2c.n3965\ : std_logic;
signal \eeprom.i2c.counter2_4\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK_N\ : std_logic;
signal \eeprom.i2c.counter2_7__N_133\ : std_logic;

signal \CS_CLK_wire\ : std_logic;
signal \CS_wire\ : std_logic;
signal \DE_wire\ : std_logic;
signal \INHA_wire\ : std_logic;
signal \INHB_wire\ : std_logic;
signal \INHC_wire\ : std_logic;
signal \INLA_wire\ : std_logic;
signal \INLB_wire\ : std_logic;
signal \INLC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \NEOPXL_wire\ : std_logic;
signal \TX_wire\ : std_logic;
signal \USBPU_wire\ : std_logic;
signal \CLK_wire\ : std_logic;

begin
    CS_CLK <= \CS_CLK_wire\;
    CS <= \CS_wire\;
    DE <= \DE_wire\;
    INHA <= \INHA_wire\;
    INHB <= \INHB_wire\;
    INHC <= \INHC_wire\;
    INLA <= \INLA_wire\;
    INLB <= \INLB_wire\;
    INLC <= \INLC_wire\;
    LED <= \LED_wire\;
    NEOPXL <= \NEOPXL_wire\;
    TX <= \TX_wire\;
    USBPU <= \USBPU_wire\;
    \CLK_wire\ <= CLK;

    \CS_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30138\,
            DIN => \N__30137\,
            DOUT => \N__30136\,
            PACKAGEPIN => \CS_CLK_wire\
        );

    \CS_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30138\,
            PADOUT => \N__30137\,
            PADIN => \N__30136\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \CS_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30129\,
            DIN => \N__30128\,
            DOUT => \N__30127\,
            PACKAGEPIN => \CS_wire\
        );

    \CS_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30129\,
            PADOUT => \N__30128\,
            PADIN => \N__30127\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \DE_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30120\,
            DIN => \N__30119\,
            DOUT => \N__30118\,
            PACKAGEPIN => \DE_wire\
        );

    \DE_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30120\,
            PADOUT => \N__30119\,
            PADIN => \N__30118\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30111\,
            DIN => \N__30110\,
            DOUT => \N__30109\,
            PACKAGEPIN => \INHA_wire\
        );

    \INHA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30111\,
            PADOUT => \N__30110\,
            PADIN => \N__30109\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30102\,
            DIN => \N__30101\,
            DOUT => \N__30100\,
            PACKAGEPIN => \INHB_wire\
        );

    \INHB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30102\,
            PADOUT => \N__30101\,
            PADIN => \N__30100\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INHC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30093\,
            DIN => \N__30092\,
            DOUT => \N__30091\,
            PACKAGEPIN => \INHC_wire\
        );

    \INHC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30093\,
            PADOUT => \N__30092\,
            PADIN => \N__30091\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLA_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30084\,
            DIN => \N__30083\,
            DOUT => \N__30082\,
            PACKAGEPIN => \INLA_wire\
        );

    \INLA_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30084\,
            PADOUT => \N__30083\,
            PADIN => \N__30082\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLB_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30075\,
            DIN => \N__30074\,
            DOUT => \N__30073\,
            PACKAGEPIN => \INLB_wire\
        );

    \INLB_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30075\,
            PADOUT => \N__30074\,
            PADIN => \N__30073\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \INLC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30066\,
            DIN => \N__30065\,
            DOUT => \N__30064\,
            PACKAGEPIN => \INLC_wire\
        );

    \INLC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30066\,
            PADOUT => \N__30065\,
            PADIN => \N__30064\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30057\,
            DIN => \N__30056\,
            DOUT => \N__30055\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30057\,
            PADOUT => \N__30056\,
            PADIN => \N__30055\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__11906\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \NEOPXL_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30048\,
            DIN => \N__30047\,
            DOUT => \N__30046\,
            PACKAGEPIN => \NEOPXL_wire\
        );

    \NEOPXL_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30048\,
            PADOUT => \N__30047\,
            PADIN => \N__30046\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \TX_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30039\,
            DIN => \N__30038\,
            DOUT => \N__30037\,
            PACKAGEPIN => \TX_wire\
        );

    \TX_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30039\,
            PADOUT => \N__30038\,
            PADIN => \N__30037\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \USBPU_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30030\,
            DIN => \N__30029\,
            DOUT => \N__30028\,
            PACKAGEPIN => \USBPU_wire\
        );

    \USBPU_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30030\,
            PADOUT => \N__30029\,
            PADIN => \N__30028\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \scl_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__30021\,
            DIN => \N__30020\,
            DOUT => \N__30019\,
            PACKAGEPIN => SCL
        );

    \scl_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30021\,
            PADOUT => \N__30020\,
            PADIN => \N__30019\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__29558\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__29585\
        );

    \sda_output_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__30012\,
            DIN => \N__30011\,
            DOUT => \N__30010\,
            PACKAGEPIN => SDA
        );

    \sda_output_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30012\,
            PADOUT => \N__30011\,
            PADIN => \N__30010\,
            CLOCKENABLE => 'H',
            DIN0 => OPEN,
            DIN1 => OPEN,
            DOUT0 => \N__26531\,
            DOUT1 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => \N__27311\
        );

    \CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__30003\,
            DIN => \N__30002\,
            DOUT => \N__30001\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__30003\,
            PADOUT => \N__30002\,
            PADIN => \N__30001\,
            CLOCKENABLE => 'H',
            DIN0 => \CLK_pad_gb_input\,
            DIN1 => OPEN,
            DOUT0 => '0',
            DOUT1 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0'
        );

    \I__7050\ : InMux
    port map (
            O => \N__29984\,
            I => \N__29980\
        );

    \I__7049\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29977\
        );

    \I__7048\ : LocalMux
    port map (
            O => \N__29980\,
            I => \N__29973\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__29977\,
            I => \N__29970\
        );

    \I__7046\ : InMux
    port map (
            O => \N__29976\,
            I => \N__29967\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__29973\,
            I => \N__29962\
        );

    \I__7044\ : Span4Mux_h
    port map (
            O => \N__29970\,
            I => \N__29962\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__29967\,
            I => \eeprom.eeprom_counter_15\
        );

    \I__7042\ : Odrv4
    port map (
            O => \N__29962\,
            I => \eeprom.eeprom_counter_15\
        );

    \I__7041\ : CascadeMux
    port map (
            O => \N__29957\,
            I => \N__29954\
        );

    \I__7040\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29951\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__29951\,
            I => \N__29948\
        );

    \I__7038\ : Span4Mux_v
    port map (
            O => \N__29948\,
            I => \N__29945\
        );

    \I__7037\ : Odrv4
    port map (
            O => \N__29945\,
            I => \eeprom.n18_adj_293\
        );

    \I__7036\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29938\
        );

    \I__7035\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29935\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__29938\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__7033\ : LocalMux
    port map (
            O => \N__29935\,
            I => \eeprom.i2c.counter2_0\
        );

    \I__7032\ : InMux
    port map (
            O => \N__29930\,
            I => \bfn_30_20_0_\
        );

    \I__7031\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29923\
        );

    \I__7030\ : InMux
    port map (
            O => \N__29926\,
            I => \N__29920\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__29923\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__29920\,
            I => \eeprom.i2c.counter2_1\
        );

    \I__7027\ : InMux
    port map (
            O => \N__29915\,
            I => \eeprom.i2c.n3962\
        );

    \I__7026\ : InMux
    port map (
            O => \N__29912\,
            I => \N__29908\
        );

    \I__7025\ : InMux
    port map (
            O => \N__29911\,
            I => \N__29905\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__29908\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__29905\,
            I => \eeprom.i2c.counter2_2\
        );

    \I__7022\ : InMux
    port map (
            O => \N__29900\,
            I => \eeprom.i2c.n3963\
        );

    \I__7021\ : InMux
    port map (
            O => \N__29897\,
            I => \N__29893\
        );

    \I__7020\ : InMux
    port map (
            O => \N__29896\,
            I => \N__29890\
        );

    \I__7019\ : LocalMux
    port map (
            O => \N__29893\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__7018\ : LocalMux
    port map (
            O => \N__29890\,
            I => \eeprom.i2c.counter2_3\
        );

    \I__7017\ : InMux
    port map (
            O => \N__29885\,
            I => \eeprom.i2c.n3964\
        );

    \I__7016\ : InMux
    port map (
            O => \N__29882\,
            I => \eeprom.i2c.n3965\
        );

    \I__7015\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29875\
        );

    \I__7014\ : InMux
    port map (
            O => \N__29878\,
            I => \N__29872\
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__29875\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__7012\ : LocalMux
    port map (
            O => \N__29872\,
            I => \eeprom.i2c.counter2_4\
        );

    \I__7011\ : ClkMux
    port map (
            O => \N__29867\,
            I => \N__29831\
        );

    \I__7010\ : ClkMux
    port map (
            O => \N__29866\,
            I => \N__29831\
        );

    \I__7009\ : ClkMux
    port map (
            O => \N__29865\,
            I => \N__29831\
        );

    \I__7008\ : ClkMux
    port map (
            O => \N__29864\,
            I => \N__29831\
        );

    \I__7007\ : ClkMux
    port map (
            O => \N__29863\,
            I => \N__29831\
        );

    \I__7006\ : ClkMux
    port map (
            O => \N__29862\,
            I => \N__29831\
        );

    \I__7005\ : ClkMux
    port map (
            O => \N__29861\,
            I => \N__29831\
        );

    \I__7004\ : ClkMux
    port map (
            O => \N__29860\,
            I => \N__29831\
        );

    \I__7003\ : ClkMux
    port map (
            O => \N__29859\,
            I => \N__29831\
        );

    \I__7002\ : ClkMux
    port map (
            O => \N__29858\,
            I => \N__29831\
        );

    \I__7001\ : ClkMux
    port map (
            O => \N__29857\,
            I => \N__29831\
        );

    \I__7000\ : ClkMux
    port map (
            O => \N__29856\,
            I => \N__29831\
        );

    \I__6999\ : GlobalMux
    port map (
            O => \N__29831\,
            I => \N__29828\
        );

    \I__6998\ : gio2CtrlBuf
    port map (
            O => \N__29828\,
            I => \CLK_N\
        );

    \I__6997\ : SRMux
    port map (
            O => \N__29825\,
            I => \N__29821\
        );

    \I__6996\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29818\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__29821\,
            I => \N__29813\
        );

    \I__6994\ : LocalMux
    port map (
            O => \N__29818\,
            I => \N__29810\
        );

    \I__6993\ : InMux
    port map (
            O => \N__29817\,
            I => \N__29805\
        );

    \I__6992\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29805\
        );

    \I__6991\ : Odrv4
    port map (
            O => \N__29813\,
            I => \eeprom.i2c.counter2_7__N_133\
        );

    \I__6990\ : Odrv4
    port map (
            O => \N__29810\,
            I => \eeprom.i2c.counter2_7__N_133\
        );

    \I__6989\ : LocalMux
    port map (
            O => \N__29805\,
            I => \eeprom.i2c.counter2_7__N_133\
        );

    \I__6988\ : InMux
    port map (
            O => \N__29798\,
            I => \N__29794\
        );

    \I__6987\ : InMux
    port map (
            O => \N__29797\,
            I => \N__29791\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__29794\,
            I => \state_7_N_146_0\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__29791\,
            I => \state_7_N_146_0\
        );

    \I__6984\ : SRMux
    port map (
            O => \N__29786\,
            I => \N__29782\
        );

    \I__6983\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29778\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__29782\,
            I => \N__29775\
        );

    \I__6981\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29772\
        );

    \I__6980\ : LocalMux
    port map (
            O => \N__29778\,
            I => \N__29769\
        );

    \I__6979\ : Span4Mux_v
    port map (
            O => \N__29775\,
            I => \N__29764\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__29772\,
            I => \N__29764\
        );

    \I__6977\ : Span4Mux_v
    port map (
            O => \N__29769\,
            I => \N__29759\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__29764\,
            I => \N__29759\
        );

    \I__6975\ : Span4Mux_h
    port map (
            O => \N__29759\,
            I => \N__29756\
        );

    \I__6974\ : Odrv4
    port map (
            O => \N__29756\,
            I => \eeprom.enable\
        );

    \I__6973\ : CEMux
    port map (
            O => \N__29753\,
            I => \N__29750\
        );

    \I__6972\ : LocalMux
    port map (
            O => \N__29750\,
            I => \N__29747\
        );

    \I__6971\ : Span4Mux_h
    port map (
            O => \N__29747\,
            I => \N__29744\
        );

    \I__6970\ : Odrv4
    port map (
            O => \N__29744\,
            I => \eeprom.i2c.n1832\
        );

    \I__6969\ : CascadeMux
    port map (
            O => \N__29741\,
            I => \eeprom.i2c.n6_adj_255_cascade_\
        );

    \I__6968\ : InMux
    port map (
            O => \N__29738\,
            I => \N__29734\
        );

    \I__6967\ : InMux
    port map (
            O => \N__29737\,
            I => \N__29731\
        );

    \I__6966\ : LocalMux
    port map (
            O => \N__29734\,
            I => \N__29727\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__29731\,
            I => \N__29724\
        );

    \I__6964\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29721\
        );

    \I__6963\ : Span4Mux_v
    port map (
            O => \N__29727\,
            I => \N__29716\
        );

    \I__6962\ : Span4Mux_v
    port map (
            O => \N__29724\,
            I => \N__29716\
        );

    \I__6961\ : LocalMux
    port map (
            O => \N__29721\,
            I => \eeprom.eeprom_counter_9\
        );

    \I__6960\ : Odrv4
    port map (
            O => \N__29716\,
            I => \eeprom.eeprom_counter_9\
        );

    \I__6959\ : CascadeMux
    port map (
            O => \N__29711\,
            I => \N__29708\
        );

    \I__6958\ : InMux
    port map (
            O => \N__29708\,
            I => \N__29705\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29702\
        );

    \I__6956\ : Span4Mux_h
    port map (
            O => \N__29702\,
            I => \N__29699\
        );

    \I__6955\ : Odrv4
    port map (
            O => \N__29699\,
            I => \eeprom.n24_adj_270\
        );

    \I__6954\ : ClkMux
    port map (
            O => \N__29696\,
            I => \N__29690\
        );

    \I__6953\ : ClkMux
    port map (
            O => \N__29695\,
            I => \N__29684\
        );

    \I__6952\ : ClkMux
    port map (
            O => \N__29694\,
            I => \N__29680\
        );

    \I__6951\ : ClkMux
    port map (
            O => \N__29693\,
            I => \N__29677\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__29690\,
            I => \N__29674\
        );

    \I__6949\ : ClkMux
    port map (
            O => \N__29689\,
            I => \N__29671\
        );

    \I__6948\ : ClkMux
    port map (
            O => \N__29688\,
            I => \N__29668\
        );

    \I__6947\ : ClkMux
    port map (
            O => \N__29687\,
            I => \N__29665\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__29684\,
            I => \N__29662\
        );

    \I__6945\ : ClkMux
    port map (
            O => \N__29683\,
            I => \N__29659\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__29680\,
            I => \N__29651\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__29677\,
            I => \N__29651\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__29674\,
            I => \N__29646\
        );

    \I__6941\ : LocalMux
    port map (
            O => \N__29671\,
            I => \N__29646\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29641\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__29665\,
            I => \N__29641\
        );

    \I__6938\ : Span4Mux_h
    port map (
            O => \N__29662\,
            I => \N__29636\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__29659\,
            I => \N__29636\
        );

    \I__6936\ : ClkMux
    port map (
            O => \N__29658\,
            I => \N__29633\
        );

    \I__6935\ : InMux
    port map (
            O => \N__29657\,
            I => \N__29629\
        );

    \I__6934\ : ClkMux
    port map (
            O => \N__29656\,
            I => \N__29626\
        );

    \I__6933\ : Span4Mux_v
    port map (
            O => \N__29651\,
            I => \N__29619\
        );

    \I__6932\ : Span4Mux_v
    port map (
            O => \N__29646\,
            I => \N__29619\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__29641\,
            I => \N__29616\
        );

    \I__6930\ : Span4Mux_v
    port map (
            O => \N__29636\,
            I => \N__29611\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__29633\,
            I => \N__29611\
        );

    \I__6928\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29608\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__29629\,
            I => \N__29603\
        );

    \I__6926\ : LocalMux
    port map (
            O => \N__29626\,
            I => \N__29603\
        );

    \I__6925\ : InMux
    port map (
            O => \N__29625\,
            I => \N__29598\
        );

    \I__6924\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29598\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__29619\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__6922\ : Odrv4
    port map (
            O => \N__29616\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__29611\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__6920\ : LocalMux
    port map (
            O => \N__29608\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__29603\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__29598\,
            I => \eeprom.i2c.i2c_clk\
        );

    \I__6917\ : IoInMux
    port map (
            O => \N__29585\,
            I => \N__29582\
        );

    \I__6916\ : LocalMux
    port map (
            O => \N__29582\,
            I => \N__29579\
        );

    \I__6915\ : IoSpan4Mux
    port map (
            O => \N__29579\,
            I => \N__29575\
        );

    \I__6914\ : InMux
    port map (
            O => \N__29578\,
            I => \N__29572\
        );

    \I__6913\ : Span4Mux_s2_h
    port map (
            O => \N__29575\,
            I => \N__29569\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__29572\,
            I => \N__29566\
        );

    \I__6911\ : Span4Mux_v
    port map (
            O => \N__29569\,
            I => \N__29561\
        );

    \I__6910\ : Span4Mux_v
    port map (
            O => \N__29566\,
            I => \N__29561\
        );

    \I__6909\ : Odrv4
    port map (
            O => \N__29561\,
            I => scl_enable
        );

    \I__6908\ : IoInMux
    port map (
            O => \N__29558\,
            I => \N__29555\
        );

    \I__6907\ : LocalMux
    port map (
            O => \N__29555\,
            I => \N__29552\
        );

    \I__6906\ : Odrv12
    port map (
            O => \N__29552\,
            I => scl_c
        );

    \I__6905\ : InMux
    port map (
            O => \N__29549\,
            I => \N__29546\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__29546\,
            I => \N__29541\
        );

    \I__6903\ : InMux
    port map (
            O => \N__29545\,
            I => \N__29538\
        );

    \I__6902\ : InMux
    port map (
            O => \N__29544\,
            I => \N__29535\
        );

    \I__6901\ : Span4Mux_h
    port map (
            O => \N__29541\,
            I => \N__29532\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__29538\,
            I => \N__29529\
        );

    \I__6899\ : LocalMux
    port map (
            O => \N__29535\,
            I => \eeprom.eeprom_counter_11\
        );

    \I__6898\ : Odrv4
    port map (
            O => \N__29532\,
            I => \eeprom.eeprom_counter_11\
        );

    \I__6897\ : Odrv4
    port map (
            O => \N__29529\,
            I => \eeprom.eeprom_counter_11\
        );

    \I__6896\ : CascadeMux
    port map (
            O => \N__29522\,
            I => \N__29519\
        );

    \I__6895\ : InMux
    port map (
            O => \N__29519\,
            I => \N__29516\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__29516\,
            I => \N__29513\
        );

    \I__6893\ : Span4Mux_h
    port map (
            O => \N__29513\,
            I => \N__29510\
        );

    \I__6892\ : Odrv4
    port map (
            O => \N__29510\,
            I => \eeprom.n22_adj_266\
        );

    \I__6891\ : CascadeMux
    port map (
            O => \N__29507\,
            I => \N__29504\
        );

    \I__6890\ : InMux
    port map (
            O => \N__29504\,
            I => \N__29500\
        );

    \I__6889\ : InMux
    port map (
            O => \N__29503\,
            I => \N__29497\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__29500\,
            I => \N__29491\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__29497\,
            I => \N__29491\
        );

    \I__6886\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29488\
        );

    \I__6885\ : Span4Mux_h
    port map (
            O => \N__29491\,
            I => \N__29485\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__29488\,
            I => \eeprom.eeprom_counter_25\
        );

    \I__6883\ : Odrv4
    port map (
            O => \N__29485\,
            I => \eeprom.eeprom_counter_25\
        );

    \I__6882\ : CascadeMux
    port map (
            O => \N__29480\,
            I => \N__29477\
        );

    \I__6881\ : InMux
    port map (
            O => \N__29477\,
            I => \N__29474\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__29474\,
            I => \N__29471\
        );

    \I__6879\ : Span4Mux_v
    port map (
            O => \N__29471\,
            I => \N__29468\
        );

    \I__6878\ : Odrv4
    port map (
            O => \N__29468\,
            I => \eeprom.n8\
        );

    \I__6877\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29462\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__29462\,
            I => \eeprom.n25_adj_271\
        );

    \I__6875\ : InMux
    port map (
            O => \N__29459\,
            I => \N__29454\
        );

    \I__6874\ : InMux
    port map (
            O => \N__29458\,
            I => \N__29451\
        );

    \I__6873\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29448\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29445\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__29451\,
            I => \N__29442\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__29448\,
            I => \N__29439\
        );

    \I__6869\ : Span4Mux_v
    port map (
            O => \N__29445\,
            I => \N__29436\
        );

    \I__6868\ : Span4Mux_v
    port map (
            O => \N__29442\,
            I => \N__29431\
        );

    \I__6867\ : Span4Mux_h
    port map (
            O => \N__29439\,
            I => \N__29431\
        );

    \I__6866\ : Sp12to4
    port map (
            O => \N__29436\,
            I => \N__29428\
        );

    \I__6865\ : Span4Mux_h
    port map (
            O => \N__29431\,
            I => \N__29425\
        );

    \I__6864\ : Span12Mux_h
    port map (
            O => \N__29428\,
            I => \N__29422\
        );

    \I__6863\ : Span4Mux_h
    port map (
            O => \N__29425\,
            I => \N__29419\
        );

    \I__6862\ : Odrv12
    port map (
            O => \N__29422\,
            I => \eeprom.n3519\
        );

    \I__6861\ : Odrv4
    port map (
            O => \N__29419\,
            I => \eeprom.n3519\
        );

    \I__6860\ : InMux
    port map (
            O => \N__29414\,
            I => \N__29411\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__29411\,
            I => \eeprom.n27_adj_281\
        );

    \I__6858\ : InMux
    port map (
            O => \N__29408\,
            I => \N__29405\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__29405\,
            I => \N__29401\
        );

    \I__6856\ : InMux
    port map (
            O => \N__29404\,
            I => \N__29398\
        );

    \I__6855\ : Span4Mux_h
    port map (
            O => \N__29401\,
            I => \N__29395\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__29398\,
            I => \N__29391\
        );

    \I__6853\ : Span4Mux_v
    port map (
            O => \N__29395\,
            I => \N__29387\
        );

    \I__6852\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29384\
        );

    \I__6851\ : Span4Mux_h
    port map (
            O => \N__29391\,
            I => \N__29381\
        );

    \I__6850\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29378\
        );

    \I__6849\ : Odrv4
    port map (
            O => \N__29387\,
            I => \eeprom.eeprom_counter_6\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__29384\,
            I => \eeprom.eeprom_counter_6\
        );

    \I__6847\ : Odrv4
    port map (
            O => \N__29381\,
            I => \eeprom.eeprom_counter_6\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__29378\,
            I => \eeprom.eeprom_counter_6\
        );

    \I__6845\ : CascadeMux
    port map (
            O => \N__29369\,
            I => \N__29366\
        );

    \I__6844\ : InMux
    port map (
            O => \N__29366\,
            I => \N__29363\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__29363\,
            I => \N__29360\
        );

    \I__6842\ : Span4Mux_h
    port map (
            O => \N__29360\,
            I => \N__29357\
        );

    \I__6841\ : Span4Mux_h
    port map (
            O => \N__29357\,
            I => \N__29354\
        );

    \I__6840\ : Span4Mux_v
    port map (
            O => \N__29354\,
            I => \N__29351\
        );

    \I__6839\ : Odrv4
    port map (
            O => \N__29351\,
            I => \eeprom.n3719\
        );

    \I__6838\ : InMux
    port map (
            O => \N__29348\,
            I => \N__29344\
        );

    \I__6837\ : InMux
    port map (
            O => \N__29347\,
            I => \N__29341\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__29344\,
            I => \N__29337\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__29341\,
            I => \N__29334\
        );

    \I__6834\ : InMux
    port map (
            O => \N__29340\,
            I => \N__29331\
        );

    \I__6833\ : Span4Mux_v
    port map (
            O => \N__29337\,
            I => \N__29328\
        );

    \I__6832\ : Span4Mux_h
    port map (
            O => \N__29334\,
            I => \N__29325\
        );

    \I__6831\ : LocalMux
    port map (
            O => \N__29331\,
            I => \eeprom.eeprom_counter_19\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__29328\,
            I => \eeprom.eeprom_counter_19\
        );

    \I__6829\ : Odrv4
    port map (
            O => \N__29325\,
            I => \eeprom.eeprom_counter_19\
        );

    \I__6828\ : InMux
    port map (
            O => \N__29318\,
            I => \N__29315\
        );

    \I__6827\ : LocalMux
    port map (
            O => \N__29315\,
            I => \eeprom.n14_adj_297\
        );

    \I__6826\ : InMux
    port map (
            O => \N__29312\,
            I => \N__29308\
        );

    \I__6825\ : InMux
    port map (
            O => \N__29311\,
            I => \N__29305\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__29308\,
            I => \N__29299\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__29305\,
            I => \N__29299\
        );

    \I__6822\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29296\
        );

    \I__6821\ : Odrv4
    port map (
            O => \N__29299\,
            I => \eeprom.eeprom_counter_26\
        );

    \I__6820\ : LocalMux
    port map (
            O => \N__29296\,
            I => \eeprom.eeprom_counter_26\
        );

    \I__6819\ : InMux
    port map (
            O => \N__29291\,
            I => \N__29288\
        );

    \I__6818\ : LocalMux
    port map (
            O => \N__29288\,
            I => \N__29284\
        );

    \I__6817\ : InMux
    port map (
            O => \N__29287\,
            I => \N__29281\
        );

    \I__6816\ : Span4Mux_v
    port map (
            O => \N__29284\,
            I => \N__29276\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__29281\,
            I => \N__29276\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__29276\,
            I => \eeprom.n7_adj_309\
        );

    \I__6813\ : CascadeMux
    port map (
            O => \N__29273\,
            I => \N__29269\
        );

    \I__6812\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29266\
        );

    \I__6811\ : InMux
    port map (
            O => \N__29269\,
            I => \N__29263\
        );

    \I__6810\ : LocalMux
    port map (
            O => \N__29266\,
            I => \N__29260\
        );

    \I__6809\ : LocalMux
    port map (
            O => \N__29263\,
            I => \N__29257\
        );

    \I__6808\ : Odrv4
    port map (
            O => \N__29260\,
            I => \eeprom.n1140\
        );

    \I__6807\ : Odrv4
    port map (
            O => \N__29257\,
            I => \eeprom.n1140\
        );

    \I__6806\ : InMux
    port map (
            O => \N__29252\,
            I => \N__29248\
        );

    \I__6805\ : InMux
    port map (
            O => \N__29251\,
            I => \N__29245\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__29248\,
            I => \N__29241\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__29245\,
            I => \N__29238\
        );

    \I__6802\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29235\
        );

    \I__6801\ : Span4Mux_h
    port map (
            O => \N__29241\,
            I => \N__29232\
        );

    \I__6800\ : Span4Mux_h
    port map (
            O => \N__29238\,
            I => \N__29229\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__29235\,
            I => \eeprom.eeprom_counter_8\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__29232\,
            I => \eeprom.eeprom_counter_8\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__29229\,
            I => \eeprom.eeprom_counter_8\
        );

    \I__6796\ : CascadeMux
    port map (
            O => \N__29222\,
            I => \N__29219\
        );

    \I__6795\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29216\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__29216\,
            I => \eeprom.n25_adj_272\
        );

    \I__6793\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29200\
        );

    \I__6792\ : InMux
    port map (
            O => \N__29212\,
            I => \N__29187\
        );

    \I__6791\ : InMux
    port map (
            O => \N__29211\,
            I => \N__29187\
        );

    \I__6790\ : InMux
    port map (
            O => \N__29210\,
            I => \N__29187\
        );

    \I__6789\ : InMux
    port map (
            O => \N__29209\,
            I => \N__29187\
        );

    \I__6788\ : InMux
    port map (
            O => \N__29208\,
            I => \N__29187\
        );

    \I__6787\ : InMux
    port map (
            O => \N__29207\,
            I => \N__29181\
        );

    \I__6786\ : InMux
    port map (
            O => \N__29206\,
            I => \N__29165\
        );

    \I__6785\ : InMux
    port map (
            O => \N__29205\,
            I => \N__29162\
        );

    \I__6784\ : InMux
    port map (
            O => \N__29204\,
            I => \N__29159\
        );

    \I__6783\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29156\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__29200\,
            I => \N__29153\
        );

    \I__6781\ : InMux
    port map (
            O => \N__29199\,
            I => \N__29150\
        );

    \I__6780\ : InMux
    port map (
            O => \N__29198\,
            I => \N__29147\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__29187\,
            I => \N__29144\
        );

    \I__6778\ : InMux
    port map (
            O => \N__29186\,
            I => \N__29141\
        );

    \I__6777\ : InMux
    port map (
            O => \N__29185\,
            I => \N__29138\
        );

    \I__6776\ : CascadeMux
    port map (
            O => \N__29184\,
            I => \N__29134\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__29181\,
            I => \N__29131\
        );

    \I__6774\ : InMux
    port map (
            O => \N__29180\,
            I => \N__29124\
        );

    \I__6773\ : InMux
    port map (
            O => \N__29179\,
            I => \N__29124\
        );

    \I__6772\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29124\
        );

    \I__6771\ : InMux
    port map (
            O => \N__29177\,
            I => \N__29117\
        );

    \I__6770\ : InMux
    port map (
            O => \N__29176\,
            I => \N__29117\
        );

    \I__6769\ : InMux
    port map (
            O => \N__29175\,
            I => \N__29117\
        );

    \I__6768\ : InMux
    port map (
            O => \N__29174\,
            I => \N__29112\
        );

    \I__6767\ : InMux
    port map (
            O => \N__29173\,
            I => \N__29112\
        );

    \I__6766\ : InMux
    port map (
            O => \N__29172\,
            I => \N__29105\
        );

    \I__6765\ : InMux
    port map (
            O => \N__29171\,
            I => \N__29105\
        );

    \I__6764\ : InMux
    port map (
            O => \N__29170\,
            I => \N__29105\
        );

    \I__6763\ : InMux
    port map (
            O => \N__29169\,
            I => \N__29102\
        );

    \I__6762\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29099\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__29165\,
            I => \N__29091\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__29162\,
            I => \N__29087\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__29159\,
            I => \N__29084\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__29156\,
            I => \N__29081\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__29153\,
            I => \N__29072\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__29150\,
            I => \N__29072\
        );

    \I__6755\ : LocalMux
    port map (
            O => \N__29147\,
            I => \N__29072\
        );

    \I__6754\ : Span4Mux_h
    port map (
            O => \N__29144\,
            I => \N__29072\
        );

    \I__6753\ : LocalMux
    port map (
            O => \N__29141\,
            I => \N__29069\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__29138\,
            I => \N__29066\
        );

    \I__6751\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29061\
        );

    \I__6750\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29061\
        );

    \I__6749\ : Span4Mux_v
    port map (
            O => \N__29131\,
            I => \N__29054\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__29124\,
            I => \N__29054\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__29117\,
            I => \N__29054\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__29112\,
            I => \N__29049\
        );

    \I__6745\ : LocalMux
    port map (
            O => \N__29105\,
            I => \N__29049\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__29102\,
            I => \N__29044\
        );

    \I__6743\ : LocalMux
    port map (
            O => \N__29099\,
            I => \N__29044\
        );

    \I__6742\ : InMux
    port map (
            O => \N__29098\,
            I => \N__29037\
        );

    \I__6741\ : InMux
    port map (
            O => \N__29097\,
            I => \N__29037\
        );

    \I__6740\ : InMux
    port map (
            O => \N__29096\,
            I => \N__29037\
        );

    \I__6739\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29034\
        );

    \I__6738\ : InMux
    port map (
            O => \N__29094\,
            I => \N__29031\
        );

    \I__6737\ : Span12Mux_h
    port map (
            O => \N__29091\,
            I => \N__29028\
        );

    \I__6736\ : InMux
    port map (
            O => \N__29090\,
            I => \N__29025\
        );

    \I__6735\ : Span4Mux_v
    port map (
            O => \N__29087\,
            I => \N__29010\
        );

    \I__6734\ : Span4Mux_h
    port map (
            O => \N__29084\,
            I => \N__29010\
        );

    \I__6733\ : Span4Mux_v
    port map (
            O => \N__29081\,
            I => \N__29010\
        );

    \I__6732\ : Span4Mux_v
    port map (
            O => \N__29072\,
            I => \N__29010\
        );

    \I__6731\ : Span4Mux_v
    port map (
            O => \N__29069\,
            I => \N__29010\
        );

    \I__6730\ : Span4Mux_v
    port map (
            O => \N__29066\,
            I => \N__29010\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__29061\,
            I => \N__29010\
        );

    \I__6728\ : Span4Mux_h
    port map (
            O => \N__29054\,
            I => \N__29001\
        );

    \I__6727\ : Span4Mux_v
    port map (
            O => \N__29049\,
            I => \N__29001\
        );

    \I__6726\ : Span4Mux_h
    port map (
            O => \N__29044\,
            I => \N__29001\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__29037\,
            I => \N__29001\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__29034\,
            I => \N__28998\
        );

    \I__6723\ : LocalMux
    port map (
            O => \N__29031\,
            I => \eeprom.eeprom_counter_31\
        );

    \I__6722\ : Odrv12
    port map (
            O => \N__29028\,
            I => \eeprom.eeprom_counter_31\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__29025\,
            I => \eeprom.eeprom_counter_31\
        );

    \I__6720\ : Odrv4
    port map (
            O => \N__29010\,
            I => \eeprom.eeprom_counter_31\
        );

    \I__6719\ : Odrv4
    port map (
            O => \N__29001\,
            I => \eeprom.eeprom_counter_31\
        );

    \I__6718\ : Odrv4
    port map (
            O => \N__28998\,
            I => \eeprom.eeprom_counter_31\
        );

    \I__6717\ : CascadeMux
    port map (
            O => \N__28985\,
            I => \N__28982\
        );

    \I__6716\ : InMux
    port map (
            O => \N__28982\,
            I => \N__28977\
        );

    \I__6715\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28974\
        );

    \I__6714\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28971\
        );

    \I__6713\ : LocalMux
    port map (
            O => \N__28977\,
            I => \N__28968\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__28974\,
            I => \N__28962\
        );

    \I__6711\ : LocalMux
    port map (
            O => \N__28971\,
            I => \N__28962\
        );

    \I__6710\ : Span4Mux_v
    port map (
            O => \N__28968\,
            I => \N__28959\
        );

    \I__6709\ : InMux
    port map (
            O => \N__28967\,
            I => \N__28956\
        );

    \I__6708\ : Span4Mux_v
    port map (
            O => \N__28962\,
            I => \N__28953\
        );

    \I__6707\ : Odrv4
    port map (
            O => \N__28959\,
            I => \eeprom.n2_adj_307\
        );

    \I__6706\ : LocalMux
    port map (
            O => \N__28956\,
            I => \eeprom.n2_adj_307\
        );

    \I__6705\ : Odrv4
    port map (
            O => \N__28953\,
            I => \eeprom.n2_adj_307\
        );

    \I__6704\ : InMux
    port map (
            O => \N__28946\,
            I => \N__28943\
        );

    \I__6703\ : LocalMux
    port map (
            O => \N__28943\,
            I => \N__28940\
        );

    \I__6702\ : Odrv12
    port map (
            O => \N__28940\,
            I => \eeprom.n1135\
        );

    \I__6701\ : CascadeMux
    port map (
            O => \N__28937\,
            I => \N__28916\
        );

    \I__6700\ : CascadeMux
    port map (
            O => \N__28936\,
            I => \N__28912\
        );

    \I__6699\ : CascadeMux
    port map (
            O => \N__28935\,
            I => \N__28909\
        );

    \I__6698\ : CascadeMux
    port map (
            O => \N__28934\,
            I => \N__28905\
        );

    \I__6697\ : CascadeMux
    port map (
            O => \N__28933\,
            I => \N__28901\
        );

    \I__6696\ : CascadeMux
    port map (
            O => \N__28932\,
            I => \N__28898\
        );

    \I__6695\ : CascadeMux
    port map (
            O => \N__28931\,
            I => \N__28893\
        );

    \I__6694\ : CascadeMux
    port map (
            O => \N__28930\,
            I => \N__28889\
        );

    \I__6693\ : CascadeMux
    port map (
            O => \N__28929\,
            I => \N__28886\
        );

    \I__6692\ : CascadeMux
    port map (
            O => \N__28928\,
            I => \N__28879\
        );

    \I__6691\ : CascadeMux
    port map (
            O => \N__28927\,
            I => \N__28870\
        );

    \I__6690\ : CascadeMux
    port map (
            O => \N__28926\,
            I => \N__28867\
        );

    \I__6689\ : CascadeMux
    port map (
            O => \N__28925\,
            I => \N__28864\
        );

    \I__6688\ : CascadeMux
    port map (
            O => \N__28924\,
            I => \N__28861\
        );

    \I__6687\ : CascadeMux
    port map (
            O => \N__28923\,
            I => \N__28858\
        );

    \I__6686\ : CascadeMux
    port map (
            O => \N__28922\,
            I => \N__28855\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__28921\,
            I => \N__28852\
        );

    \I__6684\ : CascadeMux
    port map (
            O => \N__28920\,
            I => \N__28849\
        );

    \I__6683\ : CascadeMux
    port map (
            O => \N__28919\,
            I => \N__28846\
        );

    \I__6682\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28838\
        );

    \I__6681\ : InMux
    port map (
            O => \N__28915\,
            I => \N__28833\
        );

    \I__6680\ : InMux
    port map (
            O => \N__28912\,
            I => \N__28833\
        );

    \I__6679\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28824\
        );

    \I__6678\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28824\
        );

    \I__6677\ : InMux
    port map (
            O => \N__28905\,
            I => \N__28824\
        );

    \I__6676\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28824\
        );

    \I__6675\ : InMux
    port map (
            O => \N__28901\,
            I => \N__28815\
        );

    \I__6674\ : InMux
    port map (
            O => \N__28898\,
            I => \N__28815\
        );

    \I__6673\ : InMux
    port map (
            O => \N__28897\,
            I => \N__28815\
        );

    \I__6672\ : InMux
    port map (
            O => \N__28896\,
            I => \N__28815\
        );

    \I__6671\ : InMux
    port map (
            O => \N__28893\,
            I => \N__28808\
        );

    \I__6670\ : InMux
    port map (
            O => \N__28892\,
            I => \N__28808\
        );

    \I__6669\ : InMux
    port map (
            O => \N__28889\,
            I => \N__28808\
        );

    \I__6668\ : InMux
    port map (
            O => \N__28886\,
            I => \N__28803\
        );

    \I__6667\ : InMux
    port map (
            O => \N__28885\,
            I => \N__28803\
        );

    \I__6666\ : InMux
    port map (
            O => \N__28884\,
            I => \N__28792\
        );

    \I__6665\ : InMux
    port map (
            O => \N__28883\,
            I => \N__28792\
        );

    \I__6664\ : InMux
    port map (
            O => \N__28882\,
            I => \N__28792\
        );

    \I__6663\ : InMux
    port map (
            O => \N__28879\,
            I => \N__28792\
        );

    \I__6662\ : InMux
    port map (
            O => \N__28878\,
            I => \N__28792\
        );

    \I__6661\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28785\
        );

    \I__6660\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28785\
        );

    \I__6659\ : InMux
    port map (
            O => \N__28875\,
            I => \N__28785\
        );

    \I__6658\ : CascadeMux
    port map (
            O => \N__28874\,
            I => \N__28778\
        );

    \I__6657\ : CascadeMux
    port map (
            O => \N__28873\,
            I => \N__28774\
        );

    \I__6656\ : InMux
    port map (
            O => \N__28870\,
            I => \N__28756\
        );

    \I__6655\ : InMux
    port map (
            O => \N__28867\,
            I => \N__28747\
        );

    \I__6654\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28747\
        );

    \I__6653\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28747\
        );

    \I__6652\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28747\
        );

    \I__6651\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28738\
        );

    \I__6650\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28738\
        );

    \I__6649\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28738\
        );

    \I__6648\ : InMux
    port map (
            O => \N__28846\,
            I => \N__28738\
        );

    \I__6647\ : CascadeMux
    port map (
            O => \N__28845\,
            I => \N__28734\
        );

    \I__6646\ : CascadeMux
    port map (
            O => \N__28844\,
            I => \N__28730\
        );

    \I__6645\ : CascadeMux
    port map (
            O => \N__28843\,
            I => \N__28726\
        );

    \I__6644\ : CascadeMux
    port map (
            O => \N__28842\,
            I => \N__28722\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__28841\,
            I => \N__28718\
        );

    \I__6642\ : LocalMux
    port map (
            O => \N__28838\,
            I => \N__28699\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__28833\,
            I => \N__28699\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__28824\,
            I => \N__28699\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__28815\,
            I => \N__28699\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__28808\,
            I => \N__28690\
        );

    \I__6637\ : LocalMux
    port map (
            O => \N__28803\,
            I => \N__28690\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__28792\,
            I => \N__28690\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__28785\,
            I => \N__28690\
        );

    \I__6634\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28685\
        );

    \I__6633\ : InMux
    port map (
            O => \N__28783\,
            I => \N__28685\
        );

    \I__6632\ : InMux
    port map (
            O => \N__28782\,
            I => \N__28676\
        );

    \I__6631\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28676\
        );

    \I__6630\ : InMux
    port map (
            O => \N__28778\,
            I => \N__28676\
        );

    \I__6629\ : InMux
    port map (
            O => \N__28777\,
            I => \N__28676\
        );

    \I__6628\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28669\
        );

    \I__6627\ : InMux
    port map (
            O => \N__28773\,
            I => \N__28669\
        );

    \I__6626\ : InMux
    port map (
            O => \N__28772\,
            I => \N__28669\
        );

    \I__6625\ : InMux
    port map (
            O => \N__28771\,
            I => \N__28660\
        );

    \I__6624\ : InMux
    port map (
            O => \N__28770\,
            I => \N__28660\
        );

    \I__6623\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28660\
        );

    \I__6622\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28660\
        );

    \I__6621\ : InMux
    port map (
            O => \N__28767\,
            I => \N__28651\
        );

    \I__6620\ : InMux
    port map (
            O => \N__28766\,
            I => \N__28651\
        );

    \I__6619\ : InMux
    port map (
            O => \N__28765\,
            I => \N__28651\
        );

    \I__6618\ : InMux
    port map (
            O => \N__28764\,
            I => \N__28651\
        );

    \I__6617\ : CascadeMux
    port map (
            O => \N__28763\,
            I => \N__28648\
        );

    \I__6616\ : CascadeMux
    port map (
            O => \N__28762\,
            I => \N__28645\
        );

    \I__6615\ : CascadeMux
    port map (
            O => \N__28761\,
            I => \N__28641\
        );

    \I__6614\ : CascadeMux
    port map (
            O => \N__28760\,
            I => \N__28638\
        );

    \I__6613\ : CascadeMux
    port map (
            O => \N__28759\,
            I => \N__28635\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__28756\,
            I => \N__28625\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__28747\,
            I => \N__28625\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__28738\,
            I => \N__28625\
        );

    \I__6609\ : InMux
    port map (
            O => \N__28737\,
            I => \N__28616\
        );

    \I__6608\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28616\
        );

    \I__6607\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28616\
        );

    \I__6606\ : InMux
    port map (
            O => \N__28730\,
            I => \N__28616\
        );

    \I__6605\ : InMux
    port map (
            O => \N__28729\,
            I => \N__28607\
        );

    \I__6604\ : InMux
    port map (
            O => \N__28726\,
            I => \N__28607\
        );

    \I__6603\ : InMux
    port map (
            O => \N__28725\,
            I => \N__28607\
        );

    \I__6602\ : InMux
    port map (
            O => \N__28722\,
            I => \N__28607\
        );

    \I__6601\ : InMux
    port map (
            O => \N__28721\,
            I => \N__28604\
        );

    \I__6600\ : InMux
    port map (
            O => \N__28718\,
            I => \N__28601\
        );

    \I__6599\ : CascadeMux
    port map (
            O => \N__28717\,
            I => \N__28596\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__28716\,
            I => \N__28590\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__28715\,
            I => \N__28587\
        );

    \I__6596\ : CascadeMux
    port map (
            O => \N__28714\,
            I => \N__28583\
        );

    \I__6595\ : CascadeMux
    port map (
            O => \N__28713\,
            I => \N__28580\
        );

    \I__6594\ : CascadeMux
    port map (
            O => \N__28712\,
            I => \N__28577\
        );

    \I__6593\ : CascadeMux
    port map (
            O => \N__28711\,
            I => \N__28573\
        );

    \I__6592\ : CascadeMux
    port map (
            O => \N__28710\,
            I => \N__28570\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__28709\,
            I => \N__28567\
        );

    \I__6590\ : CascadeMux
    port map (
            O => \N__28708\,
            I => \N__28564\
        );

    \I__6589\ : Span4Mux_s3_v
    port map (
            O => \N__28699\,
            I => \N__28540\
        );

    \I__6588\ : Span4Mux_v
    port map (
            O => \N__28690\,
            I => \N__28524\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__28685\,
            I => \N__28524\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__28676\,
            I => \N__28524\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__28669\,
            I => \N__28524\
        );

    \I__6584\ : LocalMux
    port map (
            O => \N__28660\,
            I => \N__28524\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__28651\,
            I => \N__28524\
        );

    \I__6582\ : InMux
    port map (
            O => \N__28648\,
            I => \N__28517\
        );

    \I__6581\ : InMux
    port map (
            O => \N__28645\,
            I => \N__28517\
        );

    \I__6580\ : InMux
    port map (
            O => \N__28644\,
            I => \N__28517\
        );

    \I__6579\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28506\
        );

    \I__6578\ : InMux
    port map (
            O => \N__28638\,
            I => \N__28506\
        );

    \I__6577\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28506\
        );

    \I__6576\ : InMux
    port map (
            O => \N__28634\,
            I => \N__28506\
        );

    \I__6575\ : InMux
    port map (
            O => \N__28633\,
            I => \N__28506\
        );

    \I__6574\ : CascadeMux
    port map (
            O => \N__28632\,
            I => \N__28501\
        );

    \I__6573\ : Span4Mux_v
    port map (
            O => \N__28625\,
            I => \N__28489\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__28616\,
            I => \N__28489\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__28607\,
            I => \N__28489\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__28604\,
            I => \N__28489\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28489\
        );

    \I__6568\ : InMux
    port map (
            O => \N__28600\,
            I => \N__28480\
        );

    \I__6567\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28480\
        );

    \I__6566\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28480\
        );

    \I__6565\ : InMux
    port map (
            O => \N__28595\,
            I => \N__28480\
        );

    \I__6564\ : CascadeMux
    port map (
            O => \N__28594\,
            I => \N__28474\
        );

    \I__6563\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28469\
        );

    \I__6562\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28469\
        );

    \I__6561\ : InMux
    port map (
            O => \N__28587\,
            I => \N__28460\
        );

    \I__6560\ : InMux
    port map (
            O => \N__28586\,
            I => \N__28460\
        );

    \I__6559\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28460\
        );

    \I__6558\ : InMux
    port map (
            O => \N__28580\,
            I => \N__28460\
        );

    \I__6557\ : InMux
    port map (
            O => \N__28577\,
            I => \N__28451\
        );

    \I__6556\ : InMux
    port map (
            O => \N__28576\,
            I => \N__28451\
        );

    \I__6555\ : InMux
    port map (
            O => \N__28573\,
            I => \N__28451\
        );

    \I__6554\ : InMux
    port map (
            O => \N__28570\,
            I => \N__28451\
        );

    \I__6553\ : InMux
    port map (
            O => \N__28567\,
            I => \N__28446\
        );

    \I__6552\ : InMux
    port map (
            O => \N__28564\,
            I => \N__28446\
        );

    \I__6551\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28441\
        );

    \I__6550\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28441\
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__28561\,
            I => \N__28437\
        );

    \I__6548\ : CascadeMux
    port map (
            O => \N__28560\,
            I => \N__28434\
        );

    \I__6547\ : CascadeMux
    port map (
            O => \N__28559\,
            I => \N__28430\
        );

    \I__6546\ : CascadeMux
    port map (
            O => \N__28558\,
            I => \N__28425\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__28557\,
            I => \N__28422\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__28556\,
            I => \N__28419\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__28555\,
            I => \N__28415\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__28554\,
            I => \N__28412\
        );

    \I__6541\ : CascadeMux
    port map (
            O => \N__28553\,
            I => \N__28408\
        );

    \I__6540\ : CascadeMux
    port map (
            O => \N__28552\,
            I => \N__28404\
        );

    \I__6539\ : CascadeMux
    port map (
            O => \N__28551\,
            I => \N__28401\
        );

    \I__6538\ : CascadeMux
    port map (
            O => \N__28550\,
            I => \N__28397\
        );

    \I__6537\ : CascadeMux
    port map (
            O => \N__28549\,
            I => \N__28394\
        );

    \I__6536\ : CascadeMux
    port map (
            O => \N__28548\,
            I => \N__28387\
        );

    \I__6535\ : CascadeMux
    port map (
            O => \N__28547\,
            I => \N__28383\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__28546\,
            I => \N__28380\
        );

    \I__6533\ : CascadeMux
    port map (
            O => \N__28545\,
            I => \N__28376\
        );

    \I__6532\ : CascadeMux
    port map (
            O => \N__28544\,
            I => \N__28372\
        );

    \I__6531\ : CascadeMux
    port map (
            O => \N__28543\,
            I => \N__28367\
        );

    \I__6530\ : Span4Mux_v
    port map (
            O => \N__28540\,
            I => \N__28362\
        );

    \I__6529\ : InMux
    port map (
            O => \N__28539\,
            I => \N__28357\
        );

    \I__6528\ : InMux
    port map (
            O => \N__28538\,
            I => \N__28357\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__28537\,
            I => \N__28353\
        );

    \I__6526\ : Span4Mux_v
    port map (
            O => \N__28524\,
            I => \N__28345\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__28517\,
            I => \N__28345\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__28506\,
            I => \N__28345\
        );

    \I__6523\ : InMux
    port map (
            O => \N__28505\,
            I => \N__28340\
        );

    \I__6522\ : InMux
    port map (
            O => \N__28504\,
            I => \N__28340\
        );

    \I__6521\ : InMux
    port map (
            O => \N__28501\,
            I => \N__28335\
        );

    \I__6520\ : InMux
    port map (
            O => \N__28500\,
            I => \N__28335\
        );

    \I__6519\ : Span4Mux_v
    port map (
            O => \N__28489\,
            I => \N__28330\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__28480\,
            I => \N__28330\
        );

    \I__6517\ : InMux
    port map (
            O => \N__28479\,
            I => \N__28325\
        );

    \I__6516\ : InMux
    port map (
            O => \N__28478\,
            I => \N__28325\
        );

    \I__6515\ : InMux
    port map (
            O => \N__28477\,
            I => \N__28320\
        );

    \I__6514\ : InMux
    port map (
            O => \N__28474\,
            I => \N__28320\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__28469\,
            I => \N__28311\
        );

    \I__6512\ : LocalMux
    port map (
            O => \N__28460\,
            I => \N__28311\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__28451\,
            I => \N__28311\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28306\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__28441\,
            I => \N__28306\
        );

    \I__6508\ : InMux
    port map (
            O => \N__28440\,
            I => \N__28303\
        );

    \I__6507\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28298\
        );

    \I__6506\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28298\
        );

    \I__6505\ : InMux
    port map (
            O => \N__28433\,
            I => \N__28295\
        );

    \I__6504\ : InMux
    port map (
            O => \N__28430\,
            I => \N__28292\
        );

    \I__6503\ : InMux
    port map (
            O => \N__28429\,
            I => \N__28278\
        );

    \I__6502\ : InMux
    port map (
            O => \N__28428\,
            I => \N__28278\
        );

    \I__6501\ : InMux
    port map (
            O => \N__28425\,
            I => \N__28278\
        );

    \I__6500\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28278\
        );

    \I__6499\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28269\
        );

    \I__6498\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28269\
        );

    \I__6497\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28269\
        );

    \I__6496\ : InMux
    port map (
            O => \N__28412\,
            I => \N__28269\
        );

    \I__6495\ : CascadeMux
    port map (
            O => \N__28411\,
            I => \N__28265\
        );

    \I__6494\ : InMux
    port map (
            O => \N__28408\,
            I => \N__28261\
        );

    \I__6493\ : InMux
    port map (
            O => \N__28407\,
            I => \N__28252\
        );

    \I__6492\ : InMux
    port map (
            O => \N__28404\,
            I => \N__28252\
        );

    \I__6491\ : InMux
    port map (
            O => \N__28401\,
            I => \N__28252\
        );

    \I__6490\ : InMux
    port map (
            O => \N__28400\,
            I => \N__28252\
        );

    \I__6489\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28247\
        );

    \I__6488\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28247\
        );

    \I__6487\ : CascadeMux
    port map (
            O => \N__28393\,
            I => \N__28244\
        );

    \I__6486\ : InMux
    port map (
            O => \N__28392\,
            I => \N__28237\
        );

    \I__6485\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28237\
        );

    \I__6484\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28230\
        );

    \I__6483\ : InMux
    port map (
            O => \N__28387\,
            I => \N__28230\
        );

    \I__6482\ : InMux
    port map (
            O => \N__28386\,
            I => \N__28230\
        );

    \I__6481\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28219\
        );

    \I__6480\ : InMux
    port map (
            O => \N__28380\,
            I => \N__28219\
        );

    \I__6479\ : InMux
    port map (
            O => \N__28379\,
            I => \N__28219\
        );

    \I__6478\ : InMux
    port map (
            O => \N__28376\,
            I => \N__28219\
        );

    \I__6477\ : InMux
    port map (
            O => \N__28375\,
            I => \N__28219\
        );

    \I__6476\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28216\
        );

    \I__6475\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28213\
        );

    \I__6474\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28204\
        );

    \I__6473\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28204\
        );

    \I__6472\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28204\
        );

    \I__6471\ : InMux
    port map (
            O => \N__28365\,
            I => \N__28204\
        );

    \I__6470\ : Span4Mux_v
    port map (
            O => \N__28362\,
            I => \N__28199\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__28357\,
            I => \N__28199\
        );

    \I__6468\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28194\
        );

    \I__6467\ : InMux
    port map (
            O => \N__28353\,
            I => \N__28194\
        );

    \I__6466\ : CascadeMux
    port map (
            O => \N__28352\,
            I => \N__28191\
        );

    \I__6465\ : Span4Mux_h
    port map (
            O => \N__28345\,
            I => \N__28185\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28185\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__28335\,
            I => \N__28178\
        );

    \I__6462\ : Span4Mux_h
    port map (
            O => \N__28330\,
            I => \N__28178\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__28325\,
            I => \N__28178\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__28320\,
            I => \N__28175\
        );

    \I__6459\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28170\
        );

    \I__6458\ : InMux
    port map (
            O => \N__28318\,
            I => \N__28170\
        );

    \I__6457\ : Span4Mux_s3_v
    port map (
            O => \N__28311\,
            I => \N__28164\
        );

    \I__6456\ : Span4Mux_s3_v
    port map (
            O => \N__28306\,
            I => \N__28164\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__28303\,
            I => \N__28161\
        );

    \I__6454\ : LocalMux
    port map (
            O => \N__28298\,
            I => \N__28154\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__28295\,
            I => \N__28154\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__28292\,
            I => \N__28154\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__28291\,
            I => \N__28150\
        );

    \I__6450\ : CascadeMux
    port map (
            O => \N__28290\,
            I => \N__28146\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__28289\,
            I => \N__28142\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__28288\,
            I => \N__28138\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__28287\,
            I => \N__28135\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__28278\,
            I => \N__28129\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__28269\,
            I => \N__28129\
        );

    \I__6444\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28122\
        );

    \I__6443\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28122\
        );

    \I__6442\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28122\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__28261\,
            I => \N__28115\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__28252\,
            I => \N__28115\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__28247\,
            I => \N__28115\
        );

    \I__6438\ : InMux
    port map (
            O => \N__28244\,
            I => \N__28112\
        );

    \I__6437\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28109\
        );

    \I__6436\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28106\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__28237\,
            I => \N__28090\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__28230\,
            I => \N__28090\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__28219\,
            I => \N__28090\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__28216\,
            I => \N__28090\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__28213\,
            I => \N__28090\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__28204\,
            I => \N__28090\
        );

    \I__6429\ : Span4Mux_v
    port map (
            O => \N__28199\,
            I => \N__28085\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__28194\,
            I => \N__28085\
        );

    \I__6427\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28082\
        );

    \I__6426\ : InMux
    port map (
            O => \N__28190\,
            I => \N__28079\
        );

    \I__6425\ : Span4Mux_v
    port map (
            O => \N__28185\,
            I => \N__28076\
        );

    \I__6424\ : Span4Mux_v
    port map (
            O => \N__28178\,
            I => \N__28069\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__28175\,
            I => \N__28069\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28069\
        );

    \I__6421\ : InMux
    port map (
            O => \N__28169\,
            I => \N__28066\
        );

    \I__6420\ : Sp12to4
    port map (
            O => \N__28164\,
            I => \N__28063\
        );

    \I__6419\ : Span4Mux_s3_v
    port map (
            O => \N__28161\,
            I => \N__28058\
        );

    \I__6418\ : Span4Mux_h
    port map (
            O => \N__28154\,
            I => \N__28058\
        );

    \I__6417\ : InMux
    port map (
            O => \N__28153\,
            I => \N__28055\
        );

    \I__6416\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28048\
        );

    \I__6415\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28048\
        );

    \I__6414\ : InMux
    port map (
            O => \N__28146\,
            I => \N__28048\
        );

    \I__6413\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28039\
        );

    \I__6412\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28039\
        );

    \I__6411\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28039\
        );

    \I__6410\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28039\
        );

    \I__6409\ : InMux
    port map (
            O => \N__28135\,
            I => \N__28036\
        );

    \I__6408\ : InMux
    port map (
            O => \N__28134\,
            I => \N__28033\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__28129\,
            I => \N__28026\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__28122\,
            I => \N__28026\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__28115\,
            I => \N__28021\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__28112\,
            I => \N__28021\
        );

    \I__6403\ : LocalMux
    port map (
            O => \N__28109\,
            I => \N__28016\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__28106\,
            I => \N__28016\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__28105\,
            I => \N__28012\
        );

    \I__6400\ : CascadeMux
    port map (
            O => \N__28104\,
            I => \N__28008\
        );

    \I__6399\ : CascadeMux
    port map (
            O => \N__28103\,
            I => \N__28004\
        );

    \I__6398\ : Span12Mux_v
    port map (
            O => \N__28090\,
            I => \N__28000\
        );

    \I__6397\ : Span4Mux_h
    port map (
            O => \N__28085\,
            I => \N__27993\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__28082\,
            I => \N__27993\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__28079\,
            I => \N__27993\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__28076\,
            I => \N__27988\
        );

    \I__6393\ : Span4Mux_v
    port map (
            O => \N__28069\,
            I => \N__27988\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__27985\
        );

    \I__6391\ : Span12Mux_s11_h
    port map (
            O => \N__28063\,
            I => \N__27970\
        );

    \I__6390\ : Sp12to4
    port map (
            O => \N__28058\,
            I => \N__27970\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__28055\,
            I => \N__27970\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__28048\,
            I => \N__27970\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__28039\,
            I => \N__27970\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__28036\,
            I => \N__27970\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__28033\,
            I => \N__27970\
        );

    \I__6384\ : InMux
    port map (
            O => \N__28032\,
            I => \N__27965\
        );

    \I__6383\ : InMux
    port map (
            O => \N__28031\,
            I => \N__27965\
        );

    \I__6382\ : Span4Mux_v
    port map (
            O => \N__28026\,
            I => \N__27960\
        );

    \I__6381\ : Span4Mux_v
    port map (
            O => \N__28021\,
            I => \N__27960\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__28016\,
            I => \N__27957\
        );

    \I__6379\ : InMux
    port map (
            O => \N__28015\,
            I => \N__27942\
        );

    \I__6378\ : InMux
    port map (
            O => \N__28012\,
            I => \N__27942\
        );

    \I__6377\ : InMux
    port map (
            O => \N__28011\,
            I => \N__27942\
        );

    \I__6376\ : InMux
    port map (
            O => \N__28008\,
            I => \N__27942\
        );

    \I__6375\ : InMux
    port map (
            O => \N__28007\,
            I => \N__27942\
        );

    \I__6374\ : InMux
    port map (
            O => \N__28004\,
            I => \N__27942\
        );

    \I__6373\ : InMux
    port map (
            O => \N__28003\,
            I => \N__27942\
        );

    \I__6372\ : Span12Mux_h
    port map (
            O => \N__28000\,
            I => \N__27939\
        );

    \I__6371\ : Span4Mux_h
    port map (
            O => \N__27993\,
            I => \N__27936\
        );

    \I__6370\ : Span4Mux_h
    port map (
            O => \N__27988\,
            I => \N__27931\
        );

    \I__6369\ : Span4Mux_v
    port map (
            O => \N__27985\,
            I => \N__27931\
        );

    \I__6368\ : Span12Mux_v
    port map (
            O => \N__27970\,
            I => \N__27926\
        );

    \I__6367\ : LocalMux
    port map (
            O => \N__27965\,
            I => \N__27926\
        );

    \I__6366\ : Span4Mux_h
    port map (
            O => \N__27960\,
            I => \N__27919\
        );

    \I__6365\ : Span4Mux_h
    port map (
            O => \N__27957\,
            I => \N__27919\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__27942\,
            I => \N__27919\
        );

    \I__6363\ : Odrv12
    port map (
            O => \N__27939\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6362\ : Odrv4
    port map (
            O => \N__27936\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6361\ : Odrv4
    port map (
            O => \N__27931\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6360\ : Odrv12
    port map (
            O => \N__27926\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6359\ : Odrv4
    port map (
            O => \N__27919\,
            I => \CONSTANT_ONE_NET\
        );

    \I__6358\ : InMux
    port map (
            O => \N__27908\,
            I => \N__27905\
        );

    \I__6357\ : LocalMux
    port map (
            O => \N__27905\,
            I => n174
        );

    \I__6356\ : CascadeMux
    port map (
            O => \N__27902\,
            I => \N__27899\
        );

    \I__6355\ : InMux
    port map (
            O => \N__27899\,
            I => \N__27896\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__27896\,
            I => \N__27892\
        );

    \I__6353\ : InMux
    port map (
            O => \N__27895\,
            I => \N__27889\
        );

    \I__6352\ : Odrv12
    port map (
            O => \N__27892\,
            I => rw
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__27889\,
            I => rw
        );

    \I__6350\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27881\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__27881\,
            I => \N__27876\
        );

    \I__6348\ : InMux
    port map (
            O => \N__27880\,
            I => \N__27873\
        );

    \I__6347\ : InMux
    port map (
            O => \N__27879\,
            I => \N__27870\
        );

    \I__6346\ : Span4Mux_v
    port map (
            O => \N__27876\,
            I => \N__27867\
        );

    \I__6345\ : LocalMux
    port map (
            O => \N__27873\,
            I => \N__27864\
        );

    \I__6344\ : LocalMux
    port map (
            O => \N__27870\,
            I => saved_addr_0
        );

    \I__6343\ : Odrv4
    port map (
            O => \N__27867\,
            I => saved_addr_0
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__27864\,
            I => saved_addr_0
        );

    \I__6341\ : InMux
    port map (
            O => \N__27857\,
            I => \eeprom.n4278\
        );

    \I__6340\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27851\
        );

    \I__6339\ : LocalMux
    port map (
            O => \N__27851\,
            I => \N__27848\
        );

    \I__6338\ : Odrv4
    port map (
            O => \N__27848\,
            I => \eeprom.n1192\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__27845\,
            I => \N__27840\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__27844\,
            I => \N__27837\
        );

    \I__6335\ : InMux
    port map (
            O => \N__27843\,
            I => \N__27834\
        );

    \I__6334\ : InMux
    port map (
            O => \N__27840\,
            I => \N__27831\
        );

    \I__6333\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27828\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__27834\,
            I => \N__27823\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__27831\,
            I => \N__27823\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__27828\,
            I => \eeprom.n1256\
        );

    \I__6329\ : Odrv4
    port map (
            O => \N__27823\,
            I => \eeprom.n1256\
        );

    \I__6328\ : CascadeMux
    port map (
            O => \N__27818\,
            I => \eeprom.n1843_cascade_\
        );

    \I__6327\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27812\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__27812\,
            I => \eeprom.n1195\
        );

    \I__6325\ : CascadeMux
    port map (
            O => \N__27809\,
            I => \N__27805\
        );

    \I__6324\ : InMux
    port map (
            O => \N__27808\,
            I => \N__27802\
        );

    \I__6323\ : InMux
    port map (
            O => \N__27805\,
            I => \N__27799\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__27802\,
            I => \N__27794\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__27799\,
            I => \N__27794\
        );

    \I__6320\ : Span4Mux_v
    port map (
            O => \N__27794\,
            I => \N__27790\
        );

    \I__6319\ : InMux
    port map (
            O => \N__27793\,
            I => \N__27787\
        );

    \I__6318\ : Odrv4
    port map (
            O => \N__27790\,
            I => \eeprom.n1915\
        );

    \I__6317\ : LocalMux
    port map (
            O => \N__27787\,
            I => \eeprom.n1915\
        );

    \I__6316\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27779\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27775\
        );

    \I__6314\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27771\
        );

    \I__6313\ : Span4Mux_h
    port map (
            O => \N__27775\,
            I => \N__27768\
        );

    \I__6312\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27765\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__27771\,
            I => \eeprom.eeprom_counter_29\
        );

    \I__6310\ : Odrv4
    port map (
            O => \N__27768\,
            I => \eeprom.eeprom_counter_29\
        );

    \I__6309\ : LocalMux
    port map (
            O => \N__27765\,
            I => \eeprom.eeprom_counter_29\
        );

    \I__6308\ : InMux
    port map (
            O => \N__27758\,
            I => \N__27755\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__27755\,
            I => \N__27752\
        );

    \I__6306\ : Span4Mux_h
    port map (
            O => \N__27752\,
            I => \N__27749\
        );

    \I__6305\ : Odrv4
    port map (
            O => \N__27749\,
            I => \eeprom.n4_adj_310\
        );

    \I__6304\ : CascadeMux
    port map (
            O => \N__27746\,
            I => \N__27743\
        );

    \I__6303\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27738\
        );

    \I__6302\ : InMux
    port map (
            O => \N__27742\,
            I => \N__27733\
        );

    \I__6301\ : InMux
    port map (
            O => \N__27741\,
            I => \N__27733\
        );

    \I__6300\ : LocalMux
    port map (
            O => \N__27738\,
            I => \eeprom.n1138\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__27733\,
            I => \eeprom.n1138\
        );

    \I__6298\ : CascadeMux
    port map (
            O => \N__27728\,
            I => \eeprom.n1137_cascade_\
        );

    \I__6297\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27721\
        );

    \I__6296\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27718\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__27721\,
            I => \eeprom.n4977\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__27718\,
            I => \eeprom.n4977\
        );

    \I__6293\ : InMux
    port map (
            O => \N__27713\,
            I => \N__27710\
        );

    \I__6292\ : LocalMux
    port map (
            O => \N__27710\,
            I => \eeprom.n4983\
        );

    \I__6291\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27704\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__27704\,
            I => \eeprom.n1197\
        );

    \I__6289\ : CascadeMux
    port map (
            O => \N__27701\,
            I => \N__27697\
        );

    \I__6288\ : CascadeMux
    port map (
            O => \N__27700\,
            I => \N__27694\
        );

    \I__6287\ : InMux
    port map (
            O => \N__27697\,
            I => \N__27691\
        );

    \I__6286\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27688\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__27691\,
            I => \N__27685\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__27688\,
            I => \N__27682\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__27685\,
            I => \N__27678\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__27682\,
            I => \N__27675\
        );

    \I__6281\ : InMux
    port map (
            O => \N__27681\,
            I => \N__27672\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__27678\,
            I => \eeprom.n1917\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__27675\,
            I => \eeprom.n1917\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__27672\,
            I => \eeprom.n1917\
        );

    \I__6277\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27662\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__27662\,
            I => \eeprom.n1194\
        );

    \I__6275\ : CascadeMux
    port map (
            O => \N__27659\,
            I => \N__27656\
        );

    \I__6274\ : InMux
    port map (
            O => \N__27656\,
            I => \N__27651\
        );

    \I__6273\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27648\
        );

    \I__6272\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27645\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__27651\,
            I => \eeprom.n1137\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__27648\,
            I => \eeprom.n1137\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__27645\,
            I => \eeprom.n1137\
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__27638\,
            I => \N__27632\
        );

    \I__6267\ : InMux
    port map (
            O => \N__27637\,
            I => \N__27624\
        );

    \I__6266\ : InMux
    port map (
            O => \N__27636\,
            I => \N__27624\
        );

    \I__6265\ : InMux
    port map (
            O => \N__27635\,
            I => \N__27624\
        );

    \I__6264\ : InMux
    port map (
            O => \N__27632\,
            I => \N__27619\
        );

    \I__6263\ : InMux
    port map (
            O => \N__27631\,
            I => \N__27619\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__27624\,
            I => \eeprom.n1843\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__27619\,
            I => \eeprom.n1843\
        );

    \I__6260\ : CascadeMux
    port map (
            O => \N__27614\,
            I => \N__27610\
        );

    \I__6259\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27607\
        );

    \I__6258\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27604\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__27607\,
            I => \N__27601\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__27604\,
            I => \N__27598\
        );

    \I__6255\ : Span4Mux_v
    port map (
            O => \N__27601\,
            I => \N__27594\
        );

    \I__6254\ : Span4Mux_h
    port map (
            O => \N__27598\,
            I => \N__27591\
        );

    \I__6253\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27588\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__27594\,
            I => \eeprom.n1914\
        );

    \I__6251\ : Odrv4
    port map (
            O => \N__27591\,
            I => \eeprom.n1914\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__27588\,
            I => \eeprom.n1914\
        );

    \I__6249\ : InMux
    port map (
            O => \N__27581\,
            I => \N__27577\
        );

    \I__6248\ : InMux
    port map (
            O => \N__27580\,
            I => \N__27574\
        );

    \I__6247\ : LocalMux
    port map (
            O => \N__27577\,
            I => \N__27570\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__27574\,
            I => \N__27567\
        );

    \I__6245\ : InMux
    port map (
            O => \N__27573\,
            I => \N__27564\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__27570\,
            I => \N__27561\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__27567\,
            I => \N__27558\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__27564\,
            I => \eeprom.eeprom_counter_14\
        );

    \I__6241\ : Odrv4
    port map (
            O => \N__27561\,
            I => \eeprom.eeprom_counter_14\
        );

    \I__6240\ : Odrv4
    port map (
            O => \N__27558\,
            I => \eeprom.eeprom_counter_14\
        );

    \I__6239\ : CascadeMux
    port map (
            O => \N__27551\,
            I => \N__27548\
        );

    \I__6238\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27545\
        );

    \I__6237\ : LocalMux
    port map (
            O => \N__27545\,
            I => \eeprom.n19\
        );

    \I__6236\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27535\
        );

    \I__6235\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27528\
        );

    \I__6234\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27528\
        );

    \I__6233\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27528\
        );

    \I__6232\ : CascadeMux
    port map (
            O => \N__27538\,
            I => \N__27517\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__27535\,
            I => \N__27508\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27508\
        );

    \I__6229\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27503\
        );

    \I__6228\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27503\
        );

    \I__6227\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27496\
        );

    \I__6226\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27496\
        );

    \I__6225\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27496\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__27522\,
            I => \N__27490\
        );

    \I__6223\ : InMux
    port map (
            O => \N__27521\,
            I => \N__27485\
        );

    \I__6222\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27485\
        );

    \I__6221\ : InMux
    port map (
            O => \N__27517\,
            I => \N__27482\
        );

    \I__6220\ : InMux
    port map (
            O => \N__27516\,
            I => \N__27475\
        );

    \I__6219\ : InMux
    port map (
            O => \N__27515\,
            I => \N__27475\
        );

    \I__6218\ : InMux
    port map (
            O => \N__27514\,
            I => \N__27475\
        );

    \I__6217\ : InMux
    port map (
            O => \N__27513\,
            I => \N__27472\
        );

    \I__6216\ : Span4Mux_v
    port map (
            O => \N__27508\,
            I => \N__27465\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__27503\,
            I => \N__27465\
        );

    \I__6214\ : LocalMux
    port map (
            O => \N__27496\,
            I => \N__27465\
        );

    \I__6213\ : InMux
    port map (
            O => \N__27495\,
            I => \N__27456\
        );

    \I__6212\ : InMux
    port map (
            O => \N__27494\,
            I => \N__27456\
        );

    \I__6211\ : InMux
    port map (
            O => \N__27493\,
            I => \N__27456\
        );

    \I__6210\ : InMux
    port map (
            O => \N__27490\,
            I => \N__27456\
        );

    \I__6209\ : LocalMux
    port map (
            O => \N__27485\,
            I => state_1
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__27482\,
            I => state_1
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__27475\,
            I => state_1
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__27472\,
            I => state_1
        );

    \I__6205\ : Odrv4
    port map (
            O => \N__27465\,
            I => state_1
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__27456\,
            I => state_1
        );

    \I__6203\ : InMux
    port map (
            O => \N__27443\,
            I => \N__27440\
        );

    \I__6202\ : LocalMux
    port map (
            O => \N__27440\,
            I => n3581
        );

    \I__6201\ : InMux
    port map (
            O => \N__27437\,
            I => \N__27433\
        );

    \I__6200\ : InMux
    port map (
            O => \N__27436\,
            I => \N__27430\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__27433\,
            I => \eeprom.i2c.n407\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__27430\,
            I => \eeprom.i2c.n407\
        );

    \I__6197\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27420\
        );

    \I__6196\ : CascadeMux
    port map (
            O => \N__27424\,
            I => \N__27415\
        );

    \I__6195\ : InMux
    port map (
            O => \N__27423\,
            I => \N__27412\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__27420\,
            I => \N__27397\
        );

    \I__6193\ : InMux
    port map (
            O => \N__27419\,
            I => \N__27390\
        );

    \I__6192\ : InMux
    port map (
            O => \N__27418\,
            I => \N__27390\
        );

    \I__6191\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27390\
        );

    \I__6190\ : LocalMux
    port map (
            O => \N__27412\,
            I => \N__27387\
        );

    \I__6189\ : InMux
    port map (
            O => \N__27411\,
            I => \N__27382\
        );

    \I__6188\ : InMux
    port map (
            O => \N__27410\,
            I => \N__27375\
        );

    \I__6187\ : InMux
    port map (
            O => \N__27409\,
            I => \N__27375\
        );

    \I__6186\ : InMux
    port map (
            O => \N__27408\,
            I => \N__27375\
        );

    \I__6185\ : InMux
    port map (
            O => \N__27407\,
            I => \N__27370\
        );

    \I__6184\ : InMux
    port map (
            O => \N__27406\,
            I => \N__27370\
        );

    \I__6183\ : InMux
    port map (
            O => \N__27405\,
            I => \N__27364\
        );

    \I__6182\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27353\
        );

    \I__6181\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27353\
        );

    \I__6180\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27353\
        );

    \I__6179\ : InMux
    port map (
            O => \N__27401\,
            I => \N__27353\
        );

    \I__6178\ : InMux
    port map (
            O => \N__27400\,
            I => \N__27353\
        );

    \I__6177\ : Span4Mux_v
    port map (
            O => \N__27397\,
            I => \N__27348\
        );

    \I__6176\ : LocalMux
    port map (
            O => \N__27390\,
            I => \N__27348\
        );

    \I__6175\ : Span4Mux_h
    port map (
            O => \N__27387\,
            I => \N__27345\
        );

    \I__6174\ : InMux
    port map (
            O => \N__27386\,
            I => \N__27340\
        );

    \I__6173\ : InMux
    port map (
            O => \N__27385\,
            I => \N__27340\
        );

    \I__6172\ : LocalMux
    port map (
            O => \N__27382\,
            I => \N__27333\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__27375\,
            I => \N__27333\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__27370\,
            I => \N__27333\
        );

    \I__6169\ : InMux
    port map (
            O => \N__27369\,
            I => \N__27326\
        );

    \I__6168\ : InMux
    port map (
            O => \N__27368\,
            I => \N__27326\
        );

    \I__6167\ : InMux
    port map (
            O => \N__27367\,
            I => \N__27326\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__27364\,
            I => state_0
        );

    \I__6165\ : LocalMux
    port map (
            O => \N__27353\,
            I => state_0
        );

    \I__6164\ : Odrv4
    port map (
            O => \N__27348\,
            I => state_0
        );

    \I__6163\ : Odrv4
    port map (
            O => \N__27345\,
            I => state_0
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__27340\,
            I => state_0
        );

    \I__6161\ : Odrv4
    port map (
            O => \N__27333\,
            I => state_0
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__27326\,
            I => state_0
        );

    \I__6159\ : IoInMux
    port map (
            O => \N__27311\,
            I => \N__27308\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__27308\,
            I => \N__27305\
        );

    \I__6157\ : Span12Mux_s4_h
    port map (
            O => \N__27305\,
            I => \N__27302\
        );

    \I__6156\ : Span12Mux_v
    port map (
            O => \N__27302\,
            I => \N__27298\
        );

    \I__6155\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27295\
        );

    \I__6154\ : Odrv12
    port map (
            O => \N__27298\,
            I => sda_enable
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__27295\,
            I => sda_enable
        );

    \I__6152\ : CEMux
    port map (
            O => \N__27290\,
            I => \N__27287\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__27287\,
            I => \N__27284\
        );

    \I__6150\ : Span4Mux_h
    port map (
            O => \N__27284\,
            I => \N__27281\
        );

    \I__6149\ : Odrv4
    port map (
            O => \N__27281\,
            I => \eeprom.i2c.n524\
        );

    \I__6148\ : SRMux
    port map (
            O => \N__27278\,
            I => \N__27275\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__27275\,
            I => \N__27272\
        );

    \I__6146\ : Odrv4
    port map (
            O => \N__27272\,
            I => \eeprom.i2c.n1901\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__27269\,
            I => \N__27265\
        );

    \I__6144\ : InMux
    port map (
            O => \N__27268\,
            I => \N__27262\
        );

    \I__6143\ : InMux
    port map (
            O => \N__27265\,
            I => \N__27259\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__27262\,
            I => \eeprom.n892\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__27259\,
            I => \eeprom.n892\
        );

    \I__6140\ : CascadeMux
    port map (
            O => \N__27254\,
            I => \N__27251\
        );

    \I__6139\ : InMux
    port map (
            O => \N__27251\,
            I => \N__27248\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__27248\,
            I => \eeprom.n1198\
        );

    \I__6137\ : InMux
    port map (
            O => \N__27245\,
            I => \bfn_28_21_0_\
        );

    \I__6136\ : InMux
    port map (
            O => \N__27242\,
            I => \eeprom.n4273\
        );

    \I__6135\ : CascadeMux
    port map (
            O => \N__27239\,
            I => \N__27236\
        );

    \I__6134\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27233\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__27233\,
            I => \eeprom.n1139\
        );

    \I__6132\ : InMux
    port map (
            O => \N__27230\,
            I => \N__27227\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__27227\,
            I => \eeprom.n1196\
        );

    \I__6130\ : InMux
    port map (
            O => \N__27224\,
            I => \eeprom.n4274\
        );

    \I__6129\ : InMux
    port map (
            O => \N__27221\,
            I => \eeprom.n4275\
        );

    \I__6128\ : InMux
    port map (
            O => \N__27218\,
            I => \eeprom.n4276\
        );

    \I__6127\ : InMux
    port map (
            O => \N__27215\,
            I => \N__27212\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__27212\,
            I => \eeprom.n5327\
        );

    \I__6125\ : CascadeMux
    port map (
            O => \N__27209\,
            I => \N__27205\
        );

    \I__6124\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27202\
        );

    \I__6123\ : InMux
    port map (
            O => \N__27205\,
            I => \N__27199\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__27202\,
            I => \eeprom.n5328\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__27199\,
            I => \eeprom.n5328\
        );

    \I__6120\ : InMux
    port map (
            O => \N__27194\,
            I => \eeprom.n4277\
        );

    \I__6119\ : InMux
    port map (
            O => \N__27191\,
            I => \N__27188\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__27188\,
            I => n11_adj_359
        );

    \I__6117\ : InMux
    port map (
            O => \N__27185\,
            I => \N__27182\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__27182\,
            I => n5458
        );

    \I__6115\ : CascadeMux
    port map (
            O => \N__27179\,
            I => \n6_adj_365_cascade_\
        );

    \I__6114\ : InMux
    port map (
            O => \N__27176\,
            I => \N__27171\
        );

    \I__6113\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27166\
        );

    \I__6112\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27166\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__27171\,
            I => n471
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__27166\,
            I => n471
        );

    \I__6109\ : CascadeMux
    port map (
            O => \N__27161\,
            I => \N__27154\
        );

    \I__6108\ : CascadeMux
    port map (
            O => \N__27160\,
            I => \N__27145\
        );

    \I__6107\ : CascadeMux
    port map (
            O => \N__27159\,
            I => \N__27139\
        );

    \I__6106\ : InMux
    port map (
            O => \N__27158\,
            I => \N__27133\
        );

    \I__6105\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27133\
        );

    \I__6104\ : InMux
    port map (
            O => \N__27154\,
            I => \N__27126\
        );

    \I__6103\ : InMux
    port map (
            O => \N__27153\,
            I => \N__27119\
        );

    \I__6102\ : InMux
    port map (
            O => \N__27152\,
            I => \N__27119\
        );

    \I__6101\ : InMux
    port map (
            O => \N__27151\,
            I => \N__27119\
        );

    \I__6100\ : InMux
    port map (
            O => \N__27150\,
            I => \N__27112\
        );

    \I__6099\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27112\
        );

    \I__6098\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27112\
        );

    \I__6097\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27107\
        );

    \I__6096\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27107\
        );

    \I__6095\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27104\
        );

    \I__6094\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27101\
        );

    \I__6093\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27096\
        );

    \I__6092\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27096\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__27133\,
            I => \N__27093\
        );

    \I__6090\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27084\
        );

    \I__6089\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27084\
        );

    \I__6088\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27084\
        );

    \I__6087\ : InMux
    port map (
            O => \N__27129\,
            I => \N__27084\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__27126\,
            I => state_3
        );

    \I__6085\ : LocalMux
    port map (
            O => \N__27119\,
            I => state_3
        );

    \I__6084\ : LocalMux
    port map (
            O => \N__27112\,
            I => state_3
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__27107\,
            I => state_3
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__27104\,
            I => state_3
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__27101\,
            I => state_3
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__27096\,
            I => state_3
        );

    \I__6079\ : Odrv4
    port map (
            O => \N__27093\,
            I => state_3
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__27084\,
            I => state_3
        );

    \I__6077\ : InMux
    port map (
            O => \N__27065\,
            I => \N__27062\
        );

    \I__6076\ : LocalMux
    port map (
            O => \N__27062\,
            I => n3587
        );

    \I__6075\ : CascadeMux
    port map (
            O => \N__27059\,
            I => \n3587_cascade_\
        );

    \I__6074\ : InMux
    port map (
            O => \N__27056\,
            I => \N__27052\
        );

    \I__6073\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27049\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__27052\,
            I => n10
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__27049\,
            I => n10
        );

    \I__6070\ : InMux
    port map (
            O => \N__27044\,
            I => \N__27041\
        );

    \I__6069\ : LocalMux
    port map (
            O => \N__27041\,
            I => n5454
        );

    \I__6068\ : CascadeMux
    port map (
            O => \N__27038\,
            I => \N__27033\
        );

    \I__6067\ : InMux
    port map (
            O => \N__27037\,
            I => \N__27029\
        );

    \I__6066\ : InMux
    port map (
            O => \N__27036\,
            I => \N__27024\
        );

    \I__6065\ : InMux
    port map (
            O => \N__27033\,
            I => \N__27021\
        );

    \I__6064\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27018\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__27029\,
            I => \N__27015\
        );

    \I__6062\ : InMux
    port map (
            O => \N__27028\,
            I => \N__27012\
        );

    \I__6061\ : InMux
    port map (
            O => \N__27027\,
            I => \N__27009\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__27024\,
            I => \N__27006\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__27021\,
            I => \eeprom.i2c.counter_1\
        );

    \I__6058\ : LocalMux
    port map (
            O => \N__27018\,
            I => \eeprom.i2c.counter_1\
        );

    \I__6057\ : Odrv4
    port map (
            O => \N__27015\,
            I => \eeprom.i2c.counter_1\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__27012\,
            I => \eeprom.i2c.counter_1\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__27009\,
            I => \eeprom.i2c.counter_1\
        );

    \I__6054\ : Odrv4
    port map (
            O => \N__27006\,
            I => \eeprom.i2c.counter_1\
        );

    \I__6053\ : InMux
    port map (
            O => \N__26993\,
            I => \N__26990\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__26990\,
            I => \N__26983\
        );

    \I__6051\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26979\
        );

    \I__6050\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26976\
        );

    \I__6049\ : InMux
    port map (
            O => \N__26987\,
            I => \N__26971\
        );

    \I__6048\ : InMux
    port map (
            O => \N__26986\,
            I => \N__26971\
        );

    \I__6047\ : Span4Mux_v
    port map (
            O => \N__26983\,
            I => \N__26968\
        );

    \I__6046\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26965\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__26979\,
            I => \N__26962\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__26976\,
            I => \eeprom.i2c.counter_2\
        );

    \I__6043\ : LocalMux
    port map (
            O => \N__26971\,
            I => \eeprom.i2c.counter_2\
        );

    \I__6042\ : Odrv4
    port map (
            O => \N__26968\,
            I => \eeprom.i2c.counter_2\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__26965\,
            I => \eeprom.i2c.counter_2\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__26962\,
            I => \eeprom.i2c.counter_2\
        );

    \I__6039\ : CascadeMux
    port map (
            O => \N__26951\,
            I => \N__26944\
        );

    \I__6038\ : InMux
    port map (
            O => \N__26950\,
            I => \N__26941\
        );

    \I__6037\ : InMux
    port map (
            O => \N__26949\,
            I => \N__26936\
        );

    \I__6036\ : InMux
    port map (
            O => \N__26948\,
            I => \N__26936\
        );

    \I__6035\ : InMux
    port map (
            O => \N__26947\,
            I => \N__26933\
        );

    \I__6034\ : InMux
    port map (
            O => \N__26944\,
            I => \N__26930\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__26941\,
            I => \N__26927\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__26936\,
            I => \eeprom.i2c.counter_0\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__26933\,
            I => \eeprom.i2c.counter_0\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__26930\,
            I => \eeprom.i2c.counter_0\
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__26927\,
            I => \eeprom.i2c.counter_0\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__26918\,
            I => \eeprom.i2c.n5464_cascade_\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__26915\,
            I => \eeprom.i2c.n5451_cascade_\
        );

    \I__6026\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26909\
        );

    \I__6025\ : LocalMux
    port map (
            O => \N__26909\,
            I => \eeprom.i2c.sda_out\
        );

    \I__6024\ : CEMux
    port map (
            O => \N__26906\,
            I => \N__26903\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__26903\,
            I => \N__26900\
        );

    \I__6022\ : Odrv12
    port map (
            O => \N__26900\,
            I => \eeprom.i2c.n4513\
        );

    \I__6021\ : CascadeMux
    port map (
            O => \N__26897\,
            I => \N__26888\
        );

    \I__6020\ : CascadeMux
    port map (
            O => \N__26896\,
            I => \N__26882\
        );

    \I__6019\ : CascadeMux
    port map (
            O => \N__26895\,
            I => \N__26879\
        );

    \I__6018\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26872\
        );

    \I__6017\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26872\
        );

    \I__6016\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26869\
        );

    \I__6015\ : InMux
    port map (
            O => \N__26891\,
            I => \N__26866\
        );

    \I__6014\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26861\
        );

    \I__6013\ : InMux
    port map (
            O => \N__26887\,
            I => \N__26861\
        );

    \I__6012\ : InMux
    port map (
            O => \N__26886\,
            I => \N__26858\
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__26885\,
            I => \N__26855\
        );

    \I__6010\ : InMux
    port map (
            O => \N__26882\,
            I => \N__26850\
        );

    \I__6009\ : InMux
    port map (
            O => \N__26879\,
            I => \N__26847\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__26878\,
            I => \N__26844\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__26877\,
            I => \N__26841\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__26872\,
            I => \N__26836\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__26869\,
            I => \N__26833\
        );

    \I__6004\ : LocalMux
    port map (
            O => \N__26866\,
            I => \N__26828\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__26861\,
            I => \N__26828\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__26858\,
            I => \N__26825\
        );

    \I__6001\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26820\
        );

    \I__6000\ : InMux
    port map (
            O => \N__26854\,
            I => \N__26820\
        );

    \I__5999\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26812\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__26850\,
            I => \N__26807\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__26847\,
            I => \N__26807\
        );

    \I__5996\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26798\
        );

    \I__5995\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26798\
        );

    \I__5994\ : InMux
    port map (
            O => \N__26840\,
            I => \N__26798\
        );

    \I__5993\ : InMux
    port map (
            O => \N__26839\,
            I => \N__26798\
        );

    \I__5992\ : Span4Mux_h
    port map (
            O => \N__26836\,
            I => \N__26795\
        );

    \I__5991\ : Span4Mux_v
    port map (
            O => \N__26833\,
            I => \N__26790\
        );

    \I__5990\ : Span4Mux_h
    port map (
            O => \N__26828\,
            I => \N__26790\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__26825\,
            I => \N__26785\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26785\
        );

    \I__5987\ : InMux
    port map (
            O => \N__26819\,
            I => \N__26782\
        );

    \I__5986\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26775\
        );

    \I__5985\ : InMux
    port map (
            O => \N__26817\,
            I => \N__26775\
        );

    \I__5984\ : InMux
    port map (
            O => \N__26816\,
            I => \N__26775\
        );

    \I__5983\ : InMux
    port map (
            O => \N__26815\,
            I => \N__26772\
        );

    \I__5982\ : LocalMux
    port map (
            O => \N__26812\,
            I => state_2
        );

    \I__5981\ : Odrv4
    port map (
            O => \N__26807\,
            I => state_2
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__26798\,
            I => state_2
        );

    \I__5979\ : Odrv4
    port map (
            O => \N__26795\,
            I => state_2
        );

    \I__5978\ : Odrv4
    port map (
            O => \N__26790\,
            I => state_2
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__26785\,
            I => state_2
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__26782\,
            I => state_2
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__26775\,
            I => state_2
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__26772\,
            I => state_2
        );

    \I__5973\ : InMux
    port map (
            O => \N__26753\,
            I => \N__26747\
        );

    \I__5972\ : InMux
    port map (
            O => \N__26752\,
            I => \N__26747\
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__26747\,
            I => n3595
        );

    \I__5970\ : CascadeMux
    port map (
            O => \N__26744\,
            I => \N__26732\
        );

    \I__5969\ : InMux
    port map (
            O => \N__26743\,
            I => \N__26724\
        );

    \I__5968\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26724\
        );

    \I__5967\ : InMux
    port map (
            O => \N__26741\,
            I => \N__26724\
        );

    \I__5966\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26721\
        );

    \I__5965\ : CascadeMux
    port map (
            O => \N__26739\,
            I => \N__26717\
        );

    \I__5964\ : CascadeMux
    port map (
            O => \N__26738\,
            I => \N__26713\
        );

    \I__5963\ : CascadeMux
    port map (
            O => \N__26737\,
            I => \N__26709\
        );

    \I__5962\ : InMux
    port map (
            O => \N__26736\,
            I => \N__26699\
        );

    \I__5961\ : InMux
    port map (
            O => \N__26735\,
            I => \N__26699\
        );

    \I__5960\ : InMux
    port map (
            O => \N__26732\,
            I => \N__26699\
        );

    \I__5959\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26699\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__26724\,
            I => \N__26694\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__26721\,
            I => \N__26694\
        );

    \I__5956\ : InMux
    port map (
            O => \N__26720\,
            I => \N__26679\
        );

    \I__5955\ : InMux
    port map (
            O => \N__26717\,
            I => \N__26679\
        );

    \I__5954\ : InMux
    port map (
            O => \N__26716\,
            I => \N__26679\
        );

    \I__5953\ : InMux
    port map (
            O => \N__26713\,
            I => \N__26679\
        );

    \I__5952\ : InMux
    port map (
            O => \N__26712\,
            I => \N__26679\
        );

    \I__5951\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26679\
        );

    \I__5950\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26679\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26676\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__26694\,
            I => \N__26673\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__26679\,
            I => \N__26670\
        );

    \I__5946\ : Span4Mux_v
    port map (
            O => \N__26676\,
            I => \N__26663\
        );

    \I__5945\ : Span4Mux_h
    port map (
            O => \N__26673\,
            I => \N__26663\
        );

    \I__5944\ : Span4Mux_v
    port map (
            O => \N__26670\,
            I => \N__26663\
        );

    \I__5943\ : Sp12to4
    port map (
            O => \N__26663\,
            I => \N__26660\
        );

    \I__5942\ : Span12Mux_h
    port map (
            O => \N__26660\,
            I => \N__26656\
        );

    \I__5941\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26653\
        );

    \I__5940\ : Odrv12
    port map (
            O => \N__26656\,
            I => \eeprom.n2\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__26653\,
            I => \eeprom.n2\
        );

    \I__5938\ : InMux
    port map (
            O => \N__26648\,
            I => \eeprom.n4272\
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__26645\,
            I => \N__26642\
        );

    \I__5936\ : InMux
    port map (
            O => \N__26642\,
            I => \N__26638\
        );

    \I__5935\ : InMux
    port map (
            O => \N__26641\,
            I => \N__26635\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__26638\,
            I => \eeprom.i2c.counter_3\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__26635\,
            I => \eeprom.i2c.counter_3\
        );

    \I__5932\ : CascadeMux
    port map (
            O => \N__26630\,
            I => \N__26627\
        );

    \I__5931\ : InMux
    port map (
            O => \N__26627\,
            I => \N__26623\
        );

    \I__5930\ : InMux
    port map (
            O => \N__26626\,
            I => \N__26620\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__26623\,
            I => \eeprom.i2c.counter_5\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__26620\,
            I => \eeprom.i2c.counter_5\
        );

    \I__5927\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26611\
        );

    \I__5926\ : InMux
    port map (
            O => \N__26614\,
            I => \N__26608\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__26611\,
            I => \eeprom.i2c.counter_4\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__26608\,
            I => \eeprom.i2c.counter_4\
        );

    \I__5923\ : InMux
    port map (
            O => \N__26603\,
            I => \N__26599\
        );

    \I__5922\ : InMux
    port map (
            O => \N__26602\,
            I => \N__26596\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__26599\,
            I => \eeprom.i2c.counter_7\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__26596\,
            I => \eeprom.i2c.counter_7\
        );

    \I__5919\ : InMux
    port map (
            O => \N__26591\,
            I => \N__26587\
        );

    \I__5918\ : InMux
    port map (
            O => \N__26590\,
            I => \N__26584\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__26587\,
            I => \eeprom.i2c.counter_6\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__26584\,
            I => \eeprom.i2c.counter_6\
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__26579\,
            I => \eeprom.i2c.n12_cascade_\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__26576\,
            I => \N__26573\
        );

    \I__5913\ : InMux
    port map (
            O => \N__26573\,
            I => \N__26567\
        );

    \I__5912\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26567\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__26567\,
            I => \eeprom.i2c.n464\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__26564\,
            I => \N__26561\
        );

    \I__5909\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26557\
        );

    \I__5908\ : InMux
    port map (
            O => \N__26560\,
            I => \N__26554\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__26557\,
            I => \N__26551\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__26554\,
            I => \N__26547\
        );

    \I__5905\ : Span4Mux_h
    port map (
            O => \N__26551\,
            I => \N__26544\
        );

    \I__5904\ : InMux
    port map (
            O => \N__26550\,
            I => \N__26541\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__26547\,
            I => n4_adj_358
        );

    \I__5902\ : Odrv4
    port map (
            O => \N__26544\,
            I => n4_adj_358
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__26541\,
            I => n4_adj_358
        );

    \I__5900\ : CascadeMux
    port map (
            O => \N__26534\,
            I => \n10_cascade_\
        );

    \I__5899\ : IoInMux
    port map (
            O => \N__26531\,
            I => \N__26528\
        );

    \I__5898\ : LocalMux
    port map (
            O => \N__26528\,
            I => \N__26525\
        );

    \I__5897\ : Span12Mux_s5_h
    port map (
            O => \N__26525\,
            I => \N__26516\
        );

    \I__5896\ : CascadeMux
    port map (
            O => \N__26524\,
            I => \N__26510\
        );

    \I__5895\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26503\
        );

    \I__5894\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26503\
        );

    \I__5893\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26503\
        );

    \I__5892\ : CascadeMux
    port map (
            O => \N__26520\,
            I => \N__26500\
        );

    \I__5891\ : CascadeMux
    port map (
            O => \N__26519\,
            I => \N__26494\
        );

    \I__5890\ : Span12Mux_v
    port map (
            O => \N__26516\,
            I => \N__26490\
        );

    \I__5889\ : InMux
    port map (
            O => \N__26515\,
            I => \N__26481\
        );

    \I__5888\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26481\
        );

    \I__5887\ : InMux
    port map (
            O => \N__26513\,
            I => \N__26481\
        );

    \I__5886\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26481\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26478\
        );

    \I__5884\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26475\
        );

    \I__5883\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26468\
        );

    \I__5882\ : InMux
    port map (
            O => \N__26498\,
            I => \N__26468\
        );

    \I__5881\ : InMux
    port map (
            O => \N__26497\,
            I => \N__26468\
        );

    \I__5880\ : InMux
    port map (
            O => \N__26494\,
            I => \N__26465\
        );

    \I__5879\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26462\
        );

    \I__5878\ : Odrv12
    port map (
            O => \N__26490\,
            I => \state_7_N_162_3\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__26481\,
            I => \state_7_N_162_3\
        );

    \I__5876\ : Odrv4
    port map (
            O => \N__26478\,
            I => \state_7_N_162_3\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__26475\,
            I => \state_7_N_162_3\
        );

    \I__5874\ : LocalMux
    port map (
            O => \N__26468\,
            I => \state_7_N_162_3\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__26465\,
            I => \state_7_N_162_3\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__26462\,
            I => \state_7_N_162_3\
        );

    \I__5871\ : InMux
    port map (
            O => \N__26447\,
            I => \N__26441\
        );

    \I__5870\ : InMux
    port map (
            O => \N__26446\,
            I => \N__26441\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__26441\,
            I => \eeprom.i2c.n4579\
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__26438\,
            I => \N__26435\
        );

    \I__5867\ : InMux
    port map (
            O => \N__26435\,
            I => \N__26432\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__26432\,
            I => \eeprom.n10\
        );

    \I__5865\ : InMux
    port map (
            O => \N__26429\,
            I => \N__26426\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__26426\,
            I => \N__26423\
        );

    \I__5863\ : Span12Mux_h
    port map (
            O => \N__26423\,
            I => \N__26420\
        );

    \I__5862\ : Odrv12
    port map (
            O => \N__26420\,
            I => \eeprom.n10_adj_343\
        );

    \I__5861\ : InMux
    port map (
            O => \N__26417\,
            I => \eeprom.n4264\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__26414\,
            I => \N__26411\
        );

    \I__5859\ : InMux
    port map (
            O => \N__26411\,
            I => \N__26408\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__26408\,
            I => \eeprom.n9\
        );

    \I__5857\ : CascadeMux
    port map (
            O => \N__26405\,
            I => \N__26402\
        );

    \I__5856\ : InMux
    port map (
            O => \N__26402\,
            I => \N__26399\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__26399\,
            I => \eeprom.n9_adj_308\
        );

    \I__5854\ : InMux
    port map (
            O => \N__26396\,
            I => \bfn_27_26_0_\
        );

    \I__5853\ : InMux
    port map (
            O => \N__26393\,
            I => \N__26390\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26387\
        );

    \I__5851\ : Span4Mux_h
    port map (
            O => \N__26387\,
            I => \N__26384\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__26384\,
            I => \eeprom.n8_adj_311\
        );

    \I__5849\ : InMux
    port map (
            O => \N__26381\,
            I => \eeprom.n4266\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__26378\,
            I => \N__26375\
        );

    \I__5847\ : InMux
    port map (
            O => \N__26375\,
            I => \N__26372\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__26372\,
            I => \eeprom.n7\
        );

    \I__5845\ : InMux
    port map (
            O => \N__26369\,
            I => \eeprom.n4267\
        );

    \I__5844\ : CascadeMux
    port map (
            O => \N__26366\,
            I => \N__26363\
        );

    \I__5843\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26360\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__26360\,
            I => \eeprom.n6\
        );

    \I__5841\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26353\
        );

    \I__5840\ : InMux
    port map (
            O => \N__26356\,
            I => \N__26350\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__26353\,
            I => \N__26345\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__26350\,
            I => \N__26345\
        );

    \I__5837\ : Odrv12
    port map (
            O => \N__26345\,
            I => \eeprom.n6_adj_306\
        );

    \I__5836\ : InMux
    port map (
            O => \N__26342\,
            I => \eeprom.n4268\
        );

    \I__5835\ : CascadeMux
    port map (
            O => \N__26339\,
            I => \N__26336\
        );

    \I__5834\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26333\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__26333\,
            I => \eeprom.n5\
        );

    \I__5832\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26327\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__26327\,
            I => \N__26324\
        );

    \I__5830\ : Odrv12
    port map (
            O => \N__26324\,
            I => \eeprom.n5_adj_317\
        );

    \I__5829\ : InMux
    port map (
            O => \N__26321\,
            I => \eeprom.n4269\
        );

    \I__5828\ : CascadeMux
    port map (
            O => \N__26318\,
            I => \N__26315\
        );

    \I__5827\ : InMux
    port map (
            O => \N__26315\,
            I => \N__26312\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__26312\,
            I => \eeprom.n4\
        );

    \I__5825\ : InMux
    port map (
            O => \N__26309\,
            I => \eeprom.n4270\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__26306\,
            I => \N__26303\
        );

    \I__5823\ : InMux
    port map (
            O => \N__26303\,
            I => \N__26300\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__26300\,
            I => \eeprom.n3\
        );

    \I__5821\ : InMux
    port map (
            O => \N__26297\,
            I => \N__26294\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__26294\,
            I => \N__26291\
        );

    \I__5819\ : Span4Mux_v
    port map (
            O => \N__26291\,
            I => \N__26288\
        );

    \I__5818\ : Odrv4
    port map (
            O => \N__26288\,
            I => \eeprom.n3_adj_312\
        );

    \I__5817\ : InMux
    port map (
            O => \N__26285\,
            I => \eeprom.n4271\
        );

    \I__5816\ : InMux
    port map (
            O => \N__26282\,
            I => \N__26279\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__26279\,
            I => \N__26276\
        );

    \I__5814\ : Span4Mux_h
    port map (
            O => \N__26276\,
            I => \N__26273\
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__26273\,
            I => \eeprom.n18_adj_326\
        );

    \I__5812\ : InMux
    port map (
            O => \N__26270\,
            I => \eeprom.n4256\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__26267\,
            I => \N__26264\
        );

    \I__5810\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26261\
        );

    \I__5809\ : LocalMux
    port map (
            O => \N__26261\,
            I => \eeprom.n17\
        );

    \I__5808\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26255\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__26255\,
            I => \N__26252\
        );

    \I__5806\ : Odrv12
    port map (
            O => \N__26252\,
            I => \eeprom.n17_adj_324\
        );

    \I__5805\ : InMux
    port map (
            O => \N__26249\,
            I => \bfn_27_25_0_\
        );

    \I__5804\ : CascadeMux
    port map (
            O => \N__26246\,
            I => \N__26243\
        );

    \I__5803\ : InMux
    port map (
            O => \N__26243\,
            I => \N__26240\
        );

    \I__5802\ : LocalMux
    port map (
            O => \N__26240\,
            I => \eeprom.n16_adj_294\
        );

    \I__5801\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26234\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__26234\,
            I => \N__26231\
        );

    \I__5799\ : Odrv12
    port map (
            O => \N__26231\,
            I => \eeprom.n16_adj_325\
        );

    \I__5798\ : InMux
    port map (
            O => \N__26228\,
            I => \eeprom.n4258\
        );

    \I__5797\ : CascadeMux
    port map (
            O => \N__26225\,
            I => \N__26222\
        );

    \I__5796\ : InMux
    port map (
            O => \N__26222\,
            I => \N__26219\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__26219\,
            I => \eeprom.n15_adj_295\
        );

    \I__5794\ : InMux
    port map (
            O => \N__26216\,
            I => \N__26213\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__26213\,
            I => \N__26210\
        );

    \I__5792\ : Span4Mux_h
    port map (
            O => \N__26210\,
            I => \N__26207\
        );

    \I__5791\ : Odrv4
    port map (
            O => \N__26207\,
            I => \eeprom.n15\
        );

    \I__5790\ : InMux
    port map (
            O => \N__26204\,
            I => \eeprom.n4259\
        );

    \I__5789\ : InMux
    port map (
            O => \N__26201\,
            I => \N__26198\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__26198\,
            I => \N__26195\
        );

    \I__5787\ : Odrv12
    port map (
            O => \N__26195\,
            I => \eeprom.n14\
        );

    \I__5786\ : InMux
    port map (
            O => \N__26192\,
            I => \eeprom.n4260\
        );

    \I__5785\ : CascadeMux
    port map (
            O => \N__26189\,
            I => \N__26186\
        );

    \I__5784\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26183\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26180\
        );

    \I__5782\ : Span4Mux_v
    port map (
            O => \N__26180\,
            I => \N__26177\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__26177\,
            I => \eeprom.n13\
        );

    \I__5780\ : InMux
    port map (
            O => \N__26174\,
            I => \N__26171\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__26171\,
            I => \N__26168\
        );

    \I__5778\ : Span4Mux_v
    port map (
            O => \N__26168\,
            I => \N__26165\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__26165\,
            I => \eeprom.n13_adj_318\
        );

    \I__5776\ : InMux
    port map (
            O => \N__26162\,
            I => \eeprom.n4261\
        );

    \I__5775\ : CascadeMux
    port map (
            O => \N__26159\,
            I => \N__26156\
        );

    \I__5774\ : InMux
    port map (
            O => \N__26156\,
            I => \N__26153\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__26153\,
            I => \eeprom.n12_adj_298\
        );

    \I__5772\ : InMux
    port map (
            O => \N__26150\,
            I => \N__26147\
        );

    \I__5771\ : LocalMux
    port map (
            O => \N__26147\,
            I => \N__26144\
        );

    \I__5770\ : Span4Mux_v
    port map (
            O => \N__26144\,
            I => \N__26141\
        );

    \I__5769\ : Span4Mux_h
    port map (
            O => \N__26141\,
            I => \N__26138\
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__26138\,
            I => \eeprom.n12_adj_319\
        );

    \I__5767\ : InMux
    port map (
            O => \N__26135\,
            I => \eeprom.n4262\
        );

    \I__5766\ : CascadeMux
    port map (
            O => \N__26132\,
            I => \N__26129\
        );

    \I__5765\ : InMux
    port map (
            O => \N__26129\,
            I => \N__26126\
        );

    \I__5764\ : LocalMux
    port map (
            O => \N__26126\,
            I => \eeprom.n11_adj_299\
        );

    \I__5763\ : InMux
    port map (
            O => \N__26123\,
            I => \N__26120\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__26120\,
            I => \N__26117\
        );

    \I__5761\ : Span4Mux_v
    port map (
            O => \N__26117\,
            I => \N__26114\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__26114\,
            I => \eeprom.n11\
        );

    \I__5759\ : InMux
    port map (
            O => \N__26111\,
            I => \eeprom.n4263\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__26108\,
            I => \N__26105\
        );

    \I__5757\ : InMux
    port map (
            O => \N__26105\,
            I => \N__26102\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26099\
        );

    \I__5755\ : Odrv4
    port map (
            O => \N__26099\,
            I => \eeprom.n26_adj_276\
        );

    \I__5754\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26093\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26090\
        );

    \I__5752\ : Span4Mux_v
    port map (
            O => \N__26090\,
            I => \N__26087\
        );

    \I__5751\ : Odrv4
    port map (
            O => \N__26087\,
            I => \eeprom.n26_adj_275\
        );

    \I__5750\ : InMux
    port map (
            O => \N__26084\,
            I => \eeprom.n4248\
        );

    \I__5749\ : InMux
    port map (
            O => \N__26081\,
            I => \bfn_27_24_0_\
        );

    \I__5748\ : InMux
    port map (
            O => \N__26078\,
            I => \N__26075\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__26075\,
            I => \N__26072\
        );

    \I__5746\ : Span4Mux_h
    port map (
            O => \N__26072\,
            I => \N__26069\
        );

    \I__5745\ : Odrv4
    port map (
            O => \N__26069\,
            I => \eeprom.n24_adj_269\
        );

    \I__5744\ : InMux
    port map (
            O => \N__26066\,
            I => \eeprom.n4250\
        );

    \I__5743\ : CascadeMux
    port map (
            O => \N__26063\,
            I => \N__26060\
        );

    \I__5742\ : InMux
    port map (
            O => \N__26060\,
            I => \N__26057\
        );

    \I__5741\ : LocalMux
    port map (
            O => \N__26057\,
            I => \N__26054\
        );

    \I__5740\ : Odrv4
    port map (
            O => \N__26054\,
            I => \eeprom.n23_adj_268\
        );

    \I__5739\ : InMux
    port map (
            O => \N__26051\,
            I => \N__26048\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__26048\,
            I => \N__26045\
        );

    \I__5737\ : Odrv12
    port map (
            O => \N__26045\,
            I => \eeprom.n23\
        );

    \I__5736\ : InMux
    port map (
            O => \N__26042\,
            I => \eeprom.n4251\
        );

    \I__5735\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26036\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__26036\,
            I => \N__26033\
        );

    \I__5733\ : Span4Mux_h
    port map (
            O => \N__26033\,
            I => \N__26030\
        );

    \I__5732\ : Odrv4
    port map (
            O => \N__26030\,
            I => \eeprom.n22_adj_265\
        );

    \I__5731\ : InMux
    port map (
            O => \N__26027\,
            I => \eeprom.n4252\
        );

    \I__5730\ : CascadeMux
    port map (
            O => \N__26024\,
            I => \N__26021\
        );

    \I__5729\ : InMux
    port map (
            O => \N__26021\,
            I => \N__26018\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__26018\,
            I => \N__26015\
        );

    \I__5727\ : Odrv4
    port map (
            O => \N__26015\,
            I => \eeprom.n21_adj_264\
        );

    \I__5726\ : InMux
    port map (
            O => \N__26012\,
            I => \N__26009\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__26009\,
            I => \N__26006\
        );

    \I__5724\ : Span4Mux_v
    port map (
            O => \N__26006\,
            I => \N__26003\
        );

    \I__5723\ : Odrv4
    port map (
            O => \N__26003\,
            I => \eeprom.n21\
        );

    \I__5722\ : InMux
    port map (
            O => \N__26000\,
            I => \eeprom.n4253\
        );

    \I__5721\ : CascadeMux
    port map (
            O => \N__25997\,
            I => \N__25994\
        );

    \I__5720\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25991\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__25991\,
            I => \N__25988\
        );

    \I__5718\ : Span4Mux_v
    port map (
            O => \N__25988\,
            I => \N__25985\
        );

    \I__5717\ : Odrv4
    port map (
            O => \N__25985\,
            I => \eeprom.n20_adj_259\
        );

    \I__5716\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25979\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__25979\,
            I => \N__25976\
        );

    \I__5714\ : Span4Mux_h
    port map (
            O => \N__25976\,
            I => \N__25973\
        );

    \I__5713\ : Odrv4
    port map (
            O => \N__25973\,
            I => \eeprom.n20\
        );

    \I__5712\ : InMux
    port map (
            O => \N__25970\,
            I => \eeprom.n4254\
        );

    \I__5711\ : InMux
    port map (
            O => \N__25967\,
            I => \N__25964\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__25964\,
            I => \N__25961\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__25961\,
            I => \N__25958\
        );

    \I__5708\ : Odrv4
    port map (
            O => \N__25958\,
            I => \eeprom.n19_adj_320\
        );

    \I__5707\ : InMux
    port map (
            O => \N__25955\,
            I => \eeprom.n4255\
        );

    \I__5706\ : CascadeMux
    port map (
            O => \N__25952\,
            I => \eeprom.n1138_cascade_\
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__25949\,
            I => \N__25946\
        );

    \I__5704\ : InMux
    port map (
            O => \N__25946\,
            I => \N__25943\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__25943\,
            I => \N__25940\
        );

    \I__5702\ : Odrv4
    port map (
            O => \N__25940\,
            I => \eeprom.n33_adj_289\
        );

    \I__5701\ : InMux
    port map (
            O => \N__25937\,
            I => \N__25934\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__25934\,
            I => \N__25931\
        );

    \I__5699\ : Odrv12
    port map (
            O => \N__25931\,
            I => \eeprom.n33\
        );

    \I__5698\ : InMux
    port map (
            O => \N__25928\,
            I => \bfn_27_23_0_\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__25925\,
            I => \N__25922\
        );

    \I__5696\ : InMux
    port map (
            O => \N__25922\,
            I => \N__25919\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__25919\,
            I => \eeprom.n32_adj_288\
        );

    \I__5694\ : InMux
    port map (
            O => \N__25916\,
            I => \N__25913\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__25913\,
            I => \N__25910\
        );

    \I__5692\ : Span4Mux_v
    port map (
            O => \N__25910\,
            I => \N__25907\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__25907\,
            I => \N__25904\
        );

    \I__5690\ : Odrv4
    port map (
            O => \N__25904\,
            I => \eeprom.n32_adj_287\
        );

    \I__5689\ : InMux
    port map (
            O => \N__25901\,
            I => \eeprom.n4242\
        );

    \I__5688\ : CascadeMux
    port map (
            O => \N__25898\,
            I => \N__25895\
        );

    \I__5687\ : InMux
    port map (
            O => \N__25895\,
            I => \N__25892\
        );

    \I__5686\ : LocalMux
    port map (
            O => \N__25892\,
            I => \N__25889\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__25889\,
            I => \N__25886\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__25886\,
            I => \eeprom.n31_adj_286\
        );

    \I__5683\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25880\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__25880\,
            I => \N__25877\
        );

    \I__5681\ : Span4Mux_v
    port map (
            O => \N__25877\,
            I => \N__25874\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__25874\,
            I => \eeprom.n31_adj_285\
        );

    \I__5679\ : InMux
    port map (
            O => \N__25871\,
            I => \eeprom.n4243\
        );

    \I__5678\ : InMux
    port map (
            O => \N__25868\,
            I => \N__25865\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__25865\,
            I => \N__25862\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__25862\,
            I => \eeprom.n30_adj_277\
        );

    \I__5675\ : InMux
    port map (
            O => \N__25859\,
            I => \N__25856\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__25856\,
            I => \N__25853\
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__25853\,
            I => \eeprom.n30_adj_284\
        );

    \I__5672\ : InMux
    port map (
            O => \N__25850\,
            I => \eeprom.n4244\
        );

    \I__5671\ : CascadeMux
    port map (
            O => \N__25847\,
            I => \N__25844\
        );

    \I__5670\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25841\
        );

    \I__5669\ : LocalMux
    port map (
            O => \N__25841\,
            I => \N__25838\
        );

    \I__5668\ : Odrv4
    port map (
            O => \N__25838\,
            I => \eeprom.n29_adj_278\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__25835\,
            I => \N__25832\
        );

    \I__5666\ : InMux
    port map (
            O => \N__25832\,
            I => \N__25829\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__25829\,
            I => \N__25826\
        );

    \I__5664\ : Span4Mux_v
    port map (
            O => \N__25826\,
            I => \N__25823\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__25823\,
            I => \eeprom.n29_adj_283\
        );

    \I__5662\ : InMux
    port map (
            O => \N__25820\,
            I => \eeprom.n4245\
        );

    \I__5661\ : CascadeMux
    port map (
            O => \N__25817\,
            I => \N__25814\
        );

    \I__5660\ : InMux
    port map (
            O => \N__25814\,
            I => \N__25811\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__25811\,
            I => \N__25808\
        );

    \I__5658\ : Span4Mux_v
    port map (
            O => \N__25808\,
            I => \N__25805\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__25805\,
            I => \eeprom.n28_adj_279\
        );

    \I__5656\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25799\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__25799\,
            I => \N__25796\
        );

    \I__5654\ : Span4Mux_h
    port map (
            O => \N__25796\,
            I => \N__25793\
        );

    \I__5653\ : Span4Mux_v
    port map (
            O => \N__25793\,
            I => \N__25790\
        );

    \I__5652\ : Odrv4
    port map (
            O => \N__25790\,
            I => \eeprom.n28_adj_282\
        );

    \I__5651\ : InMux
    port map (
            O => \N__25787\,
            I => \eeprom.n4246\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__25784\,
            I => \N__25781\
        );

    \I__5649\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25778\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__25778\,
            I => \eeprom.n27_adj_280\
        );

    \I__5647\ : InMux
    port map (
            O => \N__25775\,
            I => \eeprom.n4247\
        );

    \I__5646\ : InMux
    port map (
            O => \N__25772\,
            I => \N__25769\
        );

    \I__5645\ : LocalMux
    port map (
            O => \N__25769\,
            I => \N__25766\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__25766\,
            I => \N__25763\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__25763\,
            I => \N__25757\
        );

    \I__5642\ : InMux
    port map (
            O => \N__25762\,
            I => \N__25754\
        );

    \I__5641\ : InMux
    port map (
            O => \N__25761\,
            I => \N__25751\
        );

    \I__5640\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25748\
        );

    \I__5639\ : Odrv4
    port map (
            O => \N__25757\,
            I => \eeprom.eeprom_counter_3\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__25754\,
            I => \eeprom.eeprom_counter_3\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__25751\,
            I => \eeprom.eeprom_counter_3\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__25748\,
            I => \eeprom.eeprom_counter_3\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__25739\,
            I => \N__25736\
        );

    \I__5634\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25732\
        );

    \I__5633\ : InMux
    port map (
            O => \N__25735\,
            I => \N__25729\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__25732\,
            I => \N__25726\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__25729\,
            I => \N__25723\
        );

    \I__5630\ : Span4Mux_v
    port map (
            O => \N__25726\,
            I => \N__25719\
        );

    \I__5629\ : Span4Mux_h
    port map (
            O => \N__25723\,
            I => \N__25716\
        );

    \I__5628\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25713\
        );

    \I__5627\ : Odrv4
    port map (
            O => \N__25719\,
            I => \eeprom.n1916\
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__25716\,
            I => \eeprom.n1916\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__25713\,
            I => \eeprom.n1916\
        );

    \I__5624\ : CascadeMux
    port map (
            O => \N__25706\,
            I => \eeprom.n5035_cascade_\
        );

    \I__5623\ : InMux
    port map (
            O => \N__25703\,
            I => \N__25700\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__25700\,
            I => \N__25697\
        );

    \I__5621\ : Span4Mux_h
    port map (
            O => \N__25697\,
            I => \N__25694\
        );

    \I__5620\ : Odrv4
    port map (
            O => \N__25694\,
            I => \eeprom.n5039\
        );

    \I__5619\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25688\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__25688\,
            I => \N__25684\
        );

    \I__5617\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25680\
        );

    \I__5616\ : Span4Mux_v
    port map (
            O => \N__25684\,
            I => \N__25677\
        );

    \I__5615\ : InMux
    port map (
            O => \N__25683\,
            I => \N__25674\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__25680\,
            I => \eeprom.eeprom_counter_12\
        );

    \I__5613\ : Odrv4
    port map (
            O => \N__25677\,
            I => \eeprom.eeprom_counter_12\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__25674\,
            I => \eeprom.eeprom_counter_12\
        );

    \I__5611\ : InMux
    port map (
            O => \N__25667\,
            I => \N__25664\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__25664\,
            I => \N__25660\
        );

    \I__5609\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25657\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__25660\,
            I => \N__25654\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__25657\,
            I => \N__25650\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__25654\,
            I => \N__25646\
        );

    \I__5605\ : InMux
    port map (
            O => \N__25653\,
            I => \N__25643\
        );

    \I__5604\ : Span4Mux_h
    port map (
            O => \N__25650\,
            I => \N__25640\
        );

    \I__5603\ : InMux
    port map (
            O => \N__25649\,
            I => \N__25637\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__25646\,
            I => \eeprom.eeprom_counter_1\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__25643\,
            I => \eeprom.eeprom_counter_1\
        );

    \I__5600\ : Odrv4
    port map (
            O => \N__25640\,
            I => \eeprom.eeprom_counter_1\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__25637\,
            I => \eeprom.eeprom_counter_1\
        );

    \I__5598\ : CascadeMux
    port map (
            O => \N__25628\,
            I => \eeprom.n892_cascade_\
        );

    \I__5597\ : InMux
    port map (
            O => \N__25625\,
            I => \N__25622\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__25622\,
            I => \N__25618\
        );

    \I__5595\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25614\
        );

    \I__5594\ : Span12Mux_h
    port map (
            O => \N__25618\,
            I => \N__25611\
        );

    \I__5593\ : InMux
    port map (
            O => \N__25617\,
            I => \N__25608\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__25614\,
            I => \eeprom.eeprom_counter_10\
        );

    \I__5591\ : Odrv12
    port map (
            O => \N__25611\,
            I => \eeprom.eeprom_counter_10\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__25608\,
            I => \eeprom.eeprom_counter_10\
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__25601\,
            I => \N__25597\
        );

    \I__5588\ : CascadeMux
    port map (
            O => \N__25600\,
            I => \N__25594\
        );

    \I__5587\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25590\
        );

    \I__5586\ : InMux
    port map (
            O => \N__25594\,
            I => \N__25587\
        );

    \I__5585\ : InMux
    port map (
            O => \N__25593\,
            I => \N__25584\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__25590\,
            I => \N__25581\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__25587\,
            I => \N__25578\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__25584\,
            I => \eeprom.eeprom_counter_28\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__25581\,
            I => \eeprom.eeprom_counter_28\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__25578\,
            I => \eeprom.eeprom_counter_28\
        );

    \I__5579\ : CascadeMux
    port map (
            O => \N__25571\,
            I => \eeprom.n1256_cascade_\
        );

    \I__5578\ : InMux
    port map (
            O => \N__25568\,
            I => \N__25565\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__25565\,
            I => \N__25561\
        );

    \I__5576\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25558\
        );

    \I__5575\ : Span4Mux_v
    port map (
            O => \N__25561\,
            I => \N__25553\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__25558\,
            I => \N__25553\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__25553\,
            I => \eeprom.n1913\
        );

    \I__5572\ : InMux
    port map (
            O => \N__25550\,
            I => \N__25547\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__25547\,
            I => \eeprom.i2c.n13\
        );

    \I__5570\ : InMux
    port map (
            O => \N__25544\,
            I => \N__25541\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__25541\,
            I => \N__25537\
        );

    \I__5568\ : InMux
    port map (
            O => \N__25540\,
            I => \N__25533\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__25537\,
            I => \N__25530\
        );

    \I__5566\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25527\
        );

    \I__5565\ : LocalMux
    port map (
            O => \N__25533\,
            I => \eeprom.eeprom_counter_7\
        );

    \I__5564\ : Odrv4
    port map (
            O => \N__25530\,
            I => \eeprom.eeprom_counter_7\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__25527\,
            I => \eeprom.eeprom_counter_7\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__25520\,
            I => \N__25516\
        );

    \I__5561\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25510\
        );

    \I__5560\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25510\
        );

    \I__5559\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25507\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__25510\,
            I => \N__25502\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__25507\,
            I => \N__25502\
        );

    \I__5556\ : Span4Mux_v
    port map (
            O => \N__25502\,
            I => \N__25499\
        );

    \I__5555\ : Odrv4
    port map (
            O => \N__25499\,
            I => \eeprom.n1918\
        );

    \I__5554\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25493\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__25493\,
            I => \N__25490\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__25490\,
            I => \N__25486\
        );

    \I__5551\ : CascadeMux
    port map (
            O => \N__25489\,
            I => \N__25481\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__25486\,
            I => \N__25478\
        );

    \I__5549\ : InMux
    port map (
            O => \N__25485\,
            I => \N__25475\
        );

    \I__5548\ : InMux
    port map (
            O => \N__25484\,
            I => \N__25472\
        );

    \I__5547\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25469\
        );

    \I__5546\ : Odrv4
    port map (
            O => \N__25478\,
            I => \eeprom.eeprom_counter_0\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__25475\,
            I => \eeprom.eeprom_counter_0\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__25472\,
            I => \eeprom.eeprom_counter_0\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__25469\,
            I => \eeprom.eeprom_counter_0\
        );

    \I__5542\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25456\
        );

    \I__5541\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25453\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__25456\,
            I => \N__25448\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__25453\,
            I => \N__25448\
        );

    \I__5538\ : Span4Mux_v
    port map (
            O => \N__25448\,
            I => \N__25445\
        );

    \I__5537\ : Odrv4
    port map (
            O => \N__25445\,
            I => \eeprom.n1912\
        );

    \I__5536\ : InMux
    port map (
            O => \N__25442\,
            I => \N__25439\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__25439\,
            I => \N__25435\
        );

    \I__5534\ : InMux
    port map (
            O => \N__25438\,
            I => \N__25431\
        );

    \I__5533\ : Span4Mux_h
    port map (
            O => \N__25435\,
            I => \N__25428\
        );

    \I__5532\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25425\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__25431\,
            I => \eeprom.eeprom_counter_27\
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__25428\,
            I => \eeprom.eeprom_counter_27\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__25425\,
            I => \eeprom.eeprom_counter_27\
        );

    \I__5528\ : CascadeMux
    port map (
            O => \N__25418\,
            I => \eeprom.n1139_cascade_\
        );

    \I__5527\ : InMux
    port map (
            O => \N__25415\,
            I => \N__25411\
        );

    \I__5526\ : InMux
    port map (
            O => \N__25414\,
            I => \N__25408\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__25411\,
            I => \eeprom.i2c.n37\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__25408\,
            I => \eeprom.i2c.n37\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__25403\,
            I => \eeprom.i2c.n37_cascade_\
        );

    \I__5522\ : InMux
    port map (
            O => \N__25400\,
            I => \N__25394\
        );

    \I__5521\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25394\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__25394\,
            I => \eeprom.i2c.n33\
        );

    \I__5519\ : CascadeMux
    port map (
            O => \N__25391\,
            I => \eeprom.i2c.n39_cascade_\
        );

    \I__5518\ : InMux
    port map (
            O => \N__25388\,
            I => \N__25385\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__25385\,
            I => \eeprom.i2c.n39\
        );

    \I__5516\ : CascadeMux
    port map (
            O => \N__25382\,
            I => \eeprom.i2c.n407_cascade_\
        );

    \I__5515\ : CascadeMux
    port map (
            O => \N__25379\,
            I => \N__25376\
        );

    \I__5514\ : InMux
    port map (
            O => \N__25376\,
            I => \N__25373\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__25373\,
            I => \N__25370\
        );

    \I__5512\ : Span4Mux_h
    port map (
            O => \N__25370\,
            I => \N__25367\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__25367\,
            I => \N__25364\
        );

    \I__5510\ : Odrv4
    port map (
            O => \N__25364\,
            I => \eeprom.n917\
        );

    \I__5509\ : InMux
    port map (
            O => \N__25361\,
            I => \N__25357\
        );

    \I__5508\ : InMux
    port map (
            O => \N__25360\,
            I => \N__25354\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__25357\,
            I => \N__25351\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__25354\,
            I => \N__25348\
        );

    \I__5505\ : Span4Mux_h
    port map (
            O => \N__25351\,
            I => \N__25345\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__25348\,
            I => \N__25341\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__25345\,
            I => \N__25337\
        );

    \I__5502\ : InMux
    port map (
            O => \N__25344\,
            I => \N__25334\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__25341\,
            I => \N__25331\
        );

    \I__5500\ : InMux
    port map (
            O => \N__25340\,
            I => \N__25328\
        );

    \I__5499\ : Odrv4
    port map (
            O => \N__25337\,
            I => \eeprom.eeprom_counter_5\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__25334\,
            I => \eeprom.eeprom_counter_5\
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__25331\,
            I => \eeprom.eeprom_counter_5\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__25328\,
            I => \eeprom.eeprom_counter_5\
        );

    \I__5495\ : InMux
    port map (
            O => \N__25319\,
            I => \N__25316\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__25316\,
            I => \N__25313\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__25313\,
            I => \N__25310\
        );

    \I__5492\ : Span4Mux_h
    port map (
            O => \N__25310\,
            I => \N__25307\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__25307\,
            I => \eeprom.n3722\
        );

    \I__5490\ : InMux
    port map (
            O => \N__25304\,
            I => \N__25301\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__25301\,
            I => \N__25297\
        );

    \I__5488\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25293\
        );

    \I__5487\ : Span4Mux_v
    port map (
            O => \N__25297\,
            I => \N__25290\
        );

    \I__5486\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25287\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__25293\,
            I => \eeprom.eeprom_counter_30\
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__25290\,
            I => \eeprom.eeprom_counter_30\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__25287\,
            I => \eeprom.eeprom_counter_30\
        );

    \I__5482\ : InMux
    port map (
            O => \N__25280\,
            I => \N__25277\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__25277\,
            I => n4733
        );

    \I__5480\ : SRMux
    port map (
            O => \N__25274\,
            I => \N__25271\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__25271\,
            I => \N__25268\
        );

    \I__5478\ : Span4Mux_h
    port map (
            O => \N__25268\,
            I => \N__25265\
        );

    \I__5477\ : Odrv4
    port map (
            O => \N__25265\,
            I => \eeprom.i2c.n1913\
        );

    \I__5476\ : InMux
    port map (
            O => \N__25262\,
            I => \N__25259\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__25259\,
            I => \eeprom.i2c.n534\
        );

    \I__5474\ : CEMux
    port map (
            O => \N__25256\,
            I => \N__25253\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__25253\,
            I => \N__25250\
        );

    \I__5472\ : Odrv12
    port map (
            O => \N__25250\,
            I => \eeprom.i2c.n1829\
        );

    \I__5471\ : InMux
    port map (
            O => \N__25247\,
            I => \N__25241\
        );

    \I__5470\ : InMux
    port map (
            O => \N__25246\,
            I => \N__25236\
        );

    \I__5469\ : InMux
    port map (
            O => \N__25245\,
            I => \N__25236\
        );

    \I__5468\ : InMux
    port map (
            O => \N__25244\,
            I => \N__25233\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__25241\,
            I => \eeprom.i2c.n9\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__25236\,
            I => \eeprom.i2c.n9\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__25233\,
            I => \eeprom.i2c.n9\
        );

    \I__5464\ : CascadeMux
    port map (
            O => \N__25226\,
            I => \eeprom.i2c.n9_cascade_\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__25223\,
            I => \N__25220\
        );

    \I__5462\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25217\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__25217\,
            I => \N__25214\
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__25214\,
            I => n1814
        );

    \I__5459\ : CascadeMux
    port map (
            O => \N__25211\,
            I => \n1814_cascade_\
        );

    \I__5458\ : InMux
    port map (
            O => \N__25208\,
            I => \bfn_27_17_0_\
        );

    \I__5457\ : InMux
    port map (
            O => \N__25205\,
            I => \eeprom.i2c.n3899\
        );

    \I__5456\ : InMux
    port map (
            O => \N__25202\,
            I => \eeprom.i2c.n3900\
        );

    \I__5455\ : InMux
    port map (
            O => \N__25199\,
            I => \eeprom.i2c.n3901\
        );

    \I__5454\ : InMux
    port map (
            O => \N__25196\,
            I => \eeprom.i2c.n3902\
        );

    \I__5453\ : InMux
    port map (
            O => \N__25193\,
            I => \eeprom.i2c.n3903\
        );

    \I__5452\ : InMux
    port map (
            O => \N__25190\,
            I => \eeprom.i2c.n3904\
        );

    \I__5451\ : InMux
    port map (
            O => \N__25187\,
            I => \eeprom.i2c.n3905\
        );

    \I__5450\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25179\
        );

    \I__5449\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25174\
        );

    \I__5448\ : InMux
    port map (
            O => \N__25182\,
            I => \N__25174\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__25179\,
            I => n11
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__25174\,
            I => n11
        );

    \I__5445\ : InMux
    port map (
            O => \N__25169\,
            I => \N__25161\
        );

    \I__5444\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25161\
        );

    \I__5443\ : InMux
    port map (
            O => \N__25167\,
            I => \N__25158\
        );

    \I__5442\ : InMux
    port map (
            O => \N__25166\,
            I => \N__25155\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__25161\,
            I => \N__25152\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__25158\,
            I => n10_adj_360
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__25155\,
            I => n10_adj_360
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__25152\,
            I => n10_adj_360
        );

    \I__5437\ : InMux
    port map (
            O => \N__25145\,
            I => \N__25140\
        );

    \I__5436\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25137\
        );

    \I__5435\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25134\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__25140\,
            I => \N__25127\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__25137\,
            I => \N__25127\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__25134\,
            I => \N__25127\
        );

    \I__5431\ : Span12Mux_v
    port map (
            O => \N__25127\,
            I => \N__25124\
        );

    \I__5430\ : Odrv12
    port map (
            O => \N__25124\,
            I => \eeprom.n1919\
        );

    \I__5429\ : CascadeMux
    port map (
            O => \N__25121\,
            I => \N__25116\
        );

    \I__5428\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25113\
        );

    \I__5427\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25108\
        );

    \I__5426\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25108\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__25113\,
            I => \eeprom.eeprom_counter_24\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__25108\,
            I => \eeprom.eeprom_counter_24\
        );

    \I__5423\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25099\
        );

    \I__5422\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25095\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__25099\,
            I => \N__25092\
        );

    \I__5420\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25089\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__25095\,
            I => \N__25084\
        );

    \I__5418\ : Span4Mux_v
    port map (
            O => \N__25092\,
            I => \N__25084\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__25089\,
            I => \N__25081\
        );

    \I__5416\ : Odrv4
    port map (
            O => \N__25084\,
            I => \eeprom.eeprom_counter_18\
        );

    \I__5415\ : Odrv4
    port map (
            O => \N__25081\,
            I => \eeprom.eeprom_counter_18\
        );

    \I__5414\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25073\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__25073\,
            I => \N__25068\
        );

    \I__5412\ : InMux
    port map (
            O => \N__25072\,
            I => \N__25065\
        );

    \I__5411\ : InMux
    port map (
            O => \N__25071\,
            I => \N__25062\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__25068\,
            I => \N__25059\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__25065\,
            I => \N__25056\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__25062\,
            I => \eeprom.eeprom_counter_17\
        );

    \I__5407\ : Odrv4
    port map (
            O => \N__25059\,
            I => \eeprom.eeprom_counter_17\
        );

    \I__5406\ : Odrv12
    port map (
            O => \N__25056\,
            I => \eeprom.eeprom_counter_17\
        );

    \I__5405\ : InMux
    port map (
            O => \N__25049\,
            I => \N__25046\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__25046\,
            I => \N__25041\
        );

    \I__5403\ : InMux
    port map (
            O => \N__25045\,
            I => \N__25038\
        );

    \I__5402\ : InMux
    port map (
            O => \N__25044\,
            I => \N__25035\
        );

    \I__5401\ : Span4Mux_v
    port map (
            O => \N__25041\,
            I => \N__25030\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25030\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__25035\,
            I => \eeprom.eeprom_counter_22\
        );

    \I__5398\ : Odrv4
    port map (
            O => \N__25030\,
            I => \eeprom.eeprom_counter_22\
        );

    \I__5397\ : InMux
    port map (
            O => \N__25025\,
            I => \N__25022\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__25022\,
            I => \N__25017\
        );

    \I__5395\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25014\
        );

    \I__5394\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25011\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__25017\,
            I => \N__25008\
        );

    \I__5392\ : LocalMux
    port map (
            O => \N__25014\,
            I => \N__25005\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__25011\,
            I => \eeprom.eeprom_counter_21\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__25008\,
            I => \eeprom.eeprom_counter_21\
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__25005\,
            I => \eeprom.eeprom_counter_21\
        );

    \I__5388\ : InMux
    port map (
            O => \N__24998\,
            I => \eeprom.n3957\
        );

    \I__5387\ : InMux
    port map (
            O => \N__24995\,
            I => \eeprom.n3958\
        );

    \I__5386\ : InMux
    port map (
            O => \N__24992\,
            I => \eeprom.n3959\
        );

    \I__5385\ : InMux
    port map (
            O => \N__24989\,
            I => \eeprom.n3960\
        );

    \I__5384\ : InMux
    port map (
            O => \N__24986\,
            I => \eeprom.n3961\
        );

    \I__5383\ : InMux
    port map (
            O => \N__24983\,
            I => \N__24980\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__24980\,
            I => \N__24975\
        );

    \I__5381\ : InMux
    port map (
            O => \N__24979\,
            I => \N__24972\
        );

    \I__5380\ : InMux
    port map (
            O => \N__24978\,
            I => \N__24969\
        );

    \I__5379\ : Span4Mux_h
    port map (
            O => \N__24975\,
            I => \N__24966\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__24972\,
            I => \N__24963\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__24969\,
            I => \eeprom.eeprom_counter_23\
        );

    \I__5376\ : Odrv4
    port map (
            O => \N__24966\,
            I => \eeprom.eeprom_counter_23\
        );

    \I__5375\ : Odrv4
    port map (
            O => \N__24963\,
            I => \eeprom.eeprom_counter_23\
        );

    \I__5374\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24952\
        );

    \I__5373\ : CascadeMux
    port map (
            O => \N__24955\,
            I => \N__24949\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__24952\,
            I => \N__24945\
        );

    \I__5371\ : InMux
    port map (
            O => \N__24949\,
            I => \N__24942\
        );

    \I__5370\ : InMux
    port map (
            O => \N__24948\,
            I => \N__24939\
        );

    \I__5369\ : Span4Mux_h
    port map (
            O => \N__24945\,
            I => \N__24936\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__24942\,
            I => \N__24933\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__24939\,
            I => \eeprom.eeprom_counter_16\
        );

    \I__5366\ : Odrv4
    port map (
            O => \N__24936\,
            I => \eeprom.eeprom_counter_16\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__24933\,
            I => \eeprom.eeprom_counter_16\
        );

    \I__5364\ : InMux
    port map (
            O => \N__24926\,
            I => \eeprom.n3948\
        );

    \I__5363\ : InMux
    port map (
            O => \N__24923\,
            I => \eeprom.n3949\
        );

    \I__5362\ : CascadeMux
    port map (
            O => \N__24920\,
            I => \N__24916\
        );

    \I__5361\ : InMux
    port map (
            O => \N__24919\,
            I => \N__24912\
        );

    \I__5360\ : InMux
    port map (
            O => \N__24916\,
            I => \N__24909\
        );

    \I__5359\ : InMux
    port map (
            O => \N__24915\,
            I => \N__24906\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__24912\,
            I => \N__24903\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__24909\,
            I => \N__24900\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__24906\,
            I => \eeprom.eeprom_counter_20\
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__24903\,
            I => \eeprom.eeprom_counter_20\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__24900\,
            I => \eeprom.eeprom_counter_20\
        );

    \I__5353\ : InMux
    port map (
            O => \N__24893\,
            I => \eeprom.n3950\
        );

    \I__5352\ : InMux
    port map (
            O => \N__24890\,
            I => \eeprom.n3951\
        );

    \I__5351\ : InMux
    port map (
            O => \N__24887\,
            I => \eeprom.n3952\
        );

    \I__5350\ : InMux
    port map (
            O => \N__24884\,
            I => \eeprom.n3953\
        );

    \I__5349\ : InMux
    port map (
            O => \N__24881\,
            I => \bfn_26_24_0_\
        );

    \I__5348\ : InMux
    port map (
            O => \N__24878\,
            I => \eeprom.n3955\
        );

    \I__5347\ : InMux
    port map (
            O => \N__24875\,
            I => \eeprom.n3956\
        );

    \I__5346\ : InMux
    port map (
            O => \N__24872\,
            I => \eeprom.n3939\
        );

    \I__5345\ : InMux
    port map (
            O => \N__24869\,
            I => \eeprom.n3940\
        );

    \I__5344\ : InMux
    port map (
            O => \N__24866\,
            I => \eeprom.n3941\
        );

    \I__5343\ : InMux
    port map (
            O => \N__24863\,
            I => \eeprom.n3942\
        );

    \I__5342\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24857\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__24857\,
            I => \N__24852\
        );

    \I__5340\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24849\
        );

    \I__5339\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24846\
        );

    \I__5338\ : Span4Mux_v
    port map (
            O => \N__24852\,
            I => \N__24843\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24840\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__24846\,
            I => \eeprom.eeprom_counter_13\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__24843\,
            I => \eeprom.eeprom_counter_13\
        );

    \I__5334\ : Odrv4
    port map (
            O => \N__24840\,
            I => \eeprom.eeprom_counter_13\
        );

    \I__5333\ : InMux
    port map (
            O => \N__24833\,
            I => \eeprom.n3943\
        );

    \I__5332\ : InMux
    port map (
            O => \N__24830\,
            I => \eeprom.n3944\
        );

    \I__5331\ : InMux
    port map (
            O => \N__24827\,
            I => \eeprom.n3945\
        );

    \I__5330\ : InMux
    port map (
            O => \N__24824\,
            I => \bfn_26_23_0_\
        );

    \I__5329\ : InMux
    port map (
            O => \N__24821\,
            I => \eeprom.n3947\
        );

    \I__5328\ : InMux
    port map (
            O => \N__24818\,
            I => \bfn_26_21_0_\
        );

    \I__5327\ : InMux
    port map (
            O => \N__24815\,
            I => \eeprom.n3931\
        );

    \I__5326\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24805\
        );

    \I__5324\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24802\
        );

    \I__5323\ : Span4Mux_h
    port map (
            O => \N__24805\,
            I => \N__24799\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__24802\,
            I => \N__24795\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__24799\,
            I => \N__24791\
        );

    \I__5320\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24788\
        );

    \I__5319\ : Span4Mux_h
    port map (
            O => \N__24795\,
            I => \N__24785\
        );

    \I__5318\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24782\
        );

    \I__5317\ : Odrv4
    port map (
            O => \N__24791\,
            I => \eeprom.eeprom_counter_2\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__24788\,
            I => \eeprom.eeprom_counter_2\
        );

    \I__5315\ : Odrv4
    port map (
            O => \N__24785\,
            I => \eeprom.eeprom_counter_2\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__24782\,
            I => \eeprom.eeprom_counter_2\
        );

    \I__5313\ : InMux
    port map (
            O => \N__24773\,
            I => \eeprom.n3932\
        );

    \I__5312\ : InMux
    port map (
            O => \N__24770\,
            I => \eeprom.n3933\
        );

    \I__5311\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24764\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__24764\,
            I => \N__24760\
        );

    \I__5309\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24757\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__24760\,
            I => \N__24754\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24750\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__24754\,
            I => \N__24746\
        );

    \I__5305\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24743\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__24750\,
            I => \N__24740\
        );

    \I__5303\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24737\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__24746\,
            I => \eeprom.eeprom_counter_4\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__24743\,
            I => \eeprom.eeprom_counter_4\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__24740\,
            I => \eeprom.eeprom_counter_4\
        );

    \I__5299\ : LocalMux
    port map (
            O => \N__24737\,
            I => \eeprom.eeprom_counter_4\
        );

    \I__5298\ : InMux
    port map (
            O => \N__24728\,
            I => \eeprom.n3934\
        );

    \I__5297\ : InMux
    port map (
            O => \N__24725\,
            I => \eeprom.n3935\
        );

    \I__5296\ : InMux
    port map (
            O => \N__24722\,
            I => \eeprom.n3936\
        );

    \I__5295\ : InMux
    port map (
            O => \N__24719\,
            I => \eeprom.n3937\
        );

    \I__5294\ : InMux
    port map (
            O => \N__24716\,
            I => \bfn_26_22_0_\
        );

    \I__5293\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24709\
        );

    \I__5292\ : InMux
    port map (
            O => \N__24712\,
            I => \N__24706\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__24709\,
            I => \N__24700\
        );

    \I__5290\ : LocalMux
    port map (
            O => \N__24706\,
            I => \N__24700\
        );

    \I__5289\ : InMux
    port map (
            O => \N__24705\,
            I => \N__24697\
        );

    \I__5288\ : Odrv4
    port map (
            O => \N__24700\,
            I => n1805
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__24697\,
            I => n1805
        );

    \I__5286\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24689\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__24689\,
            I => n158
        );

    \I__5284\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24683\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__24683\,
            I => n8
        );

    \I__5282\ : CascadeMux
    port map (
            O => \N__24680\,
            I => \n5461_cascade_\
        );

    \I__5281\ : InMux
    port map (
            O => \N__24677\,
            I => \N__24671\
        );

    \I__5280\ : InMux
    port map (
            O => \N__24676\,
            I => \N__24671\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__24671\,
            I => \N__24667\
        );

    \I__5278\ : InMux
    port map (
            O => \N__24670\,
            I => \N__24664\
        );

    \I__5277\ : Odrv4
    port map (
            O => \N__24667\,
            I => n1800
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__24664\,
            I => n1800
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__24659\,
            I => \N__24655\
        );

    \I__5274\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24650\
        );

    \I__5273\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24650\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__24650\,
            I => \N__24647\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__24647\,
            I => n3585
        );

    \I__5270\ : InMux
    port map (
            O => \N__24644\,
            I => \N__24641\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__24641\,
            I => n160
        );

    \I__5268\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24635\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__24635\,
            I => \N__24630\
        );

    \I__5266\ : InMux
    port map (
            O => \N__24634\,
            I => \N__24627\
        );

    \I__5265\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24624\
        );

    \I__5264\ : Span4Mux_h
    port map (
            O => \N__24630\,
            I => \N__24619\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__24627\,
            I => \N__24619\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__24624\,
            I => \N__24616\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__24619\,
            I => \N__24613\
        );

    \I__5260\ : Span4Mux_h
    port map (
            O => \N__24616\,
            I => \N__24610\
        );

    \I__5259\ : Span4Mux_h
    port map (
            O => \N__24613\,
            I => \N__24607\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__24610\,
            I => \eeprom.n2119\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__24607\,
            I => \eeprom.n2119\
        );

    \I__5256\ : InMux
    port map (
            O => \N__24602\,
            I => \N__24597\
        );

    \I__5255\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24594\
        );

    \I__5254\ : InMux
    port map (
            O => \N__24600\,
            I => \N__24591\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__24597\,
            I => \N__24584\
        );

    \I__5252\ : LocalMux
    port map (
            O => \N__24594\,
            I => \N__24584\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__24591\,
            I => \N__24584\
        );

    \I__5250\ : Odrv12
    port map (
            O => \N__24584\,
            I => \eeprom.n2319\
        );

    \I__5249\ : InMux
    port map (
            O => \N__24581\,
            I => \N__24578\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__24578\,
            I => n172
        );

    \I__5247\ : CascadeMux
    port map (
            O => \N__24575\,
            I => \n22_adj_367_cascade_\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__24572\,
            I => \n4_adj_369_cascade_\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__24569\,
            I => \n4_cascade_\
        );

    \I__5244\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24563\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__24563\,
            I => n166
        );

    \I__5242\ : CascadeMux
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__5241\ : InMux
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__24554\,
            I => n4
        );

    \I__5239\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24548\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__24548\,
            I => n168
        );

    \I__5237\ : CascadeMux
    port map (
            O => \N__24545\,
            I => \n1805_cascade_\
        );

    \I__5236\ : InMux
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__5235\ : LocalMux
    port map (
            O => \N__24539\,
            I => n170
        );

    \I__5234\ : CascadeMux
    port map (
            O => \N__24536\,
            I => \n1800_cascade_\
        );

    \I__5233\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24530\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__24530\,
            I => n164
        );

    \I__5231\ : InMux
    port map (
            O => \N__24527\,
            I => \N__24524\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__24524\,
            I => n4_adj_361
        );

    \I__5229\ : CascadeMux
    port map (
            O => \N__24521\,
            I => \n4_adj_361_cascade_\
        );

    \I__5228\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24515\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__24515\,
            I => n162
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__24512\,
            I => \n5361_cascade_\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__24509\,
            I => \N__24505\
        );

    \I__5224\ : InMux
    port map (
            O => \N__24508\,
            I => \N__24502\
        );

    \I__5223\ : InMux
    port map (
            O => \N__24505\,
            I => \N__24499\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__24502\,
            I => \N__24494\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__24499\,
            I => \N__24494\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__24494\,
            I => \N__24490\
        );

    \I__5219\ : InMux
    port map (
            O => \N__24493\,
            I => \N__24487\
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__24490\,
            I => \eeprom.n2508\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__24487\,
            I => \eeprom.n2508\
        );

    \I__5216\ : CascadeMux
    port map (
            O => \N__24482\,
            I => \N__24479\
        );

    \I__5215\ : InMux
    port map (
            O => \N__24479\,
            I => \N__24476\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__24476\,
            I => \eeprom.n2575\
        );

    \I__5213\ : InMux
    port map (
            O => \N__24473\,
            I => \eeprom.n4040\
        );

    \I__5212\ : InMux
    port map (
            O => \N__24470\,
            I => \N__24466\
        );

    \I__5211\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24463\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24457\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__24463\,
            I => \N__24457\
        );

    \I__5208\ : InMux
    port map (
            O => \N__24462\,
            I => \N__24454\
        );

    \I__5207\ : Odrv4
    port map (
            O => \N__24457\,
            I => \eeprom.n2507\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__24454\,
            I => \eeprom.n2507\
        );

    \I__5205\ : CascadeMux
    port map (
            O => \N__24449\,
            I => \N__24446\
        );

    \I__5204\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24443\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__24443\,
            I => \eeprom.n2574\
        );

    \I__5202\ : InMux
    port map (
            O => \N__24440\,
            I => \eeprom.n4041\
        );

    \I__5201\ : CascadeMux
    port map (
            O => \N__24437\,
            I => \N__24428\
        );

    \I__5200\ : CascadeMux
    port map (
            O => \N__24436\,
            I => \N__24423\
        );

    \I__5199\ : CascadeMux
    port map (
            O => \N__24435\,
            I => \N__24419\
        );

    \I__5198\ : InMux
    port map (
            O => \N__24434\,
            I => \N__24412\
        );

    \I__5197\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24412\
        );

    \I__5196\ : CascadeMux
    port map (
            O => \N__24432\,
            I => \N__24409\
        );

    \I__5195\ : InMux
    port map (
            O => \N__24431\,
            I => \N__24401\
        );

    \I__5194\ : InMux
    port map (
            O => \N__24428\,
            I => \N__24401\
        );

    \I__5193\ : InMux
    port map (
            O => \N__24427\,
            I => \N__24401\
        );

    \I__5192\ : InMux
    port map (
            O => \N__24426\,
            I => \N__24398\
        );

    \I__5191\ : InMux
    port map (
            O => \N__24423\,
            I => \N__24393\
        );

    \I__5190\ : InMux
    port map (
            O => \N__24422\,
            I => \N__24393\
        );

    \I__5189\ : InMux
    port map (
            O => \N__24419\,
            I => \N__24386\
        );

    \I__5188\ : InMux
    port map (
            O => \N__24418\,
            I => \N__24386\
        );

    \I__5187\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24386\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__24412\,
            I => \N__24383\
        );

    \I__5185\ : InMux
    port map (
            O => \N__24409\,
            I => \N__24378\
        );

    \I__5184\ : InMux
    port map (
            O => \N__24408\,
            I => \N__24378\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__24401\,
            I => \N__24373\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__24398\,
            I => \N__24373\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__24393\,
            I => \eeprom.n2539\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__24386\,
            I => \eeprom.n2539\
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__24383\,
            I => \eeprom.n2539\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__24378\,
            I => \eeprom.n2539\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__24373\,
            I => \eeprom.n2539\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__24362\,
            I => \N__24359\
        );

    \I__5175\ : InMux
    port map (
            O => \N__24359\,
            I => \N__24356\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__24356\,
            I => \N__24352\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__24355\,
            I => \N__24349\
        );

    \I__5172\ : Span4Mux_v
    port map (
            O => \N__24352\,
            I => \N__24346\
        );

    \I__5171\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24343\
        );

    \I__5170\ : Odrv4
    port map (
            O => \N__24346\,
            I => \eeprom.n2506\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__24343\,
            I => \eeprom.n2506\
        );

    \I__5168\ : InMux
    port map (
            O => \N__24338\,
            I => \eeprom.n4042\
        );

    \I__5167\ : InMux
    port map (
            O => \N__24335\,
            I => \N__24332\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__24332\,
            I => \N__24328\
        );

    \I__5165\ : InMux
    port map (
            O => \N__24331\,
            I => \N__24325\
        );

    \I__5164\ : Odrv4
    port map (
            O => \N__24328\,
            I => \eeprom.n2605\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__24325\,
            I => \eeprom.n2605\
        );

    \I__5162\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24316\
        );

    \I__5161\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24313\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__24316\,
            I => \N__24309\
        );

    \I__5159\ : LocalMux
    port map (
            O => \N__24313\,
            I => \N__24306\
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__24312\,
            I => \N__24303\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__24309\,
            I => \N__24300\
        );

    \I__5156\ : Span4Mux_h
    port map (
            O => \N__24306\,
            I => \N__24297\
        );

    \I__5155\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24294\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__24300\,
            I => \eeprom.n2519\
        );

    \I__5153\ : Odrv4
    port map (
            O => \N__24297\,
            I => \eeprom.n2519\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__24294\,
            I => \eeprom.n2519\
        );

    \I__5151\ : InMux
    port map (
            O => \N__24287\,
            I => \N__24283\
        );

    \I__5150\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24279\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__24283\,
            I => \N__24276\
        );

    \I__5148\ : InMux
    port map (
            O => \N__24282\,
            I => \N__24273\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__24279\,
            I => \N__24270\
        );

    \I__5146\ : Span4Mux_v
    port map (
            O => \N__24276\,
            I => \N__24267\
        );

    \I__5145\ : LocalMux
    port map (
            O => \N__24273\,
            I => \N__24262\
        );

    \I__5144\ : Span4Mux_v
    port map (
            O => \N__24270\,
            I => \N__24262\
        );

    \I__5143\ : Odrv4
    port map (
            O => \N__24267\,
            I => \eeprom.n2619\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__24262\,
            I => \eeprom.n2619\
        );

    \I__5141\ : InMux
    port map (
            O => \N__24257\,
            I => \N__24250\
        );

    \I__5140\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24250\
        );

    \I__5139\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24247\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__24250\,
            I => \N__24242\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__24247\,
            I => \N__24242\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__24242\,
            I => \N__24239\
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__24239\,
            I => \eeprom.n2819\
        );

    \I__5134\ : InMux
    port map (
            O => \N__24236\,
            I => \N__24232\
        );

    \I__5133\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24228\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24225\
        );

    \I__5131\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24222\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__24228\,
            I => \N__24219\
        );

    \I__5129\ : Span4Mux_v
    port map (
            O => \N__24225\,
            I => \N__24214\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__24222\,
            I => \N__24214\
        );

    \I__5127\ : Span4Mux_h
    port map (
            O => \N__24219\,
            I => \N__24211\
        );

    \I__5126\ : Span4Mux_h
    port map (
            O => \N__24214\,
            I => \N__24208\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__24211\,
            I => \N__24205\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__24208\,
            I => \N__24202\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__24205\,
            I => \eeprom.n3219\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__24202\,
            I => \eeprom.n3219\
        );

    \I__5121\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24193\
        );

    \I__5120\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24190\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__24193\,
            I => \N__24184\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24184\
        );

    \I__5117\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24181\
        );

    \I__5116\ : Span4Mux_h
    port map (
            O => \N__24184\,
            I => \N__24178\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__24181\,
            I => \N__24175\
        );

    \I__5114\ : Span4Mux_h
    port map (
            O => \N__24178\,
            I => \N__24172\
        );

    \I__5113\ : Odrv12
    port map (
            O => \N__24175\,
            I => \eeprom.n3019\
        );

    \I__5112\ : Odrv4
    port map (
            O => \N__24172\,
            I => \eeprom.n3019\
        );

    \I__5111\ : CascadeMux
    port map (
            O => \N__24167\,
            I => \N__24164\
        );

    \I__5110\ : InMux
    port map (
            O => \N__24164\,
            I => \N__24159\
        );

    \I__5109\ : InMux
    port map (
            O => \N__24163\,
            I => \N__24156\
        );

    \I__5108\ : InMux
    port map (
            O => \N__24162\,
            I => \N__24153\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__24159\,
            I => \N__24150\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__24156\,
            I => \eeprom.n2516\
        );

    \I__5105\ : LocalMux
    port map (
            O => \N__24153\,
            I => \eeprom.n2516\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__24150\,
            I => \eeprom.n2516\
        );

    \I__5103\ : InMux
    port map (
            O => \N__24143\,
            I => \N__24140\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__24140\,
            I => \eeprom.n2583\
        );

    \I__5101\ : InMux
    port map (
            O => \N__24137\,
            I => \eeprom.n4032\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__24134\,
            I => \N__24131\
        );

    \I__5099\ : InMux
    port map (
            O => \N__24131\,
            I => \N__24126\
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__24130\,
            I => \N__24123\
        );

    \I__5097\ : InMux
    port map (
            O => \N__24129\,
            I => \N__24120\
        );

    \I__5096\ : LocalMux
    port map (
            O => \N__24126\,
            I => \N__24117\
        );

    \I__5095\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24114\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__24120\,
            I => \eeprom.n2515\
        );

    \I__5093\ : Odrv4
    port map (
            O => \N__24117\,
            I => \eeprom.n2515\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__24114\,
            I => \eeprom.n2515\
        );

    \I__5091\ : InMux
    port map (
            O => \N__24107\,
            I => \N__24104\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__24104\,
            I => \eeprom.n2582\
        );

    \I__5089\ : InMux
    port map (
            O => \N__24101\,
            I => \eeprom.n4033\
        );

    \I__5088\ : CascadeMux
    port map (
            O => \N__24098\,
            I => \N__24095\
        );

    \I__5087\ : InMux
    port map (
            O => \N__24095\,
            I => \N__24090\
        );

    \I__5086\ : InMux
    port map (
            O => \N__24094\,
            I => \N__24087\
        );

    \I__5085\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24084\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__24090\,
            I => \N__24081\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__24087\,
            I => \eeprom.n2514\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__24084\,
            I => \eeprom.n2514\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__24081\,
            I => \eeprom.n2514\
        );

    \I__5080\ : InMux
    port map (
            O => \N__24074\,
            I => \N__24071\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__24071\,
            I => \eeprom.n2581\
        );

    \I__5078\ : InMux
    port map (
            O => \N__24068\,
            I => \eeprom.n4034\
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__24065\,
            I => \N__24062\
        );

    \I__5076\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24058\
        );

    \I__5075\ : InMux
    port map (
            O => \N__24061\,
            I => \N__24054\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__24058\,
            I => \N__24051\
        );

    \I__5073\ : InMux
    port map (
            O => \N__24057\,
            I => \N__24048\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__24054\,
            I => \N__24043\
        );

    \I__5071\ : Span4Mux_h
    port map (
            O => \N__24051\,
            I => \N__24043\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__24048\,
            I => \N__24040\
        );

    \I__5069\ : Odrv4
    port map (
            O => \N__24043\,
            I => \eeprom.n2513\
        );

    \I__5068\ : Odrv4
    port map (
            O => \N__24040\,
            I => \eeprom.n2513\
        );

    \I__5067\ : InMux
    port map (
            O => \N__24035\,
            I => \N__24032\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__24032\,
            I => \eeprom.n2580\
        );

    \I__5065\ : InMux
    port map (
            O => \N__24029\,
            I => \eeprom.n4035\
        );

    \I__5064\ : CascadeMux
    port map (
            O => \N__24026\,
            I => \N__24023\
        );

    \I__5063\ : InMux
    port map (
            O => \N__24023\,
            I => \N__24020\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__24020\,
            I => \N__24015\
        );

    \I__5061\ : InMux
    port map (
            O => \N__24019\,
            I => \N__24010\
        );

    \I__5060\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24010\
        );

    \I__5059\ : Span4Mux_h
    port map (
            O => \N__24015\,
            I => \N__24007\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__24010\,
            I => \eeprom.n2512\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__24007\,
            I => \eeprom.n2512\
        );

    \I__5056\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23999\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__23999\,
            I => \eeprom.n2579\
        );

    \I__5054\ : InMux
    port map (
            O => \N__23996\,
            I => \eeprom.n4036\
        );

    \I__5053\ : CascadeMux
    port map (
            O => \N__23993\,
            I => \N__23990\
        );

    \I__5052\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23986\
        );

    \I__5051\ : InMux
    port map (
            O => \N__23989\,
            I => \N__23983\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__23986\,
            I => \N__23980\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__23983\,
            I => \N__23977\
        );

    \I__5048\ : Span4Mux_h
    port map (
            O => \N__23980\,
            I => \N__23974\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__23977\,
            I => \eeprom.n2511\
        );

    \I__5046\ : Odrv4
    port map (
            O => \N__23974\,
            I => \eeprom.n2511\
        );

    \I__5045\ : InMux
    port map (
            O => \N__23969\,
            I => \N__23966\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__23966\,
            I => \N__23963\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__23963\,
            I => \N__23960\
        );

    \I__5042\ : Odrv4
    port map (
            O => \N__23960\,
            I => \eeprom.n2578\
        );

    \I__5041\ : InMux
    port map (
            O => \N__23957\,
            I => \bfn_24_24_0_\
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__23954\,
            I => \N__23951\
        );

    \I__5039\ : InMux
    port map (
            O => \N__23951\,
            I => \N__23948\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__23948\,
            I => \N__23944\
        );

    \I__5037\ : InMux
    port map (
            O => \N__23947\,
            I => \N__23941\
        );

    \I__5036\ : Sp12to4
    port map (
            O => \N__23944\,
            I => \N__23935\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__23941\,
            I => \N__23935\
        );

    \I__5034\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23932\
        );

    \I__5033\ : Odrv12
    port map (
            O => \N__23935\,
            I => \eeprom.n2510\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__23932\,
            I => \eeprom.n2510\
        );

    \I__5031\ : InMux
    port map (
            O => \N__23927\,
            I => \N__23924\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__23924\,
            I => \eeprom.n2577\
        );

    \I__5029\ : InMux
    port map (
            O => \N__23921\,
            I => \eeprom.n4038\
        );

    \I__5028\ : CascadeMux
    port map (
            O => \N__23918\,
            I => \N__23914\
        );

    \I__5027\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23911\
        );

    \I__5026\ : InMux
    port map (
            O => \N__23914\,
            I => \N__23908\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__23911\,
            I => \N__23902\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__23908\,
            I => \N__23902\
        );

    \I__5023\ : InMux
    port map (
            O => \N__23907\,
            I => \N__23899\
        );

    \I__5022\ : Odrv4
    port map (
            O => \N__23902\,
            I => \eeprom.n2509\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__23899\,
            I => \eeprom.n2509\
        );

    \I__5020\ : InMux
    port map (
            O => \N__23894\,
            I => \N__23891\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__23891\,
            I => \eeprom.n2576\
        );

    \I__5018\ : InMux
    port map (
            O => \N__23888\,
            I => \eeprom.n4039\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__23885\,
            I => \eeprom.n5173_cascade_\
        );

    \I__5016\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23879\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__23879\,
            I => \eeprom.n11_adj_328\
        );

    \I__5014\ : CascadeMux
    port map (
            O => \N__23876\,
            I => \N__23872\
        );

    \I__5013\ : CascadeMux
    port map (
            O => \N__23875\,
            I => \N__23869\
        );

    \I__5012\ : InMux
    port map (
            O => \N__23872\,
            I => \N__23866\
        );

    \I__5011\ : InMux
    port map (
            O => \N__23869\,
            I => \N__23863\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__23866\,
            I => \N__23860\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__23863\,
            I => \N__23857\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__23860\,
            I => \N__23854\
        );

    \I__5007\ : Odrv4
    port map (
            O => \N__23857\,
            I => \eeprom.n2615\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__23854\,
            I => \eeprom.n2615\
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__23849\,
            I => \eeprom.n2615_cascade_\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__23846\,
            I => \N__23843\
        );

    \I__5003\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23839\
        );

    \I__5002\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23836\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__23839\,
            I => \N__23833\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__23836\,
            I => \N__23829\
        );

    \I__4999\ : Span4Mux_v
    port map (
            O => \N__23833\,
            I => \N__23826\
        );

    \I__4998\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23823\
        );

    \I__4997\ : Odrv4
    port map (
            O => \N__23829\,
            I => \eeprom.n2613\
        );

    \I__4996\ : Odrv4
    port map (
            O => \N__23826\,
            I => \eeprom.n2613\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__23823\,
            I => \eeprom.n2613\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__23816\,
            I => \N__23813\
        );

    \I__4993\ : InMux
    port map (
            O => \N__23813\,
            I => \N__23810\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23806\
        );

    \I__4991\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23802\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__23806\,
            I => \N__23799\
        );

    \I__4989\ : InMux
    port map (
            O => \N__23805\,
            I => \N__23796\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__23802\,
            I => \eeprom.n2617\
        );

    \I__4987\ : Odrv4
    port map (
            O => \N__23799\,
            I => \eeprom.n2617\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__23796\,
            I => \eeprom.n2617\
        );

    \I__4985\ : CascadeMux
    port map (
            O => \N__23789\,
            I => \N__23786\
        );

    \I__4984\ : InMux
    port map (
            O => \N__23786\,
            I => \N__23783\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23779\
        );

    \I__4982\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23775\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__23779\,
            I => \N__23772\
        );

    \I__4980\ : InMux
    port map (
            O => \N__23778\,
            I => \N__23769\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__23775\,
            I => \eeprom.n2614\
        );

    \I__4978\ : Odrv4
    port map (
            O => \N__23772\,
            I => \eeprom.n2614\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__23769\,
            I => \eeprom.n2614\
        );

    \I__4976\ : CascadeMux
    port map (
            O => \N__23762\,
            I => \eeprom.n5101_cascade_\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__23759\,
            I => \N__23756\
        );

    \I__4974\ : InMux
    port map (
            O => \N__23756\,
            I => \N__23753\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__23753\,
            I => \N__23749\
        );

    \I__4972\ : InMux
    port map (
            O => \N__23752\,
            I => \N__23745\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__23749\,
            I => \N__23742\
        );

    \I__4970\ : InMux
    port map (
            O => \N__23748\,
            I => \N__23739\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__23745\,
            I => \eeprom.n2616\
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__23742\,
            I => \eeprom.n2616\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__23739\,
            I => \eeprom.n2616\
        );

    \I__4966\ : CascadeMux
    port map (
            O => \N__23732\,
            I => \N__23729\
        );

    \I__4965\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23726\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__23726\,
            I => \eeprom.n5105\
        );

    \I__4963\ : InMux
    port map (
            O => \N__23723\,
            I => \N__23720\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__23720\,
            I => \N__23717\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__23717\,
            I => \N__23714\
        );

    \I__4960\ : Odrv4
    port map (
            O => \N__23714\,
            I => \eeprom.n2586\
        );

    \I__4959\ : InMux
    port map (
            O => \N__23711\,
            I => \bfn_24_23_0_\
        );

    \I__4958\ : CascadeMux
    port map (
            O => \N__23708\,
            I => \N__23704\
        );

    \I__4957\ : CascadeMux
    port map (
            O => \N__23707\,
            I => \N__23701\
        );

    \I__4956\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23697\
        );

    \I__4955\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23694\
        );

    \I__4954\ : InMux
    port map (
            O => \N__23700\,
            I => \N__23691\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__23697\,
            I => \N__23688\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__23694\,
            I => \eeprom.n2518\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__23691\,
            I => \eeprom.n2518\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__23688\,
            I => \eeprom.n2518\
        );

    \I__4949\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23678\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__23678\,
            I => \eeprom.n2585\
        );

    \I__4947\ : InMux
    port map (
            O => \N__23675\,
            I => \eeprom.n4030\
        );

    \I__4946\ : CascadeMux
    port map (
            O => \N__23672\,
            I => \N__23668\
        );

    \I__4945\ : CascadeMux
    port map (
            O => \N__23671\,
            I => \N__23665\
        );

    \I__4944\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23661\
        );

    \I__4943\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23658\
        );

    \I__4942\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23655\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__23661\,
            I => \N__23652\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__23658\,
            I => \eeprom.n2517\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__23655\,
            I => \eeprom.n2517\
        );

    \I__4938\ : Odrv4
    port map (
            O => \N__23652\,
            I => \eeprom.n2517\
        );

    \I__4937\ : InMux
    port map (
            O => \N__23645\,
            I => \N__23642\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__23642\,
            I => \eeprom.n2584\
        );

    \I__4935\ : InMux
    port map (
            O => \N__23639\,
            I => \eeprom.n4031\
        );

    \I__4934\ : InMux
    port map (
            O => \N__23636\,
            I => \N__23633\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__23633\,
            I => \eeprom.n1982\
        );

    \I__4932\ : InMux
    port map (
            O => \N__23630\,
            I => \eeprom.n3976\
        );

    \I__4931\ : InMux
    port map (
            O => \N__23627\,
            I => \N__23624\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__23624\,
            I => \eeprom.n1981\
        );

    \I__4929\ : InMux
    port map (
            O => \N__23621\,
            I => \eeprom.n3977\
        );

    \I__4928\ : CascadeMux
    port map (
            O => \N__23618\,
            I => \N__23615\
        );

    \I__4927\ : InMux
    port map (
            O => \N__23615\,
            I => \N__23612\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__23612\,
            I => \eeprom.n1980\
        );

    \I__4925\ : InMux
    port map (
            O => \N__23609\,
            I => \eeprom.n3978\
        );

    \I__4924\ : CascadeMux
    port map (
            O => \N__23606\,
            I => \N__23600\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__23605\,
            I => \N__23597\
        );

    \I__4922\ : CascadeMux
    port map (
            O => \N__23604\,
            I => \N__23593\
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__23603\,
            I => \N__23589\
        );

    \I__4920\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23585\
        );

    \I__4919\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23580\
        );

    \I__4918\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23580\
        );

    \I__4917\ : InMux
    port map (
            O => \N__23593\,
            I => \N__23571\
        );

    \I__4916\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23571\
        );

    \I__4915\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23571\
        );

    \I__4914\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23571\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__23585\,
            I => \eeprom.n1945\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__23580\,
            I => \eeprom.n1945\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__23571\,
            I => \eeprom.n1945\
        );

    \I__4910\ : InMux
    port map (
            O => \N__23564\,
            I => \eeprom.n3979\
        );

    \I__4909\ : InMux
    port map (
            O => \N__23561\,
            I => \N__23557\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__23560\,
            I => \N__23554\
        );

    \I__4907\ : LocalMux
    port map (
            O => \N__23557\,
            I => \N__23551\
        );

    \I__4906\ : InMux
    port map (
            O => \N__23554\,
            I => \N__23548\
        );

    \I__4905\ : Span4Mux_h
    port map (
            O => \N__23551\,
            I => \N__23545\
        );

    \I__4904\ : LocalMux
    port map (
            O => \N__23548\,
            I => \eeprom.n2011\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__23545\,
            I => \eeprom.n2011\
        );

    \I__4902\ : InMux
    port map (
            O => \N__23540\,
            I => \N__23536\
        );

    \I__4901\ : CascadeMux
    port map (
            O => \N__23539\,
            I => \N__23533\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__23536\,
            I => \N__23530\
        );

    \I__4899\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23527\
        );

    \I__4898\ : Span4Mux_h
    port map (
            O => \N__23530\,
            I => \N__23523\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__23527\,
            I => \N__23520\
        );

    \I__4896\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23517\
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__23523\,
            I => \eeprom.n2411\
        );

    \I__4894\ : Odrv4
    port map (
            O => \N__23520\,
            I => \eeprom.n2411\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__23517\,
            I => \eeprom.n2411\
        );

    \I__4892\ : CascadeMux
    port map (
            O => \N__23510\,
            I => \N__23507\
        );

    \I__4891\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23504\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__23504\,
            I => \N__23501\
        );

    \I__4889\ : Span4Mux_h
    port map (
            O => \N__23501\,
            I => \N__23498\
        );

    \I__4888\ : Odrv4
    port map (
            O => \N__23498\,
            I => \eeprom.n2478\
        );

    \I__4887\ : InMux
    port map (
            O => \N__23495\,
            I => \N__23487\
        );

    \I__4886\ : InMux
    port map (
            O => \N__23494\,
            I => \N__23483\
        );

    \I__4885\ : CascadeMux
    port map (
            O => \N__23493\,
            I => \N__23480\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__23492\,
            I => \N__23476\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__23491\,
            I => \N__23471\
        );

    \I__4882\ : CascadeMux
    port map (
            O => \N__23490\,
            I => \N__23468\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__23487\,
            I => \N__23463\
        );

    \I__4880\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23460\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__23483\,
            I => \N__23457\
        );

    \I__4878\ : InMux
    port map (
            O => \N__23480\,
            I => \N__23452\
        );

    \I__4877\ : InMux
    port map (
            O => \N__23479\,
            I => \N__23452\
        );

    \I__4876\ : InMux
    port map (
            O => \N__23476\,
            I => \N__23437\
        );

    \I__4875\ : InMux
    port map (
            O => \N__23475\,
            I => \N__23437\
        );

    \I__4874\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23437\
        );

    \I__4873\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23437\
        );

    \I__4872\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23437\
        );

    \I__4871\ : InMux
    port map (
            O => \N__23467\,
            I => \N__23437\
        );

    \I__4870\ : InMux
    port map (
            O => \N__23466\,
            I => \N__23437\
        );

    \I__4869\ : Odrv4
    port map (
            O => \N__23463\,
            I => \eeprom.n2440\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__23460\,
            I => \eeprom.n2440\
        );

    \I__4867\ : Odrv4
    port map (
            O => \N__23457\,
            I => \eeprom.n2440\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__23452\,
            I => \eeprom.n2440\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__23437\,
            I => \eeprom.n2440\
        );

    \I__4864\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23423\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__23423\,
            I => \N__23418\
        );

    \I__4862\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23415\
        );

    \I__4861\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23412\
        );

    \I__4860\ : Span4Mux_v
    port map (
            O => \N__23418\,
            I => \N__23407\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__23415\,
            I => \N__23407\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23404\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__23407\,
            I => \N__23401\
        );

    \I__4856\ : Odrv12
    port map (
            O => \N__23404\,
            I => \eeprom.n3419\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__23401\,
            I => \eeprom.n3419\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__23396\,
            I => \eeprom.n5169_cascade_\
        );

    \I__4853\ : CascadeMux
    port map (
            O => \N__23393\,
            I => \N__23389\
        );

    \I__4852\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23386\
        );

    \I__4851\ : InMux
    port map (
            O => \N__23389\,
            I => \N__23383\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__23386\,
            I => \N__23380\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__23383\,
            I => \eeprom.n2016\
        );

    \I__4848\ : Odrv4
    port map (
            O => \N__23380\,
            I => \eeprom.n2016\
        );

    \I__4847\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23372\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__23372\,
            I => \eeprom.n2083\
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__23369\,
            I => \eeprom.n2016_cascade_\
        );

    \I__4844\ : CascadeMux
    port map (
            O => \N__23366\,
            I => \N__23360\
        );

    \I__4843\ : InMux
    port map (
            O => \N__23365\,
            I => \N__23354\
        );

    \I__4842\ : InMux
    port map (
            O => \N__23364\,
            I => \N__23345\
        );

    \I__4841\ : InMux
    port map (
            O => \N__23363\,
            I => \N__23345\
        );

    \I__4840\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23345\
        );

    \I__4839\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23345\
        );

    \I__4838\ : CascadeMux
    port map (
            O => \N__23358\,
            I => \N__23342\
        );

    \I__4837\ : InMux
    port map (
            O => \N__23357\,
            I => \N__23337\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23334\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__23345\,
            I => \N__23331\
        );

    \I__4834\ : InMux
    port map (
            O => \N__23342\,
            I => \N__23324\
        );

    \I__4833\ : InMux
    port map (
            O => \N__23341\,
            I => \N__23324\
        );

    \I__4832\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23324\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__23337\,
            I => \eeprom.n2044\
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__23334\,
            I => \eeprom.n2044\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__23331\,
            I => \eeprom.n2044\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__23324\,
            I => \eeprom.n2044\
        );

    \I__4827\ : CascadeMux
    port map (
            O => \N__23315\,
            I => \N__23311\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__23314\,
            I => \N__23308\
        );

    \I__4825\ : InMux
    port map (
            O => \N__23311\,
            I => \N__23305\
        );

    \I__4824\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23302\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__23305\,
            I => \N__23299\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__23302\,
            I => \N__23296\
        );

    \I__4821\ : Odrv4
    port map (
            O => \N__23299\,
            I => \eeprom.n2115\
        );

    \I__4820\ : Odrv4
    port map (
            O => \N__23296\,
            I => \eeprom.n2115\
        );

    \I__4819\ : CascadeMux
    port map (
            O => \N__23291\,
            I => \eeprom.n2115_cascade_\
        );

    \I__4818\ : CascadeMux
    port map (
            O => \N__23288\,
            I => \N__23285\
        );

    \I__4817\ : InMux
    port map (
            O => \N__23285\,
            I => \N__23281\
        );

    \I__4816\ : InMux
    port map (
            O => \N__23284\,
            I => \N__23277\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__23281\,
            I => \N__23274\
        );

    \I__4814\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23271\
        );

    \I__4813\ : LocalMux
    port map (
            O => \N__23277\,
            I => \eeprom.n2113\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__23274\,
            I => \eeprom.n2113\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__23271\,
            I => \eeprom.n2113\
        );

    \I__4810\ : InMux
    port map (
            O => \N__23264\,
            I => \N__23261\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__23261\,
            I => \eeprom.n5059\
        );

    \I__4808\ : InMux
    port map (
            O => \N__23258\,
            I => \N__23253\
        );

    \I__4807\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23250\
        );

    \I__4806\ : CascadeMux
    port map (
            O => \N__23256\,
            I => \N__23247\
        );

    \I__4805\ : LocalMux
    port map (
            O => \N__23253\,
            I => \N__23242\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23242\
        );

    \I__4803\ : InMux
    port map (
            O => \N__23247\,
            I => \N__23239\
        );

    \I__4802\ : Span4Mux_h
    port map (
            O => \N__23242\,
            I => \N__23236\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__23239\,
            I => \eeprom.n2013\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__23236\,
            I => \eeprom.n2013\
        );

    \I__4799\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23226\
        );

    \I__4798\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23223\
        );

    \I__4797\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23220\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__23226\,
            I => \N__23217\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__23223\,
            I => \eeprom.n2012\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__23220\,
            I => \eeprom.n2012\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__23217\,
            I => \eeprom.n2012\
        );

    \I__4792\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23207\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__23207\,
            I => \N__23204\
        );

    \I__4790\ : Odrv4
    port map (
            O => \N__23204\,
            I => \eeprom.n1986\
        );

    \I__4789\ : InMux
    port map (
            O => \N__23201\,
            I => \bfn_24_20_0_\
        );

    \I__4788\ : InMux
    port map (
            O => \N__23198\,
            I => \N__23195\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__23195\,
            I => \eeprom.n1985\
        );

    \I__4786\ : InMux
    port map (
            O => \N__23192\,
            I => \eeprom.n3973\
        );

    \I__4785\ : InMux
    port map (
            O => \N__23189\,
            I => \N__23186\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__23186\,
            I => \eeprom.n1984\
        );

    \I__4783\ : InMux
    port map (
            O => \N__23183\,
            I => \eeprom.n3974\
        );

    \I__4782\ : InMux
    port map (
            O => \N__23180\,
            I => \N__23177\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__23177\,
            I => \N__23174\
        );

    \I__4780\ : Odrv4
    port map (
            O => \N__23174\,
            I => \eeprom.n1983\
        );

    \I__4779\ : InMux
    port map (
            O => \N__23171\,
            I => \eeprom.n3975\
        );

    \I__4778\ : InMux
    port map (
            O => \N__23168\,
            I => \N__23164\
        );

    \I__4777\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23161\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__23164\,
            I => \eeprom.n2110\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__23161\,
            I => \eeprom.n2110\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__23156\,
            I => \N__23151\
        );

    \I__4773\ : CascadeMux
    port map (
            O => \N__23155\,
            I => \N__23148\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__23154\,
            I => \N__23141\
        );

    \I__4771\ : InMux
    port map (
            O => \N__23151\,
            I => \N__23134\
        );

    \I__4770\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23131\
        );

    \I__4769\ : InMux
    port map (
            O => \N__23147\,
            I => \N__23128\
        );

    \I__4768\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23121\
        );

    \I__4767\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23121\
        );

    \I__4766\ : InMux
    port map (
            O => \N__23144\,
            I => \N__23121\
        );

    \I__4765\ : InMux
    port map (
            O => \N__23141\,
            I => \N__23116\
        );

    \I__4764\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23116\
        );

    \I__4763\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23109\
        );

    \I__4762\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23109\
        );

    \I__4761\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23109\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__23134\,
            I => \N__23106\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__23131\,
            I => \eeprom.n2143\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__23128\,
            I => \eeprom.n2143\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__23121\,
            I => \eeprom.n2143\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__23116\,
            I => \eeprom.n2143\
        );

    \I__4755\ : LocalMux
    port map (
            O => \N__23109\,
            I => \eeprom.n2143\
        );

    \I__4754\ : Odrv4
    port map (
            O => \N__23106\,
            I => \eeprom.n2143\
        );

    \I__4753\ : InMux
    port map (
            O => \N__23093\,
            I => \eeprom.n3996\
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__23090\,
            I => \N__23086\
        );

    \I__4751\ : CascadeMux
    port map (
            O => \N__23089\,
            I => \N__23083\
        );

    \I__4750\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23080\
        );

    \I__4749\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23077\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__23074\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23071\
        );

    \I__4746\ : Odrv12
    port map (
            O => \N__23074\,
            I => \eeprom.n2209\
        );

    \I__4745\ : Odrv4
    port map (
            O => \N__23071\,
            I => \eeprom.n2209\
        );

    \I__4744\ : InMux
    port map (
            O => \N__23066\,
            I => \N__23063\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__23063\,
            I => \N__23060\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__23060\,
            I => \N__23057\
        );

    \I__4741\ : Odrv4
    port map (
            O => \N__23057\,
            I => \eeprom.n3724\
        );

    \I__4740\ : CascadeMux
    port map (
            O => \N__23054\,
            I => \N__23051\
        );

    \I__4739\ : InMux
    port map (
            O => \N__23051\,
            I => \N__23046\
        );

    \I__4738\ : InMux
    port map (
            O => \N__23050\,
            I => \N__23041\
        );

    \I__4737\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23041\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__23046\,
            I => \eeprom.n2015\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__23041\,
            I => \eeprom.n2015\
        );

    \I__4734\ : CascadeMux
    port map (
            O => \N__23036\,
            I => \N__23033\
        );

    \I__4733\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23030\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__23030\,
            I => \eeprom.n2079\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__23027\,
            I => \N__23022\
        );

    \I__4730\ : InMux
    port map (
            O => \N__23026\,
            I => \N__23019\
        );

    \I__4729\ : InMux
    port map (
            O => \N__23025\,
            I => \N__23016\
        );

    \I__4728\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23013\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__23019\,
            I => \N__23010\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__23016\,
            I => \eeprom.n2111\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__23013\,
            I => \eeprom.n2111\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__23010\,
            I => \eeprom.n2111\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__23003\,
            I => \N__22999\
        );

    \I__4722\ : CascadeMux
    port map (
            O => \N__23002\,
            I => \N__22995\
        );

    \I__4721\ : InMux
    port map (
            O => \N__22999\,
            I => \N__22990\
        );

    \I__4720\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22990\
        );

    \I__4719\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22987\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__22990\,
            I => \eeprom.n2018\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__22987\,
            I => \eeprom.n2018\
        );

    \I__4716\ : CascadeMux
    port map (
            O => \N__22982\,
            I => \eeprom.n1945_cascade_\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__22979\,
            I => \N__22973\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__22978\,
            I => \N__22970\
        );

    \I__4713\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22967\
        );

    \I__4712\ : CascadeMux
    port map (
            O => \N__22976\,
            I => \N__22964\
        );

    \I__4711\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22959\
        );

    \I__4710\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22959\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__22967\,
            I => \N__22956\
        );

    \I__4708\ : InMux
    port map (
            O => \N__22964\,
            I => \N__22953\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__22959\,
            I => \N__22950\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__22956\,
            I => \eeprom.n2017\
        );

    \I__4705\ : LocalMux
    port map (
            O => \N__22953\,
            I => \eeprom.n2017\
        );

    \I__4704\ : Odrv4
    port map (
            O => \N__22950\,
            I => \eeprom.n2017\
        );

    \I__4703\ : CascadeMux
    port map (
            O => \N__22943\,
            I => \N__22938\
        );

    \I__4702\ : CascadeMux
    port map (
            O => \N__22942\,
            I => \N__22935\
        );

    \I__4701\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22932\
        );

    \I__4700\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22929\
        );

    \I__4699\ : InMux
    port map (
            O => \N__22935\,
            I => \N__22926\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__22932\,
            I => \N__22923\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__22929\,
            I => \eeprom.n2014\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__22926\,
            I => \eeprom.n2014\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__22923\,
            I => \eeprom.n2014\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__22916\,
            I => \N__22913\
        );

    \I__4693\ : InMux
    port map (
            O => \N__22913\,
            I => \N__22909\
        );

    \I__4692\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22906\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22903\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__22906\,
            I => \eeprom.n2118\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__22903\,
            I => \eeprom.n2118\
        );

    \I__4688\ : InMux
    port map (
            O => \N__22898\,
            I => \N__22895\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__22895\,
            I => \N__22892\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__22892\,
            I => \N__22889\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__22889\,
            I => \eeprom.n2185\
        );

    \I__4684\ : InMux
    port map (
            O => \N__22886\,
            I => \eeprom.n3988\
        );

    \I__4683\ : CascadeMux
    port map (
            O => \N__22883\,
            I => \N__22879\
        );

    \I__4682\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22875\
        );

    \I__4681\ : InMux
    port map (
            O => \N__22879\,
            I => \N__22872\
        );

    \I__4680\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22869\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__22875\,
            I => \eeprom.n2117\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__22872\,
            I => \eeprom.n2117\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__22869\,
            I => \eeprom.n2117\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__22862\,
            I => \N__22859\
        );

    \I__4675\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22856\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__22856\,
            I => \N__22853\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__22853\,
            I => \N__22850\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__22850\,
            I => \eeprom.n2184\
        );

    \I__4671\ : InMux
    port map (
            O => \N__22847\,
            I => \eeprom.n3989\
        );

    \I__4670\ : CascadeMux
    port map (
            O => \N__22844\,
            I => \N__22841\
        );

    \I__4669\ : InMux
    port map (
            O => \N__22841\,
            I => \N__22838\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__22838\,
            I => \N__22834\
        );

    \I__4667\ : CascadeMux
    port map (
            O => \N__22837\,
            I => \N__22831\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__22834\,
            I => \N__22828\
        );

    \I__4665\ : InMux
    port map (
            O => \N__22831\,
            I => \N__22825\
        );

    \I__4664\ : Odrv4
    port map (
            O => \N__22828\,
            I => \eeprom.n2116\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__22825\,
            I => \eeprom.n2116\
        );

    \I__4662\ : InMux
    port map (
            O => \N__22820\,
            I => \N__22816\
        );

    \I__4661\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22813\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__22816\,
            I => \N__22810\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__22813\,
            I => \N__22807\
        );

    \I__4658\ : Span4Mux_v
    port map (
            O => \N__22810\,
            I => \N__22804\
        );

    \I__4657\ : Span4Mux_h
    port map (
            O => \N__22807\,
            I => \N__22801\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__22804\,
            I => \eeprom.n2183\
        );

    \I__4655\ : Odrv4
    port map (
            O => \N__22801\,
            I => \eeprom.n2183\
        );

    \I__4654\ : InMux
    port map (
            O => \N__22796\,
            I => \eeprom.n3990\
        );

    \I__4653\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22790\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__22790\,
            I => \N__22787\
        );

    \I__4651\ : Span4Mux_h
    port map (
            O => \N__22787\,
            I => \N__22784\
        );

    \I__4650\ : Odrv4
    port map (
            O => \N__22784\,
            I => \eeprom.n2182\
        );

    \I__4649\ : InMux
    port map (
            O => \N__22781\,
            I => \eeprom.n3991\
        );

    \I__4648\ : CascadeMux
    port map (
            O => \N__22778\,
            I => \N__22774\
        );

    \I__4647\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22770\
        );

    \I__4646\ : InMux
    port map (
            O => \N__22774\,
            I => \N__22767\
        );

    \I__4645\ : InMux
    port map (
            O => \N__22773\,
            I => \N__22764\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__22770\,
            I => \eeprom.n2114\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__22767\,
            I => \eeprom.n2114\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__22764\,
            I => \eeprom.n2114\
        );

    \I__4641\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22754\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__22754\,
            I => \N__22751\
        );

    \I__4639\ : Span4Mux_v
    port map (
            O => \N__22751\,
            I => \N__22748\
        );

    \I__4638\ : Odrv4
    port map (
            O => \N__22748\,
            I => \eeprom.n2181\
        );

    \I__4637\ : InMux
    port map (
            O => \N__22745\,
            I => \eeprom.n3992\
        );

    \I__4636\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22739\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__22739\,
            I => \N__22736\
        );

    \I__4634\ : Odrv4
    port map (
            O => \N__22736\,
            I => \eeprom.n2180\
        );

    \I__4633\ : InMux
    port map (
            O => \N__22733\,
            I => \eeprom.n3993\
        );

    \I__4632\ : InMux
    port map (
            O => \N__22730\,
            I => \N__22727\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__22727\,
            I => \N__22722\
        );

    \I__4630\ : CascadeMux
    port map (
            O => \N__22726\,
            I => \N__22719\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__22725\,
            I => \N__22716\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__22722\,
            I => \N__22713\
        );

    \I__4627\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22710\
        );

    \I__4626\ : InMux
    port map (
            O => \N__22716\,
            I => \N__22707\
        );

    \I__4625\ : Odrv4
    port map (
            O => \N__22713\,
            I => \eeprom.n2112\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__22710\,
            I => \eeprom.n2112\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__22707\,
            I => \eeprom.n2112\
        );

    \I__4622\ : CascadeMux
    port map (
            O => \N__22700\,
            I => \N__22697\
        );

    \I__4621\ : InMux
    port map (
            O => \N__22697\,
            I => \N__22694\
        );

    \I__4620\ : LocalMux
    port map (
            O => \N__22694\,
            I => \N__22691\
        );

    \I__4619\ : Span4Mux_h
    port map (
            O => \N__22691\,
            I => \N__22688\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__22688\,
            I => \eeprom.n2179\
        );

    \I__4617\ : InMux
    port map (
            O => \N__22685\,
            I => \eeprom.n3994\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__22682\,
            I => \N__22679\
        );

    \I__4615\ : InMux
    port map (
            O => \N__22679\,
            I => \N__22676\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__22676\,
            I => \eeprom.n2178\
        );

    \I__4613\ : InMux
    port map (
            O => \N__22673\,
            I => \bfn_24_18_0_\
        );

    \I__4612\ : InMux
    port map (
            O => \N__22670\,
            I => \N__22667\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__22667\,
            I => \N__22663\
        );

    \I__4610\ : InMux
    port map (
            O => \N__22666\,
            I => \N__22660\
        );

    \I__4609\ : Span4Mux_v
    port map (
            O => \N__22663\,
            I => \N__22654\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__22660\,
            I => \N__22654\
        );

    \I__4607\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22651\
        );

    \I__4606\ : Sp12to4
    port map (
            O => \N__22654\,
            I => \N__22646\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__22651\,
            I => \N__22646\
        );

    \I__4604\ : Odrv12
    port map (
            O => \N__22646\,
            I => \eeprom.n3319\
        );

    \I__4603\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22639\
        );

    \I__4602\ : InMux
    port map (
            O => \N__22642\,
            I => \N__22635\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__22639\,
            I => \N__22632\
        );

    \I__4600\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22629\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__22635\,
            I => \eeprom.n2608\
        );

    \I__4598\ : Odrv4
    port map (
            O => \N__22632\,
            I => \eeprom.n2608\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__22629\,
            I => \eeprom.n2608\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__22622\,
            I => \N__22619\
        );

    \I__4595\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22616\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__22616\,
            I => \N__22612\
        );

    \I__4593\ : InMux
    port map (
            O => \N__22615\,
            I => \N__22609\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__22612\,
            I => \eeprom.n2607\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__22609\,
            I => \eeprom.n2607\
        );

    \I__4590\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22598\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__22598\,
            I => \eeprom.n2674\
        );

    \I__4587\ : CascadeMux
    port map (
            O => \N__22595\,
            I => \eeprom.n2607_cascade_\
        );

    \I__4586\ : CascadeMux
    port map (
            O => \N__22592\,
            I => \N__22584\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__22591\,
            I => \N__22581\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__22590\,
            I => \N__22577\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__22589\,
            I => \N__22572\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__22588\,
            I => \N__22569\
        );

    \I__4581\ : CascadeMux
    port map (
            O => \N__22587\,
            I => \N__22565\
        );

    \I__4580\ : InMux
    port map (
            O => \N__22584\,
            I => \N__22556\
        );

    \I__4579\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22556\
        );

    \I__4578\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22551\
        );

    \I__4577\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22551\
        );

    \I__4576\ : InMux
    port map (
            O => \N__22576\,
            I => \N__22540\
        );

    \I__4575\ : InMux
    port map (
            O => \N__22575\,
            I => \N__22540\
        );

    \I__4574\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22540\
        );

    \I__4573\ : InMux
    port map (
            O => \N__22569\,
            I => \N__22540\
        );

    \I__4572\ : InMux
    port map (
            O => \N__22568\,
            I => \N__22540\
        );

    \I__4571\ : InMux
    port map (
            O => \N__22565\,
            I => \N__22535\
        );

    \I__4570\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22535\
        );

    \I__4569\ : InMux
    port map (
            O => \N__22563\,
            I => \N__22532\
        );

    \I__4568\ : InMux
    port map (
            O => \N__22562\,
            I => \N__22527\
        );

    \I__4567\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22527\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__22556\,
            I => \N__22524\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__22551\,
            I => \eeprom.n2638\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__22540\,
            I => \eeprom.n2638\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__22535\,
            I => \eeprom.n2638\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__22532\,
            I => \eeprom.n2638\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__22527\,
            I => \eeprom.n2638\
        );

    \I__4560\ : Odrv4
    port map (
            O => \N__22524\,
            I => \eeprom.n2638\
        );

    \I__4559\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22507\
        );

    \I__4558\ : InMux
    port map (
            O => \N__22510\,
            I => \N__22504\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__22507\,
            I => \N__22501\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__22504\,
            I => \N__22495\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__22501\,
            I => \N__22495\
        );

    \I__4554\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22492\
        );

    \I__4553\ : Odrv4
    port map (
            O => \N__22495\,
            I => \eeprom.n2706\
        );

    \I__4552\ : LocalMux
    port map (
            O => \N__22492\,
            I => \eeprom.n2706\
        );

    \I__4551\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22482\
        );

    \I__4550\ : InMux
    port map (
            O => \N__22486\,
            I => \N__22479\
        );

    \I__4549\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22476\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__22482\,
            I => \N__22471\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__22479\,
            I => \N__22471\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__22476\,
            I => \eeprom.n2719\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__22471\,
            I => \eeprom.n2719\
        );

    \I__4544\ : InMux
    port map (
            O => \N__22466\,
            I => \N__22461\
        );

    \I__4543\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22458\
        );

    \I__4542\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22455\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__22461\,
            I => \N__22448\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22448\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__22455\,
            I => \N__22448\
        );

    \I__4538\ : Span4Mux_v
    port map (
            O => \N__22448\,
            I => \N__22445\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__22445\,
            I => \eeprom.n2919\
        );

    \I__4536\ : InMux
    port map (
            O => \N__22442\,
            I => \N__22437\
        );

    \I__4535\ : InMux
    port map (
            O => \N__22441\,
            I => \N__22434\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__22440\,
            I => \N__22431\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22428\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__22434\,
            I => \N__22425\
        );

    \I__4531\ : InMux
    port map (
            O => \N__22431\,
            I => \N__22422\
        );

    \I__4530\ : Span4Mux_h
    port map (
            O => \N__22428\,
            I => \N__22415\
        );

    \I__4529\ : Span4Mux_h
    port map (
            O => \N__22425\,
            I => \N__22415\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__22422\,
            I => \N__22415\
        );

    \I__4527\ : Odrv4
    port map (
            O => \N__22415\,
            I => \eeprom.n2419\
        );

    \I__4526\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22408\
        );

    \I__4525\ : InMux
    port map (
            O => \N__22411\,
            I => \N__22404\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22401\
        );

    \I__4523\ : InMux
    port map (
            O => \N__22407\,
            I => \N__22398\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__22404\,
            I => \N__22395\
        );

    \I__4521\ : Span4Mux_v
    port map (
            O => \N__22401\,
            I => \N__22392\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__22398\,
            I => \N__22389\
        );

    \I__4519\ : Span4Mux_h
    port map (
            O => \N__22395\,
            I => \N__22386\
        );

    \I__4518\ : Span4Mux_h
    port map (
            O => \N__22392\,
            I => \N__22383\
        );

    \I__4517\ : Span4Mux_h
    port map (
            O => \N__22389\,
            I => \N__22378\
        );

    \I__4516\ : Span4Mux_v
    port map (
            O => \N__22386\,
            I => \N__22378\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__22383\,
            I => \eeprom.n3119\
        );

    \I__4514\ : Odrv4
    port map (
            O => \N__22378\,
            I => \eeprom.n3119\
        );

    \I__4513\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22370\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__22370\,
            I => \N__22367\
        );

    \I__4511\ : Span4Mux_h
    port map (
            O => \N__22367\,
            I => \N__22364\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__22364\,
            I => \eeprom.n2186\
        );

    \I__4509\ : InMux
    port map (
            O => \N__22361\,
            I => \bfn_24_17_0_\
        );

    \I__4508\ : InMux
    port map (
            O => \N__22358\,
            I => \N__22354\
        );

    \I__4507\ : InMux
    port map (
            O => \N__22357\,
            I => \N__22351\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__22354\,
            I => \N__22348\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__22351\,
            I => \eeprom.n2612\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__22348\,
            I => \eeprom.n2612\
        );

    \I__4503\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22339\
        );

    \I__4502\ : InMux
    port map (
            O => \N__22342\,
            I => \N__22336\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__22339\,
            I => \N__22333\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__22336\,
            I => \N__22330\
        );

    \I__4499\ : Span4Mux_v
    port map (
            O => \N__22333\,
            I => \N__22326\
        );

    \I__4498\ : Span4Mux_h
    port map (
            O => \N__22330\,
            I => \N__22323\
        );

    \I__4497\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22320\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__22326\,
            I => \eeprom.n2611\
        );

    \I__4495\ : Odrv4
    port map (
            O => \N__22323\,
            I => \eeprom.n2611\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__22320\,
            I => \eeprom.n2611\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__22313\,
            I => \eeprom.n2612_cascade_\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__22310\,
            I => \N__22305\
        );

    \I__4491\ : CascadeMux
    port map (
            O => \N__22309\,
            I => \N__22302\
        );

    \I__4490\ : InMux
    port map (
            O => \N__22308\,
            I => \N__22299\
        );

    \I__4489\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22294\
        );

    \I__4488\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22294\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__22299\,
            I => \N__22291\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__22294\,
            I => \N__22288\
        );

    \I__4485\ : Span4Mux_h
    port map (
            O => \N__22291\,
            I => \N__22285\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__22288\,
            I => \eeprom.n2610\
        );

    \I__4483\ : Odrv4
    port map (
            O => \N__22285\,
            I => \eeprom.n2610\
        );

    \I__4482\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22277\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__22277\,
            I => \eeprom.n16_adj_334\
        );

    \I__4480\ : InMux
    port map (
            O => \N__22274\,
            I => \N__22270\
        );

    \I__4479\ : CascadeMux
    port map (
            O => \N__22273\,
            I => \N__22267\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22264\
        );

    \I__4477\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22261\
        );

    \I__4476\ : Span4Mux_v
    port map (
            O => \N__22264\,
            I => \N__22258\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__22261\,
            I => \eeprom.n2618\
        );

    \I__4474\ : Odrv4
    port map (
            O => \N__22258\,
            I => \eeprom.n2618\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__22253\,
            I => \N__22250\
        );

    \I__4472\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22247\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__22247\,
            I => \eeprom.n12_adj_333\
        );

    \I__4470\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22240\
        );

    \I__4469\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22237\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__22240\,
            I => \N__22234\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22231\
        );

    \I__4466\ : Span4Mux_v
    port map (
            O => \N__22234\,
            I => \N__22228\
        );

    \I__4465\ : Odrv4
    port map (
            O => \N__22231\,
            I => \eeprom.n2606\
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__22228\,
            I => \eeprom.n2606\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__22223\,
            I => \eeprom.n2606_cascade_\
        );

    \I__4462\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22217\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__22217\,
            I => \eeprom.n10_adj_332\
        );

    \I__4460\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22210\
        );

    \I__4459\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22206\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__22210\,
            I => \N__22203\
        );

    \I__4457\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22200\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__22206\,
            I => \N__22195\
        );

    \I__4455\ : Span4Mux_v
    port map (
            O => \N__22203\,
            I => \N__22195\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__22200\,
            I => \eeprom.n2718\
        );

    \I__4453\ : Odrv4
    port map (
            O => \N__22195\,
            I => \eeprom.n2718\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__4451\ : InMux
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__22184\,
            I => \eeprom.n5213\
        );

    \I__4449\ : InMux
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__22178\,
            I => \eeprom.n5215\
        );

    \I__4447\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__22172\,
            I => \eeprom.n4830\
        );

    \I__4445\ : InMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__22166\,
            I => \N__22163\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__22163\,
            I => \N__22160\
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__22160\,
            I => \eeprom.n2682\
        );

    \I__4441\ : InMux
    port map (
            O => \N__22157\,
            I => \N__22152\
        );

    \I__4440\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22149\
        );

    \I__4439\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22146\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__22152\,
            I => \eeprom.n2714\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__22149\,
            I => \eeprom.n2714\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__22146\,
            I => \eeprom.n2714\
        );

    \I__4435\ : InMux
    port map (
            O => \N__22139\,
            I => \N__22135\
        );

    \I__4434\ : InMux
    port map (
            O => \N__22138\,
            I => \N__22131\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__22135\,
            I => \N__22128\
        );

    \I__4432\ : InMux
    port map (
            O => \N__22134\,
            I => \N__22125\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__22131\,
            I => \eeprom.n2609\
        );

    \I__4430\ : Odrv4
    port map (
            O => \N__22128\,
            I => \eeprom.n2609\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__22125\,
            I => \eeprom.n2609\
        );

    \I__4428\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__22115\,
            I => \eeprom.n2482\
        );

    \I__4426\ : CascadeMux
    port map (
            O => \N__22112\,
            I => \N__22109\
        );

    \I__4425\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22105\
        );

    \I__4424\ : CascadeMux
    port map (
            O => \N__22108\,
            I => \N__22102\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__22105\,
            I => \N__22099\
        );

    \I__4422\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22096\
        );

    \I__4421\ : Span4Mux_h
    port map (
            O => \N__22099\,
            I => \N__22092\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__22096\,
            I => \N__22089\
        );

    \I__4419\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22086\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__22092\,
            I => \eeprom.n2415\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__22089\,
            I => \eeprom.n2415\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__22086\,
            I => \eeprom.n2415\
        );

    \I__4415\ : CascadeMux
    port map (
            O => \N__22079\,
            I => \eeprom.n13_adj_329_cascade_\
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__22076\,
            I => \eeprom.n2539_cascade_\
        );

    \I__4413\ : CascadeMux
    port map (
            O => \N__22073\,
            I => \N__22070\
        );

    \I__4412\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__22061\,
            I => \eeprom.n2683\
        );

    \I__4408\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__4406\ : Span4Mux_h
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__22049\,
            I => \eeprom.n2681\
        );

    \I__4404\ : InMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__22043\,
            I => \N__22039\
        );

    \I__4402\ : InMux
    port map (
            O => \N__22042\,
            I => \N__22036\
        );

    \I__4401\ : Span4Mux_h
    port map (
            O => \N__22039\,
            I => \N__22031\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__22036\,
            I => \N__22031\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__22031\,
            I => \eeprom.n2713\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__22028\,
            I => \eeprom.n2713_cascade_\
        );

    \I__4397\ : InMux
    port map (
            O => \N__22025\,
            I => \N__22021\
        );

    \I__4396\ : InMux
    port map (
            O => \N__22024\,
            I => \N__22018\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__22015\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__22012\
        );

    \I__4393\ : Span4Mux_h
    port map (
            O => \N__22015\,
            I => \N__22006\
        );

    \I__4392\ : Span4Mux_h
    port map (
            O => \N__22012\,
            I => \N__22006\
        );

    \I__4391\ : InMux
    port map (
            O => \N__22011\,
            I => \N__22003\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__22006\,
            I => \eeprom.n2715\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__22003\,
            I => \eeprom.n2715\
        );

    \I__4388\ : CascadeMux
    port map (
            O => \N__21998\,
            I => \N__21994\
        );

    \I__4387\ : CascadeMux
    port map (
            O => \N__21997\,
            I => \N__21990\
        );

    \I__4386\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21987\
        );

    \I__4385\ : InMux
    port map (
            O => \N__21993\,
            I => \N__21982\
        );

    \I__4384\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21982\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21979\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__21982\,
            I => \eeprom.n2219\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__21979\,
            I => \eeprom.n2219\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__21974\,
            I => \N__21971\
        );

    \I__4379\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21968\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__21968\,
            I => \N__21965\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__21965\,
            I => \N__21962\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__21962\,
            I => \eeprom.n3723\
        );

    \I__4375\ : CascadeMux
    port map (
            O => \N__21959\,
            I => \N__21956\
        );

    \I__4374\ : InMux
    port map (
            O => \N__21956\,
            I => \N__21951\
        );

    \I__4373\ : InMux
    port map (
            O => \N__21955\,
            I => \N__21948\
        );

    \I__4372\ : InMux
    port map (
            O => \N__21954\,
            I => \N__21945\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__21951\,
            I => \eeprom.n2210\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__21948\,
            I => \eeprom.n2210\
        );

    \I__4369\ : LocalMux
    port map (
            O => \N__21945\,
            I => \eeprom.n2210\
        );

    \I__4368\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__21935\,
            I => \eeprom.n6_adj_321\
        );

    \I__4366\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__21929\,
            I => \eeprom.n2483\
        );

    \I__4364\ : InMux
    port map (
            O => \N__21926\,
            I => \N__21922\
        );

    \I__4363\ : CascadeMux
    port map (
            O => \N__21925\,
            I => \N__21918\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__21922\,
            I => \N__21915\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__21921\,
            I => \N__21912\
        );

    \I__4360\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21909\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__21915\,
            I => \N__21906\
        );

    \I__4358\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21903\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__21909\,
            I => \N__21900\
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__21906\,
            I => \eeprom.n2416\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__21903\,
            I => \eeprom.n2416\
        );

    \I__4354\ : Odrv4
    port map (
            O => \N__21900\,
            I => \eeprom.n2416\
        );

    \I__4353\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__21890\,
            I => \eeprom.n2485\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__4350\ : InMux
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__21881\,
            I => \N__21877\
        );

    \I__4348\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21873\
        );

    \I__4347\ : Span4Mux_h
    port map (
            O => \N__21877\,
            I => \N__21870\
        );

    \I__4346\ : InMux
    port map (
            O => \N__21876\,
            I => \N__21867\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__21873\,
            I => \N__21864\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__21870\,
            I => \eeprom.n2418\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__21867\,
            I => \eeprom.n2418\
        );

    \I__4342\ : Odrv4
    port map (
            O => \N__21864\,
            I => \eeprom.n2418\
        );

    \I__4341\ : InMux
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__21851\,
            I => \eeprom.n2477\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__4337\ : InMux
    port map (
            O => \N__21845\,
            I => \N__21841\
        );

    \I__4336\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21838\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__21841\,
            I => \N__21834\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__21838\,
            I => \N__21831\
        );

    \I__4333\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21828\
        );

    \I__4332\ : Odrv4
    port map (
            O => \N__21834\,
            I => \eeprom.n2410\
        );

    \I__4331\ : Odrv4
    port map (
            O => \N__21831\,
            I => \eeprom.n2410\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__21828\,
            I => \eeprom.n2410\
        );

    \I__4329\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21817\
        );

    \I__4328\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21814\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__21817\,
            I => \N__21810\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__21814\,
            I => \N__21807\
        );

    \I__4325\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21804\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__21810\,
            I => \eeprom.n2408\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__21807\,
            I => \eeprom.n2408\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__21804\,
            I => \eeprom.n2408\
        );

    \I__4321\ : InMux
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__21794\,
            I => \N__21791\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__21791\,
            I => \eeprom.n2475\
        );

    \I__4318\ : InMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__21782\,
            I => \eeprom.n2486\
        );

    \I__4315\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__21776\,
            I => \eeprom.n2484\
        );

    \I__4313\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21769\
        );

    \I__4312\ : CascadeMux
    port map (
            O => \N__21772\,
            I => \N__21766\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__21769\,
            I => \N__21762\
        );

    \I__4310\ : InMux
    port map (
            O => \N__21766\,
            I => \N__21759\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__21765\,
            I => \N__21756\
        );

    \I__4308\ : Span4Mux_h
    port map (
            O => \N__21762\,
            I => \N__21753\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__21759\,
            I => \N__21750\
        );

    \I__4306\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21747\
        );

    \I__4305\ : Odrv4
    port map (
            O => \N__21753\,
            I => \eeprom.n2417\
        );

    \I__4304\ : Odrv4
    port map (
            O => \N__21750\,
            I => \eeprom.n2417\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__21747\,
            I => \eeprom.n2417\
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__21740\,
            I => \N__21731\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__21739\,
            I => \N__21728\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__21738\,
            I => \N__21724\
        );

    \I__4299\ : InMux
    port map (
            O => \N__21737\,
            I => \N__21718\
        );

    \I__4298\ : InMux
    port map (
            O => \N__21736\,
            I => \N__21713\
        );

    \I__4297\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21713\
        );

    \I__4296\ : InMux
    port map (
            O => \N__21734\,
            I => \N__21710\
        );

    \I__4295\ : InMux
    port map (
            O => \N__21731\,
            I => \N__21703\
        );

    \I__4294\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21703\
        );

    \I__4293\ : InMux
    port map (
            O => \N__21727\,
            I => \N__21703\
        );

    \I__4292\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21696\
        );

    \I__4291\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21696\
        );

    \I__4290\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21696\
        );

    \I__4289\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21693\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__21718\,
            I => \eeprom.n2242\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__21713\,
            I => \eeprom.n2242\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__21710\,
            I => \eeprom.n2242\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__21703\,
            I => \eeprom.n2242\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__21696\,
            I => \eeprom.n2242\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__21693\,
            I => \eeprom.n2242\
        );

    \I__4282\ : InMux
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__21677\,
            I => \eeprom.n5501\
        );

    \I__4280\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__21671\,
            I => \eeprom.n2081\
        );

    \I__4278\ : InMux
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__21662\,
            I => \eeprom.n2086\
        );

    \I__4275\ : InMux
    port map (
            O => \N__21659\,
            I => \N__21656\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__21653\,
            I => \eeprom.n5061\
        );

    \I__4272\ : CascadeMux
    port map (
            O => \N__21650\,
            I => \eeprom.n2118_cascade_\
        );

    \I__4271\ : InMux
    port map (
            O => \N__21647\,
            I => \N__21644\
        );

    \I__4270\ : LocalMux
    port map (
            O => \N__21644\,
            I => \eeprom.n4788\
        );

    \I__4269\ : CascadeMux
    port map (
            O => \N__21641\,
            I => \N__21637\
        );

    \I__4268\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21633\
        );

    \I__4267\ : InMux
    port map (
            O => \N__21637\,
            I => \N__21630\
        );

    \I__4266\ : InMux
    port map (
            O => \N__21636\,
            I => \N__21627\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__21633\,
            I => \N__21624\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__21630\,
            I => \eeprom.n2212\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__21627\,
            I => \eeprom.n2212\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__21624\,
            I => \eeprom.n2212\
        );

    \I__4261\ : InMux
    port map (
            O => \N__21617\,
            I => \N__21612\
        );

    \I__4260\ : InMux
    port map (
            O => \N__21616\,
            I => \N__21609\
        );

    \I__4259\ : InMux
    port map (
            O => \N__21615\,
            I => \N__21606\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__21612\,
            I => \N__21603\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__21609\,
            I => \N__21600\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__21606\,
            I => \eeprom.n2019\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__21603\,
            I => \eeprom.n2019\
        );

    \I__4254\ : Odrv4
    port map (
            O => \N__21600\,
            I => \eeprom.n2019\
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__4252\ : InMux
    port map (
            O => \N__21590\,
            I => \N__21587\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__4249\ : Odrv4
    port map (
            O => \N__21581\,
            I => \eeprom.n3721\
        );

    \I__4248\ : InMux
    port map (
            O => \N__21578\,
            I => \N__21573\
        );

    \I__4247\ : InMux
    port map (
            O => \N__21577\,
            I => \N__21570\
        );

    \I__4246\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21567\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__21573\,
            I => \N__21560\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__21570\,
            I => \N__21560\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__21567\,
            I => \N__21560\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__21557\,
            I => \N__21554\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__21554\,
            I => \eeprom.n3619\
        );

    \I__4239\ : InMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__21548\,
            I => \eeprom.n2085\
        );

    \I__4237\ : InMux
    port map (
            O => \N__21545\,
            I => \eeprom.n3980\
        );

    \I__4236\ : InMux
    port map (
            O => \N__21542\,
            I => \N__21538\
        );

    \I__4235\ : InMux
    port map (
            O => \N__21541\,
            I => \N__21535\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__21538\,
            I => \eeprom.n2084\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__21535\,
            I => \eeprom.n2084\
        );

    \I__4232\ : InMux
    port map (
            O => \N__21530\,
            I => \eeprom.n3981\
        );

    \I__4231\ : InMux
    port map (
            O => \N__21527\,
            I => \eeprom.n3982\
        );

    \I__4230\ : InMux
    port map (
            O => \N__21524\,
            I => \N__21521\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__21521\,
            I => \eeprom.n2082\
        );

    \I__4228\ : InMux
    port map (
            O => \N__21518\,
            I => \eeprom.n3983\
        );

    \I__4227\ : InMux
    port map (
            O => \N__21515\,
            I => \eeprom.n3984\
        );

    \I__4226\ : InMux
    port map (
            O => \N__21512\,
            I => \N__21509\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__21509\,
            I => \eeprom.n2080\
        );

    \I__4224\ : InMux
    port map (
            O => \N__21506\,
            I => \eeprom.n3985\
        );

    \I__4223\ : InMux
    port map (
            O => \N__21503\,
            I => \eeprom.n3986\
        );

    \I__4222\ : InMux
    port map (
            O => \N__21500\,
            I => \bfn_23_19_0_\
        );

    \I__4221\ : InMux
    port map (
            O => \N__21497\,
            I => \N__21493\
        );

    \I__4220\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21490\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__21493\,
            I => \N__21484\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21484\
        );

    \I__4217\ : InMux
    port map (
            O => \N__21489\,
            I => \N__21481\
        );

    \I__4216\ : Odrv4
    port map (
            O => \N__21484\,
            I => \eeprom.n2704\
        );

    \I__4215\ : LocalMux
    port map (
            O => \N__21481\,
            I => \eeprom.n2704\
        );

    \I__4214\ : CascadeMux
    port map (
            O => \N__21476\,
            I => \N__21466\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__21475\,
            I => \N__21463\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__21474\,
            I => \N__21460\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__21473\,
            I => \N__21457\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__21472\,
            I => \N__21454\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__21471\,
            I => \N__21451\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21448\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__21469\,
            I => \N__21445\
        );

    \I__4206\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21434\
        );

    \I__4205\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21434\
        );

    \I__4204\ : InMux
    port map (
            O => \N__21460\,
            I => \N__21434\
        );

    \I__4203\ : InMux
    port map (
            O => \N__21457\,
            I => \N__21434\
        );

    \I__4202\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21425\
        );

    \I__4201\ : InMux
    port map (
            O => \N__21451\,
            I => \N__21425\
        );

    \I__4200\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21425\
        );

    \I__4199\ : InMux
    port map (
            O => \N__21445\,
            I => \N__21425\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__21444\,
            I => \N__21422\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__21443\,
            I => \N__21419\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__21434\,
            I => \N__21414\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__21425\,
            I => \N__21414\
        );

    \I__4194\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21409\
        );

    \I__4193\ : InMux
    port map (
            O => \N__21419\,
            I => \N__21409\
        );

    \I__4192\ : Odrv4
    port map (
            O => \N__21414\,
            I => \eeprom.n2737\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__21409\,
            I => \eeprom.n2737\
        );

    \I__4190\ : InMux
    port map (
            O => \N__21404\,
            I => \eeprom.n4071\
        );

    \I__4189\ : InMux
    port map (
            O => \N__21401\,
            I => \N__21397\
        );

    \I__4188\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21394\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21391\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__21394\,
            I => \N__21388\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__21391\,
            I => \N__21385\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__21388\,
            I => \eeprom.n2803\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__21385\,
            I => \eeprom.n2803\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__21380\,
            I => \eeprom.n5005_cascade_\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__21377\,
            I => \eeprom.n5009_cascade_\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__21374\,
            I => \eeprom.n2044_cascade_\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__21371\,
            I => \eeprom.n2116_cascade_\
        );

    \I__4178\ : InMux
    port map (
            O => \N__21368\,
            I => \bfn_23_18_0_\
        );

    \I__4177\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21361\
        );

    \I__4176\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21357\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__21361\,
            I => \N__21354\
        );

    \I__4174\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21351\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__21357\,
            I => \N__21348\
        );

    \I__4172\ : Span4Mux_h
    port map (
            O => \N__21354\,
            I => \N__21345\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__21351\,
            I => \N__21340\
        );

    \I__4170\ : Span4Mux_h
    port map (
            O => \N__21348\,
            I => \N__21340\
        );

    \I__4169\ : Odrv4
    port map (
            O => \N__21345\,
            I => \eeprom.n2811\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__21340\,
            I => \eeprom.n2811\
        );

    \I__4167\ : InMux
    port map (
            O => \N__21335\,
            I => \eeprom.n4063\
        );

    \I__4166\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21328\
        );

    \I__4165\ : InMux
    port map (
            O => \N__21331\,
            I => \N__21325\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21319\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__21325\,
            I => \N__21319\
        );

    \I__4162\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21316\
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__21319\,
            I => \eeprom.n2711\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__21316\,
            I => \eeprom.n2711\
        );

    \I__4159\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21305\
        );

    \I__4158\ : InMux
    port map (
            O => \N__21310\,
            I => \N__21305\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21301\
        );

    \I__4156\ : InMux
    port map (
            O => \N__21304\,
            I => \N__21298\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__21301\,
            I => \N__21293\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__21298\,
            I => \N__21293\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__21293\,
            I => \eeprom.n2810\
        );

    \I__4152\ : InMux
    port map (
            O => \N__21290\,
            I => \bfn_22_26_0_\
        );

    \I__4151\ : InMux
    port map (
            O => \N__21287\,
            I => \N__21283\
        );

    \I__4150\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21280\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__21283\,
            I => \eeprom.n2710\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__21280\,
            I => \eeprom.n2710\
        );

    \I__4147\ : InMux
    port map (
            O => \N__21275\,
            I => \N__21270\
        );

    \I__4146\ : CascadeMux
    port map (
            O => \N__21274\,
            I => \N__21267\
        );

    \I__4145\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21264\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__21270\,
            I => \N__21261\
        );

    \I__4143\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21258\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__21264\,
            I => \N__21255\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__21261\,
            I => \N__21252\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__21258\,
            I => \N__21249\
        );

    \I__4139\ : Span4Mux_h
    port map (
            O => \N__21255\,
            I => \N__21246\
        );

    \I__4138\ : Odrv4
    port map (
            O => \N__21252\,
            I => \eeprom.n2809\
        );

    \I__4137\ : Odrv4
    port map (
            O => \N__21249\,
            I => \eeprom.n2809\
        );

    \I__4136\ : Odrv4
    port map (
            O => \N__21246\,
            I => \eeprom.n2809\
        );

    \I__4135\ : InMux
    port map (
            O => \N__21239\,
            I => \eeprom.n4065\
        );

    \I__4134\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21232\
        );

    \I__4133\ : InMux
    port map (
            O => \N__21235\,
            I => \N__21229\
        );

    \I__4132\ : LocalMux
    port map (
            O => \N__21232\,
            I => \N__21224\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__21229\,
            I => \N__21224\
        );

    \I__4130\ : Span4Mux_h
    port map (
            O => \N__21224\,
            I => \N__21220\
        );

    \I__4129\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21217\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__21220\,
            I => \eeprom.n2709\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__21217\,
            I => \eeprom.n2709\
        );

    \I__4126\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21207\
        );

    \I__4125\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21204\
        );

    \I__4124\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21201\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__21207\,
            I => \N__21194\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__21204\,
            I => \N__21194\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__21201\,
            I => \N__21194\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__21191\,
            I => \eeprom.n2808\
        );

    \I__4118\ : InMux
    port map (
            O => \N__21188\,
            I => \eeprom.n4066\
        );

    \I__4117\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21181\
        );

    \I__4116\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21178\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__21181\,
            I => \N__21172\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__21178\,
            I => \N__21172\
        );

    \I__4113\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21169\
        );

    \I__4112\ : Odrv12
    port map (
            O => \N__21172\,
            I => \eeprom.n2708\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__21169\,
            I => \eeprom.n2708\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__21164\,
            I => \N__21160\
        );

    \I__4109\ : InMux
    port map (
            O => \N__21163\,
            I => \N__21156\
        );

    \I__4108\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21153\
        );

    \I__4107\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21150\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__21156\,
            I => \N__21143\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__21153\,
            I => \N__21143\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__21150\,
            I => \N__21143\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__4102\ : Odrv4
    port map (
            O => \N__21140\,
            I => \eeprom.n2807\
        );

    \I__4101\ : InMux
    port map (
            O => \N__21137\,
            I => \eeprom.n4067\
        );

    \I__4100\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21130\
        );

    \I__4099\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21127\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__21130\,
            I => \N__21123\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__21127\,
            I => \N__21120\
        );

    \I__4096\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21117\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__21123\,
            I => \eeprom.n2707\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__21120\,
            I => \eeprom.n2707\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__21117\,
            I => \eeprom.n2707\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__21110\,
            I => \N__21106\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__21109\,
            I => \N__21103\
        );

    \I__4090\ : InMux
    port map (
            O => \N__21106\,
            I => \N__21099\
        );

    \I__4089\ : InMux
    port map (
            O => \N__21103\,
            I => \N__21096\
        );

    \I__4088\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21093\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__21099\,
            I => \N__21088\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__21096\,
            I => \N__21088\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__21093\,
            I => \N__21085\
        );

    \I__4084\ : Span4Mux_h
    port map (
            O => \N__21088\,
            I => \N__21082\
        );

    \I__4083\ : Odrv4
    port map (
            O => \N__21085\,
            I => \eeprom.n2806\
        );

    \I__4082\ : Odrv4
    port map (
            O => \N__21082\,
            I => \eeprom.n2806\
        );

    \I__4081\ : InMux
    port map (
            O => \N__21077\,
            I => \eeprom.n4068\
        );

    \I__4080\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21069\
        );

    \I__4079\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21066\
        );

    \I__4078\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21063\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__21069\,
            I => \N__21060\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21057\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__21063\,
            I => \N__21052\
        );

    \I__4074\ : Span4Mux_h
    port map (
            O => \N__21060\,
            I => \N__21052\
        );

    \I__4073\ : Odrv4
    port map (
            O => \N__21057\,
            I => \eeprom.n2805\
        );

    \I__4072\ : Odrv4
    port map (
            O => \N__21052\,
            I => \eeprom.n2805\
        );

    \I__4071\ : InMux
    port map (
            O => \N__21047\,
            I => \eeprom.n4069\
        );

    \I__4070\ : InMux
    port map (
            O => \N__21044\,
            I => \N__21040\
        );

    \I__4069\ : InMux
    port map (
            O => \N__21043\,
            I => \N__21037\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__21040\,
            I => \N__21032\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__21037\,
            I => \N__21032\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__21032\,
            I => \eeprom.n2705\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__21029\,
            I => \N__21025\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__21028\,
            I => \N__21021\
        );

    \I__4063\ : InMux
    port map (
            O => \N__21025\,
            I => \N__21018\
        );

    \I__4062\ : InMux
    port map (
            O => \N__21024\,
            I => \N__21015\
        );

    \I__4061\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21012\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__21018\,
            I => \N__21007\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__21015\,
            I => \N__21007\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__21012\,
            I => \N__21004\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__21007\,
            I => \N__21001\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__21004\,
            I => \eeprom.n2804\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__21001\,
            I => \eeprom.n2804\
        );

    \I__4054\ : InMux
    port map (
            O => \N__20996\,
            I => \eeprom.n4070\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__20993\,
            I => \eeprom.n2737_cascade_\
        );

    \I__4052\ : InMux
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__20987\,
            I => \N__20983\
        );

    \I__4050\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20979\
        );

    \I__4049\ : Span4Mux_v
    port map (
            O => \N__20983\,
            I => \N__20976\
        );

    \I__4048\ : InMux
    port map (
            O => \N__20982\,
            I => \N__20973\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__20979\,
            I => \N__20970\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__20976\,
            I => \eeprom.n2818\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__20973\,
            I => \eeprom.n2818\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__20970\,
            I => \eeprom.n2818\
        );

    \I__4043\ : InMux
    port map (
            O => \N__20963\,
            I => \bfn_22_25_0_\
        );

    \I__4042\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20955\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__20959\,
            I => \N__20952\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__20958\,
            I => \N__20949\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__20955\,
            I => \N__20946\
        );

    \I__4038\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20943\
        );

    \I__4037\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20940\
        );

    \I__4036\ : Span4Mux_h
    port map (
            O => \N__20946\,
            I => \N__20935\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__20943\,
            I => \N__20935\
        );

    \I__4034\ : LocalMux
    port map (
            O => \N__20940\,
            I => \eeprom.n2817\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__20935\,
            I => \eeprom.n2817\
        );

    \I__4032\ : InMux
    port map (
            O => \N__20930\,
            I => \eeprom.n4057\
        );

    \I__4031\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20923\
        );

    \I__4030\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20920\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__20923\,
            I => \N__20917\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20913\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__20917\,
            I => \N__20910\
        );

    \I__4026\ : InMux
    port map (
            O => \N__20916\,
            I => \N__20907\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__20913\,
            I => \eeprom.n2717\
        );

    \I__4024\ : Odrv4
    port map (
            O => \N__20910\,
            I => \eeprom.n2717\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__20907\,
            I => \eeprom.n2717\
        );

    \I__4022\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__20897\,
            I => \N__20893\
        );

    \I__4020\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__4019\ : Span4Mux_h
    port map (
            O => \N__20893\,
            I => \N__20884\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__20890\,
            I => \N__20884\
        );

    \I__4017\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20881\
        );

    \I__4016\ : Odrv4
    port map (
            O => \N__20884\,
            I => \eeprom.n2816\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__20881\,
            I => \eeprom.n2816\
        );

    \I__4014\ : InMux
    port map (
            O => \N__20876\,
            I => \eeprom.n4058\
        );

    \I__4013\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20869\
        );

    \I__4012\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20866\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__20869\,
            I => \N__20861\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__20866\,
            I => \N__20861\
        );

    \I__4009\ : Odrv4
    port map (
            O => \N__20861\,
            I => \eeprom.n2716\
        );

    \I__4008\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20855\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__20855\,
            I => \N__20851\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__20854\,
            I => \N__20848\
        );

    \I__4005\ : Span4Mux_h
    port map (
            O => \N__20851\,
            I => \N__20844\
        );

    \I__4004\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20841\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__20847\,
            I => \N__20838\
        );

    \I__4002\ : Sp12to4
    port map (
            O => \N__20844\,
            I => \N__20835\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__20841\,
            I => \N__20832\
        );

    \I__4000\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20829\
        );

    \I__3999\ : Odrv12
    port map (
            O => \N__20835\,
            I => \eeprom.n2815\
        );

    \I__3998\ : Odrv4
    port map (
            O => \N__20832\,
            I => \eeprom.n2815\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__20829\,
            I => \eeprom.n2815\
        );

    \I__3996\ : InMux
    port map (
            O => \N__20822\,
            I => \eeprom.n4059\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__3994\ : InMux
    port map (
            O => \N__20816\,
            I => \N__20812\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__20815\,
            I => \N__20809\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__20812\,
            I => \N__20806\
        );

    \I__3991\ : InMux
    port map (
            O => \N__20809\,
            I => \N__20803\
        );

    \I__3990\ : Span4Mux_h
    port map (
            O => \N__20806\,
            I => \N__20797\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__20803\,
            I => \N__20797\
        );

    \I__3988\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20794\
        );

    \I__3987\ : Odrv4
    port map (
            O => \N__20797\,
            I => \eeprom.n2814\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__20794\,
            I => \eeprom.n2814\
        );

    \I__3985\ : InMux
    port map (
            O => \N__20789\,
            I => \eeprom.n4060\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__20786\,
            I => \N__20782\
        );

    \I__3983\ : InMux
    port map (
            O => \N__20785\,
            I => \N__20779\
        );

    \I__3982\ : InMux
    port map (
            O => \N__20782\,
            I => \N__20775\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__20779\,
            I => \N__20772\
        );

    \I__3980\ : InMux
    port map (
            O => \N__20778\,
            I => \N__20769\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__20775\,
            I => \eeprom.n2813\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__20772\,
            I => \eeprom.n2813\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__20769\,
            I => \eeprom.n2813\
        );

    \I__3976\ : InMux
    port map (
            O => \N__20762\,
            I => \eeprom.n4061\
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__20759\,
            I => \N__20751\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__20758\,
            I => \N__20748\
        );

    \I__3973\ : CascadeMux
    port map (
            O => \N__20757\,
            I => \N__20745\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__20756\,
            I => \N__20742\
        );

    \I__3971\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \N__20739\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__20754\,
            I => \N__20736\
        );

    \I__3969\ : InMux
    port map (
            O => \N__20751\,
            I => \N__20731\
        );

    \I__3968\ : InMux
    port map (
            O => \N__20748\,
            I => \N__20731\
        );

    \I__3967\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20722\
        );

    \I__3966\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20722\
        );

    \I__3965\ : InMux
    port map (
            O => \N__20739\,
            I => \N__20722\
        );

    \I__3964\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20722\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__20731\,
            I => \eeprom.n5575\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__20722\,
            I => \eeprom.n5575\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__20717\,
            I => \N__20714\
        );

    \I__3960\ : InMux
    port map (
            O => \N__20714\,
            I => \N__20711\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20706\
        );

    \I__3958\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20701\
        );

    \I__3957\ : InMux
    port map (
            O => \N__20709\,
            I => \N__20701\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__20706\,
            I => \eeprom.n2812\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__20701\,
            I => \eeprom.n2812\
        );

    \I__3954\ : InMux
    port map (
            O => \N__20696\,
            I => \eeprom.n4062\
        );

    \I__3953\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20688\
        );

    \I__3952\ : InMux
    port map (
            O => \N__20692\,
            I => \N__20685\
        );

    \I__3951\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20682\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__20688\,
            I => \eeprom.n2712\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__20685\,
            I => \eeprom.n2712\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__20682\,
            I => \eeprom.n2712\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__20675\,
            I => \eeprom.n2638_cascade_\
        );

    \I__3946\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20669\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__20669\,
            I => \eeprom.n2684\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__20666\,
            I => \eeprom.n2716_cascade_\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__20663\,
            I => \N__20660\
        );

    \I__3942\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20657\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__20657\,
            I => \eeprom.n2680\
        );

    \I__3940\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20651\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__20651\,
            I => \eeprom.n2679\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__20648\,
            I => \N__20645\
        );

    \I__3937\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20642\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__20642\,
            I => \eeprom.n2676\
        );

    \I__3935\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20636\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__20636\,
            I => \eeprom.n2675\
        );

    \I__3933\ : CascadeMux
    port map (
            O => \N__20633\,
            I => \N__20630\
        );

    \I__3932\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20627\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__20627\,
            I => \eeprom.n2673\
        );

    \I__3930\ : CascadeMux
    port map (
            O => \N__20624\,
            I => \eeprom.n2705_cascade_\
        );

    \I__3929\ : InMux
    port map (
            O => \N__20621\,
            I => \N__20618\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__20618\,
            I => \eeprom.n17_adj_339\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__20615\,
            I => \eeprom.n16_adj_338_cascade_\
        );

    \I__3926\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20609\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20604\
        );

    \I__3924\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20599\
        );

    \I__3923\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20599\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__20604\,
            I => \eeprom.n2413\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__20599\,
            I => \eeprom.n2413\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__20594\,
            I => \N__20591\
        );

    \I__3919\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20588\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__20588\,
            I => \eeprom.n2480\
        );

    \I__3917\ : InMux
    port map (
            O => \N__20585\,
            I => \eeprom.n4023\
        );

    \I__3916\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20578\
        );

    \I__3915\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20574\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__20578\,
            I => \N__20571\
        );

    \I__3913\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20568\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20565\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__20571\,
            I => \eeprom.n2412\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__20568\,
            I => \eeprom.n2412\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__20565\,
            I => \eeprom.n2412\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__20558\,
            I => \N__20555\
        );

    \I__3907\ : InMux
    port map (
            O => \N__20555\,
            I => \N__20552\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__20552\,
            I => \eeprom.n2479\
        );

    \I__3905\ : InMux
    port map (
            O => \N__20549\,
            I => \eeprom.n4024\
        );

    \I__3904\ : InMux
    port map (
            O => \N__20546\,
            I => \bfn_22_23_0_\
        );

    \I__3903\ : InMux
    port map (
            O => \N__20543\,
            I => \eeprom.n4026\
        );

    \I__3902\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20537\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__20537\,
            I => \N__20532\
        );

    \I__3900\ : InMux
    port map (
            O => \N__20536\,
            I => \N__20527\
        );

    \I__3899\ : InMux
    port map (
            O => \N__20535\,
            I => \N__20527\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__20532\,
            I => \eeprom.n2409\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__20527\,
            I => \eeprom.n2409\
        );

    \I__3896\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20519\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20516\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__20516\,
            I => \eeprom.n2476\
        );

    \I__3893\ : InMux
    port map (
            O => \N__20513\,
            I => \eeprom.n4027\
        );

    \I__3892\ : InMux
    port map (
            O => \N__20510\,
            I => \eeprom.n4028\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__20507\,
            I => \N__20504\
        );

    \I__3890\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20501\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__20501\,
            I => \N__20497\
        );

    \I__3888\ : InMux
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__3887\ : Odrv4
    port map (
            O => \N__20497\,
            I => \eeprom.n2407\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__20494\,
            I => \eeprom.n2407\
        );

    \I__3885\ : InMux
    port map (
            O => \N__20489\,
            I => \eeprom.n4029\
        );

    \I__3884\ : CascadeMux
    port map (
            O => \N__20486\,
            I => \eeprom.n2440_cascade_\
        );

    \I__3883\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20480\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__20480\,
            I => \eeprom.n5071\
        );

    \I__3881\ : InMux
    port map (
            O => \N__20477\,
            I => \bfn_22_22_0_\
        );

    \I__3880\ : InMux
    port map (
            O => \N__20474\,
            I => \eeprom.n4018\
        );

    \I__3879\ : InMux
    port map (
            O => \N__20471\,
            I => \eeprom.n4019\
        );

    \I__3878\ : InMux
    port map (
            O => \N__20468\,
            I => \eeprom.n4020\
        );

    \I__3877\ : InMux
    port map (
            O => \N__20465\,
            I => \eeprom.n4021\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__20462\,
            I => \N__20459\
        );

    \I__3875\ : InMux
    port map (
            O => \N__20459\,
            I => \N__20456\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__20456\,
            I => \N__20451\
        );

    \I__3873\ : InMux
    port map (
            O => \N__20455\,
            I => \N__20446\
        );

    \I__3872\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20446\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__20451\,
            I => \eeprom.n2414\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__20446\,
            I => \eeprom.n2414\
        );

    \I__3869\ : InMux
    port map (
            O => \N__20441\,
            I => \N__20438\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__20438\,
            I => \eeprom.n2481\
        );

    \I__3867\ : InMux
    port map (
            O => \N__20435\,
            I => \eeprom.n4022\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__20432\,
            I => \eeprom.n2309_cascade_\
        );

    \I__3865\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20425\
        );

    \I__3864\ : InMux
    port map (
            O => \N__20428\,
            I => \N__20422\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__20425\,
            I => \N__20416\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__20422\,
            I => \N__20416\
        );

    \I__3861\ : InMux
    port map (
            O => \N__20421\,
            I => \N__20413\
        );

    \I__3860\ : Span4Mux_h
    port map (
            O => \N__20416\,
            I => \N__20408\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__20413\,
            I => \N__20408\
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__20408\,
            I => \eeprom.n2308\
        );

    \I__3857\ : InMux
    port map (
            O => \N__20405\,
            I => \N__20401\
        );

    \I__3856\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20398\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__20401\,
            I => \N__20393\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__20398\,
            I => \N__20393\
        );

    \I__3853\ : Span4Mux_v
    port map (
            O => \N__20393\,
            I => \N__20389\
        );

    \I__3852\ : InMux
    port map (
            O => \N__20392\,
            I => \N__20386\
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__20389\,
            I => \eeprom.n2312\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__20386\,
            I => \eeprom.n2312\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__20381\,
            I => \eeprom.n8_adj_322_cascade_\
        );

    \I__3848\ : InMux
    port map (
            O => \N__20378\,
            I => \N__20375\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__20375\,
            I => \eeprom.n7_adj_323\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__20372\,
            I => \N__20364\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__20371\,
            I => \N__20361\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__20370\,
            I => \N__20358\
        );

    \I__3843\ : CascadeMux
    port map (
            O => \N__20369\,
            I => \N__20355\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__20368\,
            I => \N__20352\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__20367\,
            I => \N__20349\
        );

    \I__3840\ : InMux
    port map (
            O => \N__20364\,
            I => \N__20344\
        );

    \I__3839\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20344\
        );

    \I__3838\ : InMux
    port map (
            O => \N__20358\,
            I => \N__20339\
        );

    \I__3837\ : InMux
    port map (
            O => \N__20355\,
            I => \N__20339\
        );

    \I__3836\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20334\
        );

    \I__3835\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20334\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__20344\,
            I => \eeprom.n2341\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__20339\,
            I => \eeprom.n2341\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__20334\,
            I => \eeprom.n2341\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__20327\,
            I => \eeprom.n2341_cascade_\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__20324\,
            I => \N__20316\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__20323\,
            I => \N__20313\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__20322\,
            I => \N__20310\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__20321\,
            I => \N__20307\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__20320\,
            I => \N__20304\
        );

    \I__3825\ : CascadeMux
    port map (
            O => \N__20319\,
            I => \N__20301\
        );

    \I__3824\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20296\
        );

    \I__3823\ : InMux
    port map (
            O => \N__20313\,
            I => \N__20296\
        );

    \I__3822\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20287\
        );

    \I__3821\ : InMux
    port map (
            O => \N__20307\,
            I => \N__20287\
        );

    \I__3820\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20287\
        );

    \I__3819\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20287\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__20296\,
            I => \eeprom.n5576\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__20287\,
            I => \eeprom.n5576\
        );

    \I__3816\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__20276\,
            I => \eeprom.n2279\
        );

    \I__3813\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20268\
        );

    \I__3812\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20265\
        );

    \I__3811\ : InMux
    port map (
            O => \N__20271\,
            I => \N__20262\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__20268\,
            I => \eeprom.n2311\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__20265\,
            I => \eeprom.n2311\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__20262\,
            I => \eeprom.n2311\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__20255\,
            I => \eeprom.n5073_cascade_\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__20252\,
            I => \eeprom.n4782_cascade_\
        );

    \I__3805\ : CascadeMux
    port map (
            O => \N__20249\,
            I => \eeprom.n12_cascade_\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__20246\,
            I => \eeprom.n2242_cascade_\
        );

    \I__3803\ : InMux
    port map (
            O => \N__20243\,
            I => \N__20240\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__20240\,
            I => \N__20237\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__20237\,
            I => \eeprom.n2282\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__20234\,
            I => \eeprom.n5400_cascade_\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__20231\,
            I => \N__20227\
        );

    \I__3798\ : InMux
    port map (
            O => \N__20230\,
            I => \N__20223\
        );

    \I__3797\ : InMux
    port map (
            O => \N__20227\,
            I => \N__20220\
        );

    \I__3796\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20217\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__20223\,
            I => \eeprom.n2217\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__20220\,
            I => \eeprom.n2217\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__20217\,
            I => \eeprom.n2217\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__20210\,
            I => \N__20207\
        );

    \I__3791\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20204\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__20204\,
            I => \N__20201\
        );

    \I__3789\ : Odrv4
    port map (
            O => \N__20201\,
            I => \eeprom.n2284\
        );

    \I__3788\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20195\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__20195\,
            I => \N__20192\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__20192\,
            I => \eeprom.n2280\
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__20189\,
            I => \N__20186\
        );

    \I__3784\ : InMux
    port map (
            O => \N__20186\,
            I => \N__20181\
        );

    \I__3783\ : InMux
    port map (
            O => \N__20185\,
            I => \N__20176\
        );

    \I__3782\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20176\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__20181\,
            I => \eeprom.n2213\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__20176\,
            I => \eeprom.n2213\
        );

    \I__3779\ : InMux
    port map (
            O => \N__20171\,
            I => \N__20168\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__20168\,
            I => \eeprom.n5405\
        );

    \I__3777\ : InMux
    port map (
            O => \N__20165\,
            I => \N__20160\
        );

    \I__3776\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20157\
        );

    \I__3775\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20154\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__20160\,
            I => \eeprom.n2316\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__20157\,
            I => \eeprom.n2316\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__20154\,
            I => \eeprom.n2316\
        );

    \I__3771\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20142\
        );

    \I__3770\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20139\
        );

    \I__3769\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20136\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__20142\,
            I => \eeprom.n2317\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__20139\,
            I => \eeprom.n2317\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__20136\,
            I => \eeprom.n2317\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__20129\,
            I => \N__20124\
        );

    \I__3764\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20121\
        );

    \I__3763\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20118\
        );

    \I__3762\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20115\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__20121\,
            I => \eeprom.n2314\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__20118\,
            I => \eeprom.n2314\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__20115\,
            I => \eeprom.n2314\
        );

    \I__3758\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20103\
        );

    \I__3757\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20100\
        );

    \I__3756\ : InMux
    port map (
            O => \N__20106\,
            I => \N__20097\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__20103\,
            I => \eeprom.n2318\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__20100\,
            I => \eeprom.n2318\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__20097\,
            I => \eeprom.n2318\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__20090\,
            I => \eeprom.n5085_cascade_\
        );

    \I__3751\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20082\
        );

    \I__3750\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20079\
        );

    \I__3749\ : InMux
    port map (
            O => \N__20085\,
            I => \N__20076\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__20082\,
            I => \N__20071\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__20079\,
            I => \N__20071\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__20076\,
            I => \N__20068\
        );

    \I__3745\ : Odrv12
    port map (
            O => \N__20071\,
            I => \eeprom.n2310\
        );

    \I__3744\ : Odrv4
    port map (
            O => \N__20068\,
            I => \eeprom.n2310\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__20063\,
            I => \N__20058\
        );

    \I__3742\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20055\
        );

    \I__3741\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20052\
        );

    \I__3740\ : InMux
    port map (
            O => \N__20058\,
            I => \N__20049\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__20055\,
            I => \eeprom.n2315\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__20052\,
            I => \eeprom.n2315\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__20049\,
            I => \eeprom.n2315\
        );

    \I__3736\ : InMux
    port map (
            O => \N__20042\,
            I => \N__20037\
        );

    \I__3735\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20034\
        );

    \I__3734\ : InMux
    port map (
            O => \N__20040\,
            I => \N__20031\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__20037\,
            I => \eeprom.n2313\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__20034\,
            I => \eeprom.n2313\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__20031\,
            I => \eeprom.n2313\
        );

    \I__3730\ : InMux
    port map (
            O => \N__20024\,
            I => \N__20021\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__20021\,
            I => \eeprom.n5081\
        );

    \I__3728\ : InMux
    port map (
            O => \N__20018\,
            I => \N__20015\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__20015\,
            I => \N__20012\
        );

    \I__3726\ : Odrv12
    port map (
            O => \N__20012\,
            I => \eeprom.n2277\
        );

    \I__3725\ : InMux
    port map (
            O => \N__20009\,
            I => \N__20005\
        );

    \I__3724\ : InMux
    port map (
            O => \N__20008\,
            I => \N__20002\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__20005\,
            I => \eeprom.n2309\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__20002\,
            I => \eeprom.n2309\
        );

    \I__3721\ : InMux
    port map (
            O => \N__19997\,
            I => \eeprom.n4005\
        );

    \I__3720\ : InMux
    port map (
            O => \N__19994\,
            I => \eeprom.n4006\
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__19991\,
            I => \N__19987\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__19990\,
            I => \N__19984\
        );

    \I__3717\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19980\
        );

    \I__3716\ : InMux
    port map (
            O => \N__19984\,
            I => \N__19977\
        );

    \I__3715\ : InMux
    port map (
            O => \N__19983\,
            I => \N__19974\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__19980\,
            I => \eeprom.n2216\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__19977\,
            I => \eeprom.n2216\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__19974\,
            I => \eeprom.n2216\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__19967\,
            I => \eeprom.n2143_cascade_\
        );

    \I__3710\ : InMux
    port map (
            O => \N__19964\,
            I => \N__19961\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__19961\,
            I => \N__19958\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__19958\,
            I => \eeprom.n2286\
        );

    \I__3707\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19951\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__19954\,
            I => \N__19947\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__19951\,
            I => \N__19944\
        );

    \I__3704\ : InMux
    port map (
            O => \N__19950\,
            I => \N__19941\
        );

    \I__3703\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19938\
        );

    \I__3702\ : Odrv4
    port map (
            O => \N__19944\,
            I => \eeprom.n2218\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__19941\,
            I => \eeprom.n2218\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__19938\,
            I => \eeprom.n2218\
        );

    \I__3699\ : InMux
    port map (
            O => \N__19931\,
            I => \N__19928\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__19928\,
            I => \eeprom.n5045\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__19925\,
            I => \N__19922\
        );

    \I__3696\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19918\
        );

    \I__3695\ : InMux
    port map (
            O => \N__19921\,
            I => \N__19915\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__19918\,
            I => \eeprom.n2211\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__19915\,
            I => \eeprom.n2211\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__19910\,
            I => \eeprom.n4797_cascade_\
        );

    \I__3691\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19904\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19901\
        );

    \I__3689\ : Span4Mux_h
    port map (
            O => \N__19901\,
            I => \N__19898\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__19898\,
            I => \eeprom.n2285\
        );

    \I__3687\ : InMux
    port map (
            O => \N__19895\,
            I => \eeprom.n3997\
        );

    \I__3686\ : InMux
    port map (
            O => \N__19892\,
            I => \eeprom.n3998\
        );

    \I__3685\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__19883\,
            I => \eeprom.n2283\
        );

    \I__3682\ : InMux
    port map (
            O => \N__19880\,
            I => \eeprom.n3999\
        );

    \I__3681\ : CascadeMux
    port map (
            O => \N__19877\,
            I => \N__19874\
        );

    \I__3680\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19870\
        );

    \I__3679\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19867\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__19870\,
            I => \eeprom.n2215\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__19867\,
            I => \eeprom.n2215\
        );

    \I__3676\ : InMux
    port map (
            O => \N__19862\,
            I => \eeprom.n4000\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__19859\,
            I => \N__19856\
        );

    \I__3674\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19852\
        );

    \I__3673\ : InMux
    port map (
            O => \N__19855\,
            I => \N__19849\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__19852\,
            I => \N__19846\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__19849\,
            I => \eeprom.n2214\
        );

    \I__3670\ : Odrv4
    port map (
            O => \N__19846\,
            I => \eeprom.n2214\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__19841\,
            I => \N__19838\
        );

    \I__3668\ : InMux
    port map (
            O => \N__19838\,
            I => \N__19835\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19832\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__19832\,
            I => \eeprom.n2281\
        );

    \I__3665\ : InMux
    port map (
            O => \N__19829\,
            I => \eeprom.n4001\
        );

    \I__3664\ : InMux
    port map (
            O => \N__19826\,
            I => \eeprom.n4002\
        );

    \I__3663\ : InMux
    port map (
            O => \N__19823\,
            I => \eeprom.n4003\
        );

    \I__3662\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19817\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__19817\,
            I => \eeprom.n2278\
        );

    \I__3660\ : InMux
    port map (
            O => \N__19814\,
            I => \bfn_22_18_0_\
        );

    \I__3659\ : InMux
    port map (
            O => \N__19811\,
            I => \eeprom.n4085\
        );

    \I__3658\ : InMux
    port map (
            O => \N__19808\,
            I => \eeprom.n4086\
        );

    \I__3657\ : InMux
    port map (
            O => \N__19805\,
            I => \bfn_21_29_0_\
        );

    \I__3656\ : InMux
    port map (
            O => \N__19802\,
            I => \N__19799\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19796\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__19796\,
            I => \eeprom.n2902\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__19793\,
            I => \eeprom.n2902_cascade_\
        );

    \I__3652\ : InMux
    port map (
            O => \N__19790\,
            I => \N__19787\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__19787\,
            I => \N__19784\
        );

    \I__3650\ : Odrv4
    port map (
            O => \N__19784\,
            I => \eeprom.n19_adj_327\
        );

    \I__3649\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19778\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__19778\,
            I => \eeprom.n2872\
        );

    \I__3647\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19772\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__19772\,
            I => \N__19767\
        );

    \I__3645\ : InMux
    port map (
            O => \N__19771\,
            I => \N__19764\
        );

    \I__3644\ : InMux
    port map (
            O => \N__19770\,
            I => \N__19761\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__19767\,
            I => \eeprom.n2904\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__19764\,
            I => \eeprom.n2904\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__19761\,
            I => \eeprom.n2904\
        );

    \I__3640\ : InMux
    port map (
            O => \N__19754\,
            I => \N__19751\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__19751\,
            I => \eeprom.n2873\
        );

    \I__3638\ : InMux
    port map (
            O => \N__19748\,
            I => \N__19745\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__19745\,
            I => \N__19742\
        );

    \I__3636\ : Span4Mux_s3_v
    port map (
            O => \N__19742\,
            I => \N__19737\
        );

    \I__3635\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19734\
        );

    \I__3634\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19731\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__19737\,
            I => \eeprom.n2905\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__19734\,
            I => \eeprom.n2905\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__19731\,
            I => \eeprom.n2905\
        );

    \I__3630\ : InMux
    port map (
            O => \N__19724\,
            I => \N__19721\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__19721\,
            I => \eeprom.n2871\
        );

    \I__3628\ : InMux
    port map (
            O => \N__19718\,
            I => \N__19715\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__19715\,
            I => \N__19711\
        );

    \I__3626\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19708\
        );

    \I__3625\ : Span4Mux_v
    port map (
            O => \N__19711\,
            I => \N__19704\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__19708\,
            I => \N__19701\
        );

    \I__3623\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19698\
        );

    \I__3622\ : Odrv4
    port map (
            O => \N__19704\,
            I => \eeprom.n2903\
        );

    \I__3621\ : Odrv4
    port map (
            O => \N__19701\,
            I => \eeprom.n2903\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__19698\,
            I => \eeprom.n2903\
        );

    \I__3619\ : CascadeMux
    port map (
            O => \N__19691\,
            I => \N__19688\
        );

    \I__3618\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19685\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__19685\,
            I => \eeprom.n2875\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__19682\,
            I => \N__19675\
        );

    \I__3615\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19667\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__19680\,
            I => \N__19663\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__19679\,
            I => \N__19660\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__19678\,
            I => \N__19657\
        );

    \I__3611\ : InMux
    port map (
            O => \N__19675\,
            I => \N__19651\
        );

    \I__3610\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19651\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__19673\,
            I => \N__19648\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__19672\,
            I => \N__19645\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__19671\,
            I => \N__19639\
        );

    \I__3606\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19635\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19632\
        );

    \I__3604\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19621\
        );

    \I__3603\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19621\
        );

    \I__3602\ : InMux
    port map (
            O => \N__19660\,
            I => \N__19621\
        );

    \I__3601\ : InMux
    port map (
            O => \N__19657\,
            I => \N__19621\
        );

    \I__3600\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19621\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__19651\,
            I => \N__19618\
        );

    \I__3598\ : InMux
    port map (
            O => \N__19648\,
            I => \N__19609\
        );

    \I__3597\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19609\
        );

    \I__3596\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19609\
        );

    \I__3595\ : InMux
    port map (
            O => \N__19643\,
            I => \N__19609\
        );

    \I__3594\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19602\
        );

    \I__3593\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19602\
        );

    \I__3592\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19602\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__19635\,
            I => \eeprom.n2836\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__19632\,
            I => \eeprom.n2836\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__19621\,
            I => \eeprom.n2836\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__19618\,
            I => \eeprom.n2836\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__19609\,
            I => \eeprom.n2836\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__19602\,
            I => \eeprom.n2836\
        );

    \I__3585\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19585\
        );

    \I__3584\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19582\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__19585\,
            I => \N__19579\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__19582\,
            I => \N__19575\
        );

    \I__3581\ : Span4Mux_h
    port map (
            O => \N__19579\,
            I => \N__19572\
        );

    \I__3580\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19569\
        );

    \I__3579\ : Span4Mux_h
    port map (
            O => \N__19575\,
            I => \N__19566\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__19572\,
            I => \eeprom.n2907\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__19569\,
            I => \eeprom.n2907\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__19566\,
            I => \eeprom.n2907\
        );

    \I__3575\ : InMux
    port map (
            O => \N__19559\,
            I => \bfn_22_17_0_\
        );

    \I__3574\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19550\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__19550\,
            I => \eeprom.n2880\
        );

    \I__3571\ : InMux
    port map (
            O => \N__19547\,
            I => \eeprom.n4077\
        );

    \I__3570\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19541\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__19541\,
            I => \eeprom.n2879\
        );

    \I__3568\ : InMux
    port map (
            O => \N__19538\,
            I => \eeprom.n4078\
        );

    \I__3567\ : InMux
    port map (
            O => \N__19535\,
            I => \N__19532\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__19532\,
            I => \eeprom.n2878\
        );

    \I__3565\ : InMux
    port map (
            O => \N__19529\,
            I => \bfn_21_28_0_\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__19526\,
            I => \N__19523\
        );

    \I__3563\ : InMux
    port map (
            O => \N__19523\,
            I => \N__19520\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__19520\,
            I => \eeprom.n2877\
        );

    \I__3561\ : InMux
    port map (
            O => \N__19517\,
            I => \eeprom.n4080\
        );

    \I__3560\ : InMux
    port map (
            O => \N__19514\,
            I => \N__19511\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__3558\ : Odrv4
    port map (
            O => \N__19508\,
            I => \eeprom.n2876\
        );

    \I__3557\ : InMux
    port map (
            O => \N__19505\,
            I => \eeprom.n4081\
        );

    \I__3556\ : InMux
    port map (
            O => \N__19502\,
            I => \eeprom.n4082\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__3554\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19493\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__19493\,
            I => \eeprom.n2874\
        );

    \I__3552\ : InMux
    port map (
            O => \N__19490\,
            I => \eeprom.n4083\
        );

    \I__3551\ : InMux
    port map (
            O => \N__19487\,
            I => \eeprom.n4084\
        );

    \I__3550\ : InMux
    port map (
            O => \N__19484\,
            I => \N__19481\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__19481\,
            I => \eeprom.n5153\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__19478\,
            I => \N__19475\
        );

    \I__3547\ : InMux
    port map (
            O => \N__19475\,
            I => \N__19470\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__19474\,
            I => \N__19467\
        );

    \I__3545\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19464\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__19470\,
            I => \N__19461\
        );

    \I__3543\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19458\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__19464\,
            I => \N__19455\
        );

    \I__3541\ : Odrv12
    port map (
            O => \N__19461\,
            I => \eeprom.n2918\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__19458\,
            I => \eeprom.n2918\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__19455\,
            I => \eeprom.n2918\
        );

    \I__3538\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19444\
        );

    \I__3537\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19441\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__19444\,
            I => \N__19438\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__19438\,
            I => \N__19429\
        );

    \I__3533\ : Span4Mux_s3_v
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__3532\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19426\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__19429\,
            I => \eeprom.n2911\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__19426\,
            I => \eeprom.n2911\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__19421\,
            I => \N__19418\
        );

    \I__3528\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19415\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__19415\,
            I => \eeprom.n2886\
        );

    \I__3526\ : InMux
    port map (
            O => \N__19412\,
            I => \bfn_21_27_0_\
        );

    \I__3525\ : InMux
    port map (
            O => \N__19409\,
            I => \N__19406\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__19406\,
            I => \eeprom.n2885\
        );

    \I__3523\ : InMux
    port map (
            O => \N__19403\,
            I => \eeprom.n4072\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__19400\,
            I => \N__19397\
        );

    \I__3521\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19394\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__19394\,
            I => \eeprom.n2884\
        );

    \I__3519\ : InMux
    port map (
            O => \N__19391\,
            I => \eeprom.n4073\
        );

    \I__3518\ : InMux
    port map (
            O => \N__19388\,
            I => \N__19385\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__19385\,
            I => \eeprom.n2883\
        );

    \I__3516\ : InMux
    port map (
            O => \N__19382\,
            I => \eeprom.n4074\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__19379\,
            I => \N__19376\
        );

    \I__3514\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19373\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__19373\,
            I => \N__19370\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__19370\,
            I => \eeprom.n2882\
        );

    \I__3511\ : InMux
    port map (
            O => \N__19367\,
            I => \eeprom.n4075\
        );

    \I__3510\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19361\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__19361\,
            I => \eeprom.n2881\
        );

    \I__3508\ : InMux
    port map (
            O => \N__19358\,
            I => \eeprom.n4076\
        );

    \I__3507\ : InMux
    port map (
            O => \N__19355\,
            I => \eeprom.n4055\
        );

    \I__3506\ : InMux
    port map (
            O => \N__19352\,
            I => \eeprom.n4056\
        );

    \I__3505\ : InMux
    port map (
            O => \N__19349\,
            I => \N__19346\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__19346\,
            I => \eeprom.n2677\
        );

    \I__3503\ : InMux
    port map (
            O => \N__19343\,
            I => \N__19340\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__19340\,
            I => \eeprom.n2678\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__19337\,
            I => \eeprom.n2710_cascade_\
        );

    \I__3500\ : InMux
    port map (
            O => \N__19334\,
            I => \N__19331\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__19331\,
            I => \N__19328\
        );

    \I__3498\ : Odrv4
    port map (
            O => \N__19328\,
            I => \eeprom.n2686\
        );

    \I__3497\ : CascadeMux
    port map (
            O => \N__19325\,
            I => \N__19322\
        );

    \I__3496\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19319\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19314\
        );

    \I__3494\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19309\
        );

    \I__3493\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19309\
        );

    \I__3492\ : Span4Mux_v
    port map (
            O => \N__19314\,
            I => \N__19306\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__19309\,
            I => \eeprom.n2912\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__19306\,
            I => \eeprom.n2912\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__19301\,
            I => \eeprom.n5157_cascade_\
        );

    \I__3488\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19295\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__19295\,
            I => \N__19292\
        );

    \I__3486\ : Odrv4
    port map (
            O => \N__19292\,
            I => \eeprom.n16\
        );

    \I__3485\ : InMux
    port map (
            O => \N__19289\,
            I => \eeprom.n4046\
        );

    \I__3484\ : InMux
    port map (
            O => \N__19286\,
            I => \eeprom.n4047\
        );

    \I__3483\ : InMux
    port map (
            O => \N__19283\,
            I => \eeprom.n4048\
        );

    \I__3482\ : InMux
    port map (
            O => \N__19280\,
            I => \eeprom.n4049\
        );

    \I__3481\ : InMux
    port map (
            O => \N__19277\,
            I => \bfn_21_24_0_\
        );

    \I__3480\ : InMux
    port map (
            O => \N__19274\,
            I => \eeprom.n4051\
        );

    \I__3479\ : InMux
    port map (
            O => \N__19271\,
            I => \eeprom.n4052\
        );

    \I__3478\ : InMux
    port map (
            O => \N__19268\,
            I => \eeprom.n4053\
        );

    \I__3477\ : InMux
    port map (
            O => \N__19265\,
            I => \eeprom.n4054\
        );

    \I__3476\ : CascadeMux
    port map (
            O => \N__19262\,
            I => \N__19259\
        );

    \I__3475\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19255\
        );

    \I__3474\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19251\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__19255\,
            I => \N__19248\
        );

    \I__3472\ : InMux
    port map (
            O => \N__19254\,
            I => \N__19245\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__19251\,
            I => \eeprom.n3403\
        );

    \I__3470\ : Odrv4
    port map (
            O => \N__19248\,
            I => \eeprom.n3403\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__19245\,
            I => \eeprom.n3403\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__19238\,
            I => \N__19235\
        );

    \I__3467\ : InMux
    port map (
            O => \N__19235\,
            I => \N__19232\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__19232\,
            I => \N__19229\
        );

    \I__3465\ : Span4Mux_v
    port map (
            O => \N__19229\,
            I => \N__19226\
        );

    \I__3464\ : Odrv4
    port map (
            O => \N__19226\,
            I => \eeprom.n3470\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__19223\,
            I => \N__19216\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__19222\,
            I => \N__19211\
        );

    \I__3461\ : InMux
    port map (
            O => \N__19221\,
            I => \N__19208\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__19220\,
            I => \N__19200\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__19219\,
            I => \N__19197\
        );

    \I__3458\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19191\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__19215\,
            I => \N__19185\
        );

    \I__3456\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19180\
        );

    \I__3455\ : InMux
    port map (
            O => \N__19211\,
            I => \N__19180\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__19208\,
            I => \N__19177\
        );

    \I__3453\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19174\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__19206\,
            I => \N__19169\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__19205\,
            I => \N__19165\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__19204\,
            I => \N__19162\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__19203\,
            I => \N__19158\
        );

    \I__3448\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19151\
        );

    \I__3447\ : InMux
    port map (
            O => \N__19197\,
            I => \N__19151\
        );

    \I__3446\ : InMux
    port map (
            O => \N__19196\,
            I => \N__19151\
        );

    \I__3445\ : InMux
    port map (
            O => \N__19195\,
            I => \N__19146\
        );

    \I__3444\ : InMux
    port map (
            O => \N__19194\,
            I => \N__19146\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__19191\,
            I => \N__19143\
        );

    \I__3442\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19140\
        );

    \I__3441\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19133\
        );

    \I__3440\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19133\
        );

    \I__3439\ : InMux
    port map (
            O => \N__19185\,
            I => \N__19133\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__19180\,
            I => \N__19126\
        );

    \I__3437\ : Span4Mux_v
    port map (
            O => \N__19177\,
            I => \N__19126\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__19174\,
            I => \N__19126\
        );

    \I__3435\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19115\
        );

    \I__3434\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19115\
        );

    \I__3433\ : InMux
    port map (
            O => \N__19169\,
            I => \N__19115\
        );

    \I__3432\ : InMux
    port map (
            O => \N__19168\,
            I => \N__19115\
        );

    \I__3431\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19115\
        );

    \I__3430\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19108\
        );

    \I__3429\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19108\
        );

    \I__3428\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19108\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19101\
        );

    \I__3426\ : LocalMux
    port map (
            O => \N__19146\,
            I => \N__19101\
        );

    \I__3425\ : Span4Mux_h
    port map (
            O => \N__19143\,
            I => \N__19101\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__19140\,
            I => \eeprom.n3430\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__19133\,
            I => \eeprom.n3430\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__19126\,
            I => \eeprom.n3430\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__19115\,
            I => \eeprom.n3430\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__19108\,
            I => \eeprom.n3430\
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__19101\,
            I => \eeprom.n3430\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__19088\,
            I => \N__19085\
        );

    \I__3417\ : InMux
    port map (
            O => \N__19085\,
            I => \N__19081\
        );

    \I__3416\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19078\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__19081\,
            I => \N__19075\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__19078\,
            I => \N__19071\
        );

    \I__3413\ : Span4Mux_h
    port map (
            O => \N__19075\,
            I => \N__19068\
        );

    \I__3412\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19065\
        );

    \I__3411\ : Span4Mux_h
    port map (
            O => \N__19071\,
            I => \N__19062\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__19068\,
            I => \eeprom.n3502\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__19065\,
            I => \eeprom.n3502\
        );

    \I__3408\ : Odrv4
    port map (
            O => \N__19062\,
            I => \eeprom.n3502\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__19055\,
            I => \eeprom.n2511_cascade_\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__19052\,
            I => \eeprom.n2618_cascade_\
        );

    \I__3405\ : InMux
    port map (
            O => \N__19049\,
            I => \bfn_21_23_0_\
        );

    \I__3404\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19043\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__19043\,
            I => \eeprom.n2685\
        );

    \I__3402\ : InMux
    port map (
            O => \N__19040\,
            I => \eeprom.n4043\
        );

    \I__3401\ : InMux
    port map (
            O => \N__19037\,
            I => \eeprom.n4044\
        );

    \I__3400\ : InMux
    port map (
            O => \N__19034\,
            I => \eeprom.n4045\
        );

    \I__3399\ : InMux
    port map (
            O => \N__19031\,
            I => \eeprom.n4009\
        );

    \I__3398\ : InMux
    port map (
            O => \N__19028\,
            I => \eeprom.n4010\
        );

    \I__3397\ : InMux
    port map (
            O => \N__19025\,
            I => \eeprom.n4011\
        );

    \I__3396\ : InMux
    port map (
            O => \N__19022\,
            I => \eeprom.n4012\
        );

    \I__3395\ : InMux
    port map (
            O => \N__19019\,
            I => \eeprom.n4013\
        );

    \I__3394\ : InMux
    port map (
            O => \N__19016\,
            I => \bfn_21_21_0_\
        );

    \I__3393\ : InMux
    port map (
            O => \N__19013\,
            I => \eeprom.n4015\
        );

    \I__3392\ : InMux
    port map (
            O => \N__19010\,
            I => \eeprom.n4016\
        );

    \I__3391\ : InMux
    port map (
            O => \N__19007\,
            I => \eeprom.n4017\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__19004\,
            I => \eeprom.n2214_cascade_\
        );

    \I__3389\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18998\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__18998\,
            I => \N__18995\
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__18995\,
            I => \eeprom.n3720\
        );

    \I__3386\ : InMux
    port map (
            O => \N__18992\,
            I => \bfn_21_20_0_\
        );

    \I__3385\ : InMux
    port map (
            O => \N__18989\,
            I => \eeprom.n4007\
        );

    \I__3384\ : InMux
    port map (
            O => \N__18986\,
            I => \eeprom.n4008\
        );

    \I__3383\ : CascadeMux
    port map (
            O => \N__18983\,
            I => \eeprom.n4847_cascade_\
        );

    \I__3382\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18977\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__18977\,
            I => \eeprom.enable_N_60_5\
        );

    \I__3380\ : InMux
    port map (
            O => \N__18974\,
            I => \N__18971\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__18971\,
            I => \eeprom.enable_N_60_7\
        );

    \I__3378\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18965\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__18965\,
            I => \eeprom.enable_N_60_6\
        );

    \I__3376\ : CascadeMux
    port map (
            O => \N__18962\,
            I => \eeprom.n4853_cascade_\
        );

    \I__3375\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18956\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__18956\,
            I => \eeprom.enable_N_60_8\
        );

    \I__3373\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18950\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__18950\,
            I => \eeprom.enable_N_60_10\
        );

    \I__3371\ : InMux
    port map (
            O => \N__18947\,
            I => \N__18944\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__18944\,
            I => \eeprom.enable_N_60_9\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \eeprom.n4859_cascade_\
        );

    \I__3368\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18935\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__18935\,
            I => \eeprom.enable_N_60_11\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__18932\,
            I => \eeprom.n4865_cascade_\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__18929\,
            I => \eeprom.enable_N_59_cascade_\
        );

    \I__3364\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18920\
        );

    \I__3363\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18920\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__18920\,
            I => \eeprom.enable_N_60_12\
        );

    \I__3361\ : InMux
    port map (
            O => \N__18917\,
            I => \N__18911\
        );

    \I__3360\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18911\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__18911\,
            I => \eeprom.enable_N_60_14\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__18908\,
            I => \N__18905\
        );

    \I__3357\ : InMux
    port map (
            O => \N__18905\,
            I => \N__18901\
        );

    \I__3356\ : InMux
    port map (
            O => \N__18904\,
            I => \N__18898\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__18901\,
            I => \eeprom.enable_N_60_13\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__18898\,
            I => \eeprom.enable_N_60_13\
        );

    \I__3353\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18890\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__18890\,
            I => \eeprom.n4865\
        );

    \I__3351\ : CascadeMux
    port map (
            O => \N__18887\,
            I => \eeprom.n2211_cascade_\
        );

    \I__3350\ : InMux
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__18881\,
            I => \N__18878\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__18878\,
            I => \eeprom.n2975\
        );

    \I__3347\ : InMux
    port map (
            O => \N__18875\,
            I => \eeprom.n4098\
        );

    \I__3346\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18869\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18866\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__18866\,
            I => \eeprom.n2974\
        );

    \I__3343\ : InMux
    port map (
            O => \N__18863\,
            I => \eeprom.n4099\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__18860\,
            I => \N__18857\
        );

    \I__3341\ : InMux
    port map (
            O => \N__18857\,
            I => \N__18853\
        );

    \I__3340\ : InMux
    port map (
            O => \N__18856\,
            I => \N__18850\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__18853\,
            I => \N__18844\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__18850\,
            I => \N__18844\
        );

    \I__3337\ : InMux
    port map (
            O => \N__18849\,
            I => \N__18841\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__18844\,
            I => \eeprom.n2906\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__18841\,
            I => \eeprom.n2906\
        );

    \I__3334\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18833\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18830\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__18830\,
            I => \eeprom.n2973\
        );

    \I__3331\ : InMux
    port map (
            O => \N__18827\,
            I => \eeprom.n4100\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__18824\,
            I => \N__18821\
        );

    \I__3329\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18818\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__18815\,
            I => \eeprom.n2972\
        );

    \I__3326\ : InMux
    port map (
            O => \N__18812\,
            I => \eeprom.n4101\
        );

    \I__3325\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__18806\,
            I => \eeprom.n2971\
        );

    \I__3323\ : InMux
    port map (
            O => \N__18803\,
            I => \eeprom.n4102\
        );

    \I__3322\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18797\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__18797\,
            I => \N__18794\
        );

    \I__3320\ : Span4Mux_v
    port map (
            O => \N__18794\,
            I => \N__18791\
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__18791\,
            I => \eeprom.n2970\
        );

    \I__3318\ : InMux
    port map (
            O => \N__18788\,
            I => \bfn_20_31_0_\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__18785\,
            I => \N__18780\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__18784\,
            I => \N__18771\
        );

    \I__3315\ : CascadeMux
    port map (
            O => \N__18783\,
            I => \N__18767\
        );

    \I__3314\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18764\
        );

    \I__3313\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18761\
        );

    \I__3312\ : CascadeMux
    port map (
            O => \N__18778\,
            I => \N__18757\
        );

    \I__3311\ : CascadeMux
    port map (
            O => \N__18777\,
            I => \N__18754\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__18776\,
            I => \N__18750\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__18775\,
            I => \N__18747\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__18774\,
            I => \N__18742\
        );

    \I__3307\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18733\
        );

    \I__3306\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18733\
        );

    \I__3305\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18733\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__18764\,
            I => \N__18730\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__18761\,
            I => \N__18727\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__18760\,
            I => \N__18724\
        );

    \I__3301\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18714\
        );

    \I__3300\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18714\
        );

    \I__3299\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18714\
        );

    \I__3298\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18714\
        );

    \I__3297\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18707\
        );

    \I__3296\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18707\
        );

    \I__3295\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18707\
        );

    \I__3294\ : InMux
    port map (
            O => \N__18742\,
            I => \N__18700\
        );

    \I__3293\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18700\
        );

    \I__3292\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18700\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__18733\,
            I => \N__18693\
        );

    \I__3290\ : Span4Mux_s2_v
    port map (
            O => \N__18730\,
            I => \N__18693\
        );

    \I__3289\ : Span4Mux_h
    port map (
            O => \N__18727\,
            I => \N__18693\
        );

    \I__3288\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18688\
        );

    \I__3287\ : InMux
    port map (
            O => \N__18723\,
            I => \N__18688\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__18714\,
            I => \eeprom.n2935\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__18707\,
            I => \eeprom.n2935\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__18700\,
            I => \eeprom.n2935\
        );

    \I__3283\ : Odrv4
    port map (
            O => \N__18693\,
            I => \eeprom.n2935\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__18688\,
            I => \eeprom.n2935\
        );

    \I__3281\ : InMux
    port map (
            O => \N__18677\,
            I => \eeprom.n4104\
        );

    \I__3280\ : InMux
    port map (
            O => \N__18674\,
            I => \N__18670\
        );

    \I__3279\ : InMux
    port map (
            O => \N__18673\,
            I => \N__18667\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__18670\,
            I => \N__18664\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18661\
        );

    \I__3276\ : Span4Mux_v
    port map (
            O => \N__18664\,
            I => \N__18658\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__18661\,
            I => \eeprom.n3001\
        );

    \I__3274\ : Odrv4
    port map (
            O => \N__18658\,
            I => \eeprom.n3001\
        );

    \I__3273\ : InMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__18650\,
            I => \eeprom.enable_N_60_0\
        );

    \I__3271\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18644\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__18644\,
            I => \eeprom.enable_N_60_1\
        );

    \I__3269\ : InMux
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__18638\,
            I => \eeprom.enable_N_60_2\
        );

    \I__3267\ : InMux
    port map (
            O => \N__18635\,
            I => \N__18632\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__18629\,
            I => \eeprom.enable_N_60_3\
        );

    \I__3264\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__18623\,
            I => \eeprom.enable_N_60_4\
        );

    \I__3262\ : InMux
    port map (
            O => \N__18620\,
            I => \eeprom.n4090\
        );

    \I__3261\ : CascadeMux
    port map (
            O => \N__18617\,
            I => \N__18613\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__18616\,
            I => \N__18610\
        );

    \I__3259\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18606\
        );

    \I__3258\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18603\
        );

    \I__3257\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18600\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__18606\,
            I => \eeprom.n2915\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__18603\,
            I => \eeprom.n2915\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__18600\,
            I => \eeprom.n2915\
        );

    \I__3253\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__18590\,
            I => \N__18587\
        );

    \I__3251\ : Span4Mux_h
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__18584\,
            I => \eeprom.n2982\
        );

    \I__3249\ : InMux
    port map (
            O => \N__18581\,
            I => \eeprom.n4091\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__3247\ : InMux
    port map (
            O => \N__18575\,
            I => \N__18571\
        );

    \I__3246\ : InMux
    port map (
            O => \N__18574\,
            I => \N__18568\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__18571\,
            I => \N__18565\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__18568\,
            I => \eeprom.n2914\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__18565\,
            I => \eeprom.n2914\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__3241\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__18551\,
            I => \eeprom.n2981\
        );

    \I__3238\ : InMux
    port map (
            O => \N__18548\,
            I => \eeprom.n4092\
        );

    \I__3237\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18541\
        );

    \I__3236\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18538\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__18541\,
            I => \eeprom.n2913\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__18538\,
            I => \eeprom.n2913\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__18533\,
            I => \N__18530\
        );

    \I__3232\ : InMux
    port map (
            O => \N__18530\,
            I => \N__18527\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__18527\,
            I => \N__18524\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__18524\,
            I => \eeprom.n2980\
        );

    \I__3229\ : InMux
    port map (
            O => \N__18521\,
            I => \eeprom.n4093\
        );

    \I__3228\ : InMux
    port map (
            O => \N__18518\,
            I => \N__18515\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__18515\,
            I => \N__18512\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__18512\,
            I => \N__18509\
        );

    \I__3225\ : Odrv4
    port map (
            O => \N__18509\,
            I => \eeprom.n2979\
        );

    \I__3224\ : InMux
    port map (
            O => \N__18506\,
            I => \eeprom.n4094\
        );

    \I__3223\ : InMux
    port map (
            O => \N__18503\,
            I => \N__18500\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__18500\,
            I => \eeprom.n2978\
        );

    \I__3221\ : InMux
    port map (
            O => \N__18497\,
            I => \bfn_20_30_0_\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__18494\,
            I => \N__18490\
        );

    \I__3219\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18487\
        );

    \I__3218\ : InMux
    port map (
            O => \N__18490\,
            I => \N__18484\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__18487\,
            I => \N__18481\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__18484\,
            I => \eeprom.n2910\
        );

    \I__3215\ : Odrv12
    port map (
            O => \N__18481\,
            I => \eeprom.n2910\
        );

    \I__3214\ : InMux
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__18470\,
            I => \N__18467\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__18467\,
            I => \eeprom.n2977\
        );

    \I__3210\ : InMux
    port map (
            O => \N__18464\,
            I => \eeprom.n4096\
        );

    \I__3209\ : InMux
    port map (
            O => \N__18461\,
            I => \N__18456\
        );

    \I__3208\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18453\
        );

    \I__3207\ : InMux
    port map (
            O => \N__18459\,
            I => \N__18450\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__18456\,
            I => \N__18445\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__18453\,
            I => \N__18445\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__18450\,
            I => \eeprom.n2909\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__18445\,
            I => \eeprom.n2909\
        );

    \I__3202\ : InMux
    port map (
            O => \N__18440\,
            I => \N__18437\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__18437\,
            I => \N__18434\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__18434\,
            I => \eeprom.n2976\
        );

    \I__3199\ : InMux
    port map (
            O => \N__18431\,
            I => \eeprom.n4097\
        );

    \I__3198\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18423\
        );

    \I__3197\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18420\
        );

    \I__3196\ : InMux
    port map (
            O => \N__18426\,
            I => \N__18417\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__18423\,
            I => \N__18414\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__18420\,
            I => \eeprom.n2908\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__18417\,
            I => \eeprom.n2908\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__18414\,
            I => \eeprom.n2908\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__18407\,
            I => \eeprom.n2836_cascade_\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__18404\,
            I => \eeprom.n2913_cascade_\
        );

    \I__3189\ : InMux
    port map (
            O => \N__18401\,
            I => \N__18398\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__18398\,
            I => \eeprom.n5297\
        );

    \I__3187\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18392\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__18392\,
            I => \N__18389\
        );

    \I__3185\ : Span4Mux_h
    port map (
            O => \N__18389\,
            I => \N__18386\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__18386\,
            I => \eeprom.n2986\
        );

    \I__3183\ : InMux
    port map (
            O => \N__18383\,
            I => \bfn_20_29_0_\
        );

    \I__3182\ : InMux
    port map (
            O => \N__18380\,
            I => \N__18377\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__18377\,
            I => \N__18374\
        );

    \I__3180\ : Odrv4
    port map (
            O => \N__18374\,
            I => \eeprom.n2985\
        );

    \I__3179\ : InMux
    port map (
            O => \N__18371\,
            I => \eeprom.n4088\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__18368\,
            I => \N__18365\
        );

    \I__3177\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18360\
        );

    \I__3176\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18355\
        );

    \I__3175\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18355\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__18360\,
            I => \eeprom.n2917\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__18355\,
            I => \eeprom.n2917\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__18350\,
            I => \N__18347\
        );

    \I__3171\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18344\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__18344\,
            I => \N__18341\
        );

    \I__3169\ : Odrv4
    port map (
            O => \N__18341\,
            I => \eeprom.n2984\
        );

    \I__3168\ : InMux
    port map (
            O => \N__18338\,
            I => \eeprom.n4089\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__18335\,
            I => \N__18332\
        );

    \I__3166\ : InMux
    port map (
            O => \N__18332\,
            I => \N__18328\
        );

    \I__3165\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18324\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__18328\,
            I => \N__18321\
        );

    \I__3163\ : InMux
    port map (
            O => \N__18327\,
            I => \N__18318\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__18324\,
            I => \eeprom.n2916\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__18321\,
            I => \eeprom.n2916\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__18318\,
            I => \eeprom.n2916\
        );

    \I__3159\ : InMux
    port map (
            O => \N__18311\,
            I => \N__18308\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__18305\,
            I => \eeprom.n2983\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__18302\,
            I => \eeprom.n2910_cascade_\
        );

    \I__3155\ : InMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__18296\,
            I => \eeprom.n15_adj_300\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__18293\,
            I => \eeprom.n22_adj_331_cascade_\
        );

    \I__3152\ : InMux
    port map (
            O => \N__18290\,
            I => \N__18287\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__18287\,
            I => \eeprom.n18_adj_330\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__18284\,
            I => \eeprom.n2935_cascade_\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \N__18278\
        );

    \I__3148\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18274\
        );

    \I__3147\ : InMux
    port map (
            O => \N__18277\,
            I => \N__18271\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N__18263\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__18268\,
            I => \N__18263\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__18263\,
            I => \eeprom.n3015\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__3141\ : InMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__18254\,
            I => \N__18251\
        );

    \I__3139\ : Span4Mux_v
    port map (
            O => \N__18251\,
            I => \N__18247\
        );

    \I__3138\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18244\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__18247\,
            I => \eeprom.n3013\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__18244\,
            I => \eeprom.n3013\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__18239\,
            I => \eeprom.n3015_cascade_\
        );

    \I__3134\ : InMux
    port map (
            O => \N__18236\,
            I => \N__18233\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__18233\,
            I => \eeprom.n5143\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__18230\,
            I => \eeprom.n18_adj_290_cascade_\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__18227\,
            I => \eeprom.n20_adj_291_cascade_\
        );

    \I__3130\ : InMux
    port map (
            O => \N__18224\,
            I => \N__18220\
        );

    \I__3129\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18217\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__18220\,
            I => \N__18213\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18210\
        );

    \I__3126\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18207\
        );

    \I__3125\ : Span4Mux_h
    port map (
            O => \N__18213\,
            I => \N__18204\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__18210\,
            I => \eeprom.n3211\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__18207\,
            I => \eeprom.n3211\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__18204\,
            I => \eeprom.n3211\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__18197\,
            I => \eeprom.n3208_cascade_\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__18194\,
            I => \N__18190\
        );

    \I__3119\ : InMux
    port map (
            O => \N__18193\,
            I => \N__18187\
        );

    \I__3118\ : InMux
    port map (
            O => \N__18190\,
            I => \N__18183\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__18187\,
            I => \N__18180\
        );

    \I__3116\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18177\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__18183\,
            I => \N__18172\
        );

    \I__3114\ : Span4Mux_h
    port map (
            O => \N__18180\,
            I => \N__18172\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__18177\,
            I => \eeprom.n3210\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__18172\,
            I => \eeprom.n3210\
        );

    \I__3111\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18164\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__18164\,
            I => \eeprom.n26_adj_302\
        );

    \I__3109\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18158\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__18158\,
            I => \N__18155\
        );

    \I__3107\ : Span4Mux_h
    port map (
            O => \N__18155\,
            I => \N__18152\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__18152\,
            I => \eeprom.n3080\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__18149\,
            I => \eeprom.n3013_cascade_\
        );

    \I__3104\ : InMux
    port map (
            O => \N__18146\,
            I => \N__18139\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__18145\,
            I => \N__18135\
        );

    \I__3102\ : InMux
    port map (
            O => \N__18144\,
            I => \N__18130\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__18143\,
            I => \N__18125\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__18142\,
            I => \N__18121\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__18139\,
            I => \N__18116\
        );

    \I__3098\ : InMux
    port map (
            O => \N__18138\,
            I => \N__18111\
        );

    \I__3097\ : InMux
    port map (
            O => \N__18135\,
            I => \N__18111\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__18134\,
            I => \N__18105\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__18133\,
            I => \N__18102\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__18130\,
            I => \N__18097\
        );

    \I__3093\ : InMux
    port map (
            O => \N__18129\,
            I => \N__18092\
        );

    \I__3092\ : InMux
    port map (
            O => \N__18128\,
            I => \N__18092\
        );

    \I__3091\ : InMux
    port map (
            O => \N__18125\,
            I => \N__18089\
        );

    \I__3090\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18080\
        );

    \I__3089\ : InMux
    port map (
            O => \N__18121\,
            I => \N__18080\
        );

    \I__3088\ : InMux
    port map (
            O => \N__18120\,
            I => \N__18080\
        );

    \I__3087\ : InMux
    port map (
            O => \N__18119\,
            I => \N__18080\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__18116\,
            I => \N__18075\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__18111\,
            I => \N__18075\
        );

    \I__3084\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18068\
        );

    \I__3083\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18068\
        );

    \I__3082\ : InMux
    port map (
            O => \N__18108\,
            I => \N__18068\
        );

    \I__3081\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18059\
        );

    \I__3080\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18059\
        );

    \I__3079\ : InMux
    port map (
            O => \N__18101\,
            I => \N__18059\
        );

    \I__3078\ : InMux
    port map (
            O => \N__18100\,
            I => \N__18059\
        );

    \I__3077\ : Span4Mux_h
    port map (
            O => \N__18097\,
            I => \N__18056\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__18092\,
            I => \eeprom.n3034\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__18089\,
            I => \eeprom.n3034\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__18080\,
            I => \eeprom.n3034\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__18075\,
            I => \eeprom.n3034\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__18068\,
            I => \eeprom.n3034\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__18059\,
            I => \eeprom.n3034\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__18056\,
            I => \eeprom.n3034\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__18041\,
            I => \N__18038\
        );

    \I__3068\ : InMux
    port map (
            O => \N__18038\,
            I => \N__18035\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__18035\,
            I => \N__18030\
        );

    \I__3066\ : InMux
    port map (
            O => \N__18034\,
            I => \N__18025\
        );

    \I__3065\ : InMux
    port map (
            O => \N__18033\,
            I => \N__18025\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__18030\,
            I => \N__18022\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__18025\,
            I => \eeprom.n3112\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__18022\,
            I => \eeprom.n3112\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__18017\,
            I => \N__18014\
        );

    \I__3060\ : InMux
    port map (
            O => \N__18014\,
            I => \N__18010\
        );

    \I__3059\ : InMux
    port map (
            O => \N__18013\,
            I => \N__18006\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__18010\,
            I => \N__18003\
        );

    \I__3057\ : InMux
    port map (
            O => \N__18009\,
            I => \N__18000\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__18006\,
            I => \N__17995\
        );

    \I__3055\ : Span4Mux_v
    port map (
            O => \N__18003\,
            I => \N__17995\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__18000\,
            I => \eeprom.n3011\
        );

    \I__3053\ : Odrv4
    port map (
            O => \N__17995\,
            I => \eeprom.n3011\
        );

    \I__3052\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17987\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__17987\,
            I => \eeprom.n5301\
        );

    \I__3050\ : InMux
    port map (
            O => \N__17984\,
            I => \N__17980\
        );

    \I__3049\ : InMux
    port map (
            O => \N__17983\,
            I => \N__17976\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__17980\,
            I => \N__17973\
        );

    \I__3047\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17970\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__17976\,
            I => \N__17967\
        );

    \I__3045\ : Span4Mux_s3_v
    port map (
            O => \N__17973\,
            I => \N__17964\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__17970\,
            I => \eeprom.n3110\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__17967\,
            I => \eeprom.n3110\
        );

    \I__3042\ : Odrv4
    port map (
            O => \N__17964\,
            I => \eeprom.n3110\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__17957\,
            I => \N__17949\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__17956\,
            I => \N__17942\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \N__17938\
        );

    \I__3038\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17935\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__17953\,
            I => \N__17930\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__17952\,
            I => \N__17927\
        );

    \I__3035\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17923\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__17948\,
            I => \N__17916\
        );

    \I__3033\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17912\
        );

    \I__3032\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17907\
        );

    \I__3031\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17907\
        );

    \I__3030\ : InMux
    port map (
            O => \N__17942\,
            I => \N__17902\
        );

    \I__3029\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17902\
        );

    \I__3028\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17899\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__17935\,
            I => \N__17896\
        );

    \I__3026\ : InMux
    port map (
            O => \N__17934\,
            I => \N__17885\
        );

    \I__3025\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17885\
        );

    \I__3024\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17885\
        );

    \I__3023\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17885\
        );

    \I__3022\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17885\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__17923\,
            I => \N__17882\
        );

    \I__3020\ : InMux
    port map (
            O => \N__17922\,
            I => \N__17879\
        );

    \I__3019\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17868\
        );

    \I__3018\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17868\
        );

    \I__3017\ : InMux
    port map (
            O => \N__17919\,
            I => \N__17868\
        );

    \I__3016\ : InMux
    port map (
            O => \N__17916\,
            I => \N__17868\
        );

    \I__3015\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17868\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__17912\,
            I => \eeprom.n3133\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__17907\,
            I => \eeprom.n3133\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__17902\,
            I => \eeprom.n3133\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__17899\,
            I => \eeprom.n3133\
        );

    \I__3010\ : Odrv4
    port map (
            O => \N__17896\,
            I => \eeprom.n3133\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__17885\,
            I => \eeprom.n3133\
        );

    \I__3008\ : Odrv12
    port map (
            O => \N__17882\,
            I => \eeprom.n3133\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__17879\,
            I => \eeprom.n3133\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__17868\,
            I => \eeprom.n3133\
        );

    \I__3005\ : InMux
    port map (
            O => \N__17849\,
            I => \N__17846\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__17846\,
            I => \N__17843\
        );

    \I__3003\ : Span4Mux_v
    port map (
            O => \N__17843\,
            I => \N__17840\
        );

    \I__3002\ : Odrv4
    port map (
            O => \N__17840\,
            I => \eeprom.n3177\
        );

    \I__3001\ : InMux
    port map (
            O => \N__17837\,
            I => \N__17833\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__17836\,
            I => \N__17830\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__17833\,
            I => \N__17827\
        );

    \I__2998\ : InMux
    port map (
            O => \N__17830\,
            I => \N__17824\
        );

    \I__2997\ : Span4Mux_h
    port map (
            O => \N__17827\,
            I => \N__17821\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__17824\,
            I => \N__17817\
        );

    \I__2995\ : Span4Mux_h
    port map (
            O => \N__17821\,
            I => \N__17814\
        );

    \I__2994\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17811\
        );

    \I__2993\ : Span4Mux_h
    port map (
            O => \N__17817\,
            I => \N__17808\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__17814\,
            I => \eeprom.n3209\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__17811\,
            I => \eeprom.n3209\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__17808\,
            I => \eeprom.n3209\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__17801\,
            I => \N__17798\
        );

    \I__2988\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17795\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__17789\,
            I => \eeprom.n3283\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__17786\,
            I => \N__17783\
        );

    \I__2983\ : InMux
    port map (
            O => \N__17783\,
            I => \N__17779\
        );

    \I__2982\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17768\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__17779\,
            I => \N__17765\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__17778\,
            I => \N__17759\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__17777\,
            I => \N__17755\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__17776\,
            I => \N__17751\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__17775\,
            I => \N__17748\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__17774\,
            I => \N__17745\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__17773\,
            I => \N__17741\
        );

    \I__2974\ : InMux
    port map (
            O => \N__17772\,
            I => \N__17737\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__17771\,
            I => \N__17732\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__17768\,
            I => \N__17726\
        );

    \I__2971\ : Span4Mux_v
    port map (
            O => \N__17765\,
            I => \N__17726\
        );

    \I__2970\ : InMux
    port map (
            O => \N__17764\,
            I => \N__17721\
        );

    \I__2969\ : InMux
    port map (
            O => \N__17763\,
            I => \N__17721\
        );

    \I__2968\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17716\
        );

    \I__2967\ : InMux
    port map (
            O => \N__17759\,
            I => \N__17716\
        );

    \I__2966\ : InMux
    port map (
            O => \N__17758\,
            I => \N__17709\
        );

    \I__2965\ : InMux
    port map (
            O => \N__17755\,
            I => \N__17709\
        );

    \I__2964\ : InMux
    port map (
            O => \N__17754\,
            I => \N__17709\
        );

    \I__2963\ : InMux
    port map (
            O => \N__17751\,
            I => \N__17700\
        );

    \I__2962\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17700\
        );

    \I__2961\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17700\
        );

    \I__2960\ : InMux
    port map (
            O => \N__17744\,
            I => \N__17700\
        );

    \I__2959\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17695\
        );

    \I__2958\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17695\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__17737\,
            I => \N__17692\
        );

    \I__2956\ : InMux
    port map (
            O => \N__17736\,
            I => \N__17689\
        );

    \I__2955\ : InMux
    port map (
            O => \N__17735\,
            I => \N__17682\
        );

    \I__2954\ : InMux
    port map (
            O => \N__17732\,
            I => \N__17682\
        );

    \I__2953\ : InMux
    port map (
            O => \N__17731\,
            I => \N__17682\
        );

    \I__2952\ : Span4Mux_v
    port map (
            O => \N__17726\,
            I => \N__17679\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__17721\,
            I => \eeprom.n3232\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__17716\,
            I => \eeprom.n3232\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__17709\,
            I => \eeprom.n3232\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__17700\,
            I => \eeprom.n3232\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__17695\,
            I => \eeprom.n3232\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__17692\,
            I => \eeprom.n3232\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__17689\,
            I => \eeprom.n3232\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__17682\,
            I => \eeprom.n3232\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__17679\,
            I => \eeprom.n3232\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__17660\,
            I => \N__17656\
        );

    \I__2941\ : InMux
    port map (
            O => \N__17659\,
            I => \N__17652\
        );

    \I__2940\ : InMux
    port map (
            O => \N__17656\,
            I => \N__17649\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__17655\,
            I => \N__17646\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__17652\,
            I => \N__17643\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__17649\,
            I => \N__17640\
        );

    \I__2936\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17637\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__17643\,
            I => \eeprom.n3315\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__17640\,
            I => \eeprom.n3315\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__17637\,
            I => \eeprom.n3315\
        );

    \I__2932\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17626\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__17629\,
            I => \N__17623\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__17626\,
            I => \N__17620\
        );

    \I__2929\ : InMux
    port map (
            O => \N__17623\,
            I => \N__17617\
        );

    \I__2928\ : Span4Mux_v
    port map (
            O => \N__17620\,
            I => \N__17613\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17610\
        );

    \I__2926\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17607\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__17613\,
            I => \eeprom.n3114\
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__17610\,
            I => \eeprom.n3114\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__17607\,
            I => \eeprom.n3114\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__17600\,
            I => \N__17597\
        );

    \I__2921\ : InMux
    port map (
            O => \N__17597\,
            I => \N__17594\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__17594\,
            I => \N__17591\
        );

    \I__2919\ : Span4Mux_v
    port map (
            O => \N__17591\,
            I => \N__17588\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__17588\,
            I => \eeprom.n3181\
        );

    \I__2917\ : InMux
    port map (
            O => \N__17585\,
            I => \N__17581\
        );

    \I__2916\ : InMux
    port map (
            O => \N__17584\,
            I => \N__17578\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__17581\,
            I => \N__17575\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17572\
        );

    \I__2913\ : Span4Mux_v
    port map (
            O => \N__17575\,
            I => \N__17569\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__17572\,
            I => \N__17566\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__17569\,
            I => \eeprom.n3213\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__17566\,
            I => \eeprom.n3213\
        );

    \I__2909\ : CascadeMux
    port map (
            O => \N__17561\,
            I => \eeprom.n3213_cascade_\
        );

    \I__2908\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17555\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__17555\,
            I => \N__17552\
        );

    \I__2906\ : Span4Mux_v
    port map (
            O => \N__17552\,
            I => \N__17549\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__17549\,
            I => \eeprom.n3182\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__17546\,
            I => \N__17543\
        );

    \I__2903\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17539\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__17542\,
            I => \N__17536\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17533\
        );

    \I__2900\ : InMux
    port map (
            O => \N__17536\,
            I => \N__17530\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__17533\,
            I => \N__17526\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__17530\,
            I => \N__17523\
        );

    \I__2897\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17520\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__17526\,
            I => \eeprom.n3115\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__17523\,
            I => \eeprom.n3115\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__17520\,
            I => \eeprom.n3115\
        );

    \I__2893\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17510\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__17510\,
            I => \N__17506\
        );

    \I__2891\ : InMux
    port map (
            O => \N__17509\,
            I => \N__17503\
        );

    \I__2890\ : Span4Mux_v
    port map (
            O => \N__17506\,
            I => \N__17500\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__17503\,
            I => \eeprom.n3214\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__17500\,
            I => \eeprom.n3214\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__2886\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17488\
        );

    \I__2885\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17485\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__17488\,
            I => \N__17481\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__17485\,
            I => \N__17478\
        );

    \I__2882\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17475\
        );

    \I__2881\ : Span4Mux_h
    port map (
            O => \N__17481\,
            I => \N__17472\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__17478\,
            I => \eeprom.n3216\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__17475\,
            I => \eeprom.n3216\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__17472\,
            I => \eeprom.n3216\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__17465\,
            I => \eeprom.n3214_cascade_\
        );

    \I__2876\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17459\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__17459\,
            I => \eeprom.n5205\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__17456\,
            I => \N__17453\
        );

    \I__2873\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__17450\,
            I => \eeprom.n5209\
        );

    \I__2871\ : InMux
    port map (
            O => \N__17447\,
            I => \N__17443\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__17446\,
            I => \N__17440\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__17443\,
            I => \N__17437\
        );

    \I__2868\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17434\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__17437\,
            I => \N__17430\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__17434\,
            I => \N__17427\
        );

    \I__2865\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17424\
        );

    \I__2864\ : Odrv4
    port map (
            O => \N__17430\,
            I => \eeprom.n3116\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__17427\,
            I => \eeprom.n3116\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__17424\,
            I => \eeprom.n3116\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__17417\,
            I => \N__17414\
        );

    \I__2860\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17411\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__17411\,
            I => \N__17408\
        );

    \I__2858\ : Span4Mux_v
    port map (
            O => \N__17408\,
            I => \N__17405\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__17405\,
            I => \eeprom.n3183\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__17402\,
            I => \N__17399\
        );

    \I__2855\ : InMux
    port map (
            O => \N__17399\,
            I => \N__17395\
        );

    \I__2854\ : InMux
    port map (
            O => \N__17398\,
            I => \N__17392\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__17395\,
            I => \N__17389\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__17392\,
            I => \N__17385\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__17389\,
            I => \N__17382\
        );

    \I__2850\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17379\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__17385\,
            I => \eeprom.n3215\
        );

    \I__2848\ : Odrv4
    port map (
            O => \N__17382\,
            I => \eeprom.n3215\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__17379\,
            I => \eeprom.n3215\
        );

    \I__2846\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17369\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__17369\,
            I => \N__17366\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__17366\,
            I => \N__17363\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__17363\,
            I => \eeprom.n3185\
        );

    \I__2842\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17356\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__17359\,
            I => \N__17353\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17349\
        );

    \I__2839\ : InMux
    port map (
            O => \N__17353\,
            I => \N__17346\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__17352\,
            I => \N__17343\
        );

    \I__2837\ : Span4Mux_v
    port map (
            O => \N__17349\,
            I => \N__17340\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__17346\,
            I => \N__17337\
        );

    \I__2835\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17334\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__17340\,
            I => \eeprom.n3118\
        );

    \I__2833\ : Odrv12
    port map (
            O => \N__17337\,
            I => \eeprom.n3118\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__17334\,
            I => \eeprom.n3118\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__17327\,
            I => \N__17324\
        );

    \I__2830\ : InMux
    port map (
            O => \N__17324\,
            I => \N__17321\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__17321\,
            I => \N__17316\
        );

    \I__2828\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17313\
        );

    \I__2827\ : InMux
    port map (
            O => \N__17319\,
            I => \N__17310\
        );

    \I__2826\ : Span4Mux_h
    port map (
            O => \N__17316\,
            I => \N__17307\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__17313\,
            I => \eeprom.n3217\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__17310\,
            I => \eeprom.n3217\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__17307\,
            I => \eeprom.n3217\
        );

    \I__2822\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17296\
        );

    \I__2821\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17293\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__17296\,
            I => \N__17289\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__17293\,
            I => \N__17286\
        );

    \I__2818\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17283\
        );

    \I__2817\ : Span4Mux_h
    port map (
            O => \N__17289\,
            I => \N__17280\
        );

    \I__2816\ : Span4Mux_s2_v
    port map (
            O => \N__17286\,
            I => \N__17277\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__17283\,
            I => \N__17274\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__17280\,
            I => \eeprom.n3109\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__17277\,
            I => \eeprom.n3109\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__17274\,
            I => \eeprom.n3109\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__17267\,
            I => \N__17264\
        );

    \I__2810\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17261\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__17261\,
            I => \N__17258\
        );

    \I__2808\ : Span4Mux_v
    port map (
            O => \N__17258\,
            I => \N__17255\
        );

    \I__2807\ : Odrv4
    port map (
            O => \N__17255\,
            I => \eeprom.n3176\
        );

    \I__2806\ : InMux
    port map (
            O => \N__17252\,
            I => \N__17248\
        );

    \I__2805\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17245\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__17248\,
            I => \N__17242\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17239\
        );

    \I__2802\ : Span4Mux_h
    port map (
            O => \N__17242\,
            I => \N__17234\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__17239\,
            I => \N__17234\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__17234\,
            I => \eeprom.n3208\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__17231\,
            I => \eeprom.n3413_cascade_\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__17228\,
            I => \N__17224\
        );

    \I__2797\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17221\
        );

    \I__2796\ : InMux
    port map (
            O => \N__17224\,
            I => \N__17218\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__17221\,
            I => \N__17212\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__17218\,
            I => \N__17212\
        );

    \I__2793\ : InMux
    port map (
            O => \N__17217\,
            I => \N__17209\
        );

    \I__2792\ : Span4Mux_h
    port map (
            O => \N__17212\,
            I => \N__17206\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__17209\,
            I => \eeprom.n3415\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__17206\,
            I => \eeprom.n3415\
        );

    \I__2789\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17198\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__17198\,
            I => \eeprom.n5289\
        );

    \I__2787\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__2784\ : Span4Mux_h
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__17183\,
            I => \eeprom.n3278\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__17180\,
            I => \N__17177\
        );

    \I__2781\ : InMux
    port map (
            O => \N__17177\,
            I => \N__17174\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__17174\,
            I => \N__17171\
        );

    \I__2779\ : Span4Mux_h
    port map (
            O => \N__17171\,
            I => \N__17167\
        );

    \I__2778\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17164\
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__17167\,
            I => \eeprom.n3310\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__17164\,
            I => \eeprom.n3310\
        );

    \I__2775\ : InMux
    port map (
            O => \N__17159\,
            I => \N__17152\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__17158\,
            I => \N__17142\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__17157\,
            I => \N__17137\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__17156\,
            I => \N__17133\
        );

    \I__2771\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17129\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__17152\,
            I => \N__17126\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__17151\,
            I => \N__17120\
        );

    \I__2768\ : CascadeMux
    port map (
            O => \N__17150\,
            I => \N__17116\
        );

    \I__2767\ : InMux
    port map (
            O => \N__17149\,
            I => \N__17112\
        );

    \I__2766\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17107\
        );

    \I__2765\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17107\
        );

    \I__2764\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17096\
        );

    \I__2763\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17096\
        );

    \I__2762\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17096\
        );

    \I__2761\ : InMux
    port map (
            O => \N__17141\,
            I => \N__17096\
        );

    \I__2760\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17096\
        );

    \I__2759\ : InMux
    port map (
            O => \N__17137\,
            I => \N__17087\
        );

    \I__2758\ : InMux
    port map (
            O => \N__17136\,
            I => \N__17087\
        );

    \I__2757\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17087\
        );

    \I__2756\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17087\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__17129\,
            I => \N__17084\
        );

    \I__2754\ : Span4Mux_h
    port map (
            O => \N__17126\,
            I => \N__17081\
        );

    \I__2753\ : InMux
    port map (
            O => \N__17125\,
            I => \N__17074\
        );

    \I__2752\ : InMux
    port map (
            O => \N__17124\,
            I => \N__17074\
        );

    \I__2751\ : InMux
    port map (
            O => \N__17123\,
            I => \N__17074\
        );

    \I__2750\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17065\
        );

    \I__2749\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17065\
        );

    \I__2748\ : InMux
    port map (
            O => \N__17116\,
            I => \N__17065\
        );

    \I__2747\ : InMux
    port map (
            O => \N__17115\,
            I => \N__17065\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__17112\,
            I => \eeprom.n3331\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__17107\,
            I => \eeprom.n3331\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__17096\,
            I => \eeprom.n3331\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__17087\,
            I => \eeprom.n3331\
        );

    \I__2742\ : Odrv4
    port map (
            O => \N__17084\,
            I => \eeprom.n3331\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__17081\,
            I => \eeprom.n3331\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__17074\,
            I => \eeprom.n3331\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__17065\,
            I => \eeprom.n3331\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__17048\,
            I => \eeprom.n3310_cascade_\
        );

    \I__2737\ : InMux
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__17042\,
            I => \N__17039\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__17036\,
            I => \eeprom.n3377\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__17033\,
            I => \N__17030\
        );

    \I__2732\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17026\
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__17029\,
            I => \N__17023\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__17026\,
            I => \N__17019\
        );

    \I__2729\ : InMux
    port map (
            O => \N__17023\,
            I => \N__17014\
        );

    \I__2728\ : InMux
    port map (
            O => \N__17022\,
            I => \N__17014\
        );

    \I__2727\ : Span4Mux_h
    port map (
            O => \N__17019\,
            I => \N__17011\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__17014\,
            I => \eeprom.n3409\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__17011\,
            I => \eeprom.n3409\
        );

    \I__2724\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17003\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__17000\,
            I => \N__16997\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__16997\,
            I => \eeprom.n3284\
        );

    \I__2720\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__16991\,
            I => \N__16986\
        );

    \I__2718\ : InMux
    port map (
            O => \N__16990\,
            I => \N__16983\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__16989\,
            I => \N__16980\
        );

    \I__2716\ : Span4Mux_v
    port map (
            O => \N__16986\,
            I => \N__16977\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__16983\,
            I => \N__16974\
        );

    \I__2714\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16971\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__16977\,
            I => \eeprom.n3218\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__16974\,
            I => \eeprom.n3218\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__16971\,
            I => \eeprom.n3218\
        );

    \I__2710\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16961\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__16961\,
            I => \N__16958\
        );

    \I__2708\ : Span4Mux_h
    port map (
            O => \N__16958\,
            I => \N__16955\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__16955\,
            I => \eeprom.n3285\
        );

    \I__2706\ : InMux
    port map (
            O => \N__16952\,
            I => \N__16948\
        );

    \I__2705\ : InMux
    port map (
            O => \N__16951\,
            I => \N__16945\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__16948\,
            I => \N__16942\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__16945\,
            I => \N__16939\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__16942\,
            I => \eeprom.n3317\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__16939\,
            I => \eeprom.n3317\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__2699\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__16928\,
            I => \N__16925\
        );

    \I__2697\ : Span4Mux_h
    port map (
            O => \N__16925\,
            I => \N__16921\
        );

    \I__2696\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16918\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__16921\,
            I => \eeprom.n3314\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__16918\,
            I => \eeprom.n3314\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__16913\,
            I => \eeprom.n3317_cascade_\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__16910\,
            I => \N__16907\
        );

    \I__2691\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16902\
        );

    \I__2690\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16899\
        );

    \I__2689\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16896\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__16902\,
            I => \N__16893\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__16899\,
            I => \N__16890\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__16896\,
            I => \N__16885\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__16893\,
            I => \N__16885\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__16890\,
            I => \eeprom.n3316\
        );

    \I__2683\ : Odrv4
    port map (
            O => \N__16885\,
            I => \eeprom.n3316\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__16880\,
            I => \N__16875\
        );

    \I__2681\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16872\
        );

    \I__2680\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16869\
        );

    \I__2679\ : InMux
    port map (
            O => \N__16875\,
            I => \N__16866\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__16872\,
            I => \N__16863\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__16869\,
            I => \eeprom.n3318\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__16866\,
            I => \eeprom.n3318\
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__16863\,
            I => \eeprom.n3318\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__16856\,
            I => \eeprom.n5315_cascade_\
        );

    \I__2673\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16850\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__16850\,
            I => \eeprom.n5313\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__16847\,
            I => \N__16844\
        );

    \I__2670\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16841\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__16841\,
            I => \N__16837\
        );

    \I__2668\ : InMux
    port map (
            O => \N__16840\,
            I => \N__16833\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__16837\,
            I => \N__16830\
        );

    \I__2666\ : InMux
    port map (
            O => \N__16836\,
            I => \N__16827\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__16833\,
            I => \eeprom.n3303\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__16830\,
            I => \eeprom.n3303\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__16827\,
            I => \eeprom.n3303\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__16820\,
            I => \N__16816\
        );

    \I__2661\ : InMux
    port map (
            O => \N__16819\,
            I => \N__16813\
        );

    \I__2660\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16810\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__16813\,
            I => \N__16806\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__16810\,
            I => \N__16803\
        );

    \I__2657\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16800\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__16806\,
            I => \eeprom.n3304\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__16803\,
            I => \eeprom.n3304\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__16800\,
            I => \eeprom.n3304\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__16793\,
            I => \eeprom.n4820_cascade_\
        );

    \I__2652\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16786\
        );

    \I__2651\ : InMux
    port map (
            O => \N__16789\,
            I => \N__16782\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__16786\,
            I => \N__16779\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__16785\,
            I => \N__16776\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__16782\,
            I => \N__16773\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__16779\,
            I => \N__16770\
        );

    \I__2646\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16767\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__16773\,
            I => \N__16764\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__16770\,
            I => \eeprom.n3302\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__16767\,
            I => \eeprom.n3302\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__16764\,
            I => \eeprom.n3302\
        );

    \I__2641\ : InMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__16754\,
            I => \eeprom.n26\
        );

    \I__2639\ : CascadeMux
    port map (
            O => \N__16751\,
            I => \N__16747\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__16750\,
            I => \N__16744\
        );

    \I__2637\ : InMux
    port map (
            O => \N__16747\,
            I => \N__16741\
        );

    \I__2636\ : InMux
    port map (
            O => \N__16744\,
            I => \N__16738\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__16741\,
            I => \N__16734\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__16738\,
            I => \N__16731\
        );

    \I__2633\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16728\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__16734\,
            I => \N__16725\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__16731\,
            I => \eeprom.n3405\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__16728\,
            I => \eeprom.n3405\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__16725\,
            I => \eeprom.n3405\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__16718\,
            I => \eeprom.n4824_cascade_\
        );

    \I__2627\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16711\
        );

    \I__2626\ : InMux
    port map (
            O => \N__16714\,
            I => \N__16707\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__16711\,
            I => \N__16704\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__16710\,
            I => \N__16701\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__16707\,
            I => \N__16698\
        );

    \I__2622\ : Span4Mux_v
    port map (
            O => \N__16704\,
            I => \N__16695\
        );

    \I__2621\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16692\
        );

    \I__2620\ : Span4Mux_h
    port map (
            O => \N__16698\,
            I => \N__16689\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__16695\,
            I => \eeprom.n3404\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__16692\,
            I => \eeprom.n3404\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__16689\,
            I => \eeprom.n3404\
        );

    \I__2616\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16679\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__16679\,
            I => \eeprom.n28_adj_261\
        );

    \I__2614\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__2612\ : Span4Mux_h
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__16667\,
            I => \eeprom.n3386\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__2609\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__16658\,
            I => \N__16653\
        );

    \I__2607\ : InMux
    port map (
            O => \N__16657\,
            I => \N__16650\
        );

    \I__2606\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16647\
        );

    \I__2605\ : Span4Mux_h
    port map (
            O => \N__16653\,
            I => \N__16644\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__16650\,
            I => \eeprom.n3418\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__16647\,
            I => \eeprom.n3418\
        );

    \I__2602\ : Odrv4
    port map (
            O => \N__16644\,
            I => \eeprom.n3418\
        );

    \I__2601\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16634\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__16634\,
            I => \N__16631\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__16631\,
            I => \N__16628\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__16628\,
            I => \eeprom.n3384\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__16625\,
            I => \N__16622\
        );

    \I__2596\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__16619\,
            I => \N__16614\
        );

    \I__2594\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16611\
        );

    \I__2593\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16608\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__16614\,
            I => \N__16605\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__16611\,
            I => \eeprom.n3416\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__16608\,
            I => \eeprom.n3416\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__16605\,
            I => \eeprom.n3416\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__2587\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__2585\ : Span4Mux_v
    port map (
            O => \N__16589\,
            I => \N__16586\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__16586\,
            I => \eeprom.n3383\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__16583\,
            I => \N__16579\
        );

    \I__2582\ : InMux
    port map (
            O => \N__16582\,
            I => \N__16576\
        );

    \I__2581\ : InMux
    port map (
            O => \N__16579\,
            I => \N__16573\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__16576\,
            I => \N__16569\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__16573\,
            I => \N__16566\
        );

    \I__2578\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16563\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__16569\,
            I => \eeprom.n3313\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__16566\,
            I => \eeprom.n3313\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__16563\,
            I => \eeprom.n3313\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__16556\,
            I => \N__16553\
        );

    \I__2573\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16550\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__16550\,
            I => \N__16547\
        );

    \I__2571\ : Span4Mux_h
    port map (
            O => \N__16547\,
            I => \N__16544\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__16544\,
            I => \eeprom.n3371\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__16541\,
            I => \N__16538\
        );

    \I__2568\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__16532\,
            I => \N__16529\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__16529\,
            I => \eeprom.n3282\
        );

    \I__2564\ : InMux
    port map (
            O => \N__16526\,
            I => \N__16523\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__16517\,
            I => \eeprom.n3381\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__16514\,
            I => \eeprom.n3314_cascade_\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__16511\,
            I => \N__16507\
        );

    \I__2558\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16504\
        );

    \I__2557\ : InMux
    port map (
            O => \N__16507\,
            I => \N__16501\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__16504\,
            I => \N__16496\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__16501\,
            I => \N__16496\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__16496\,
            I => \N__16493\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__16493\,
            I => \eeprom.n3413\
        );

    \I__2552\ : InMux
    port map (
            O => \N__16490\,
            I => \eeprom.n4222\
        );

    \I__2551\ : CascadeMux
    port map (
            O => \N__16487\,
            I => \N__16482\
        );

    \I__2550\ : InMux
    port map (
            O => \N__16486\,
            I => \N__16479\
        );

    \I__2549\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16476\
        );

    \I__2548\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16473\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__16479\,
            I => \eeprom.n3500\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__16476\,
            I => \eeprom.n3500\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__16473\,
            I => \eeprom.n3500\
        );

    \I__2544\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__16460\,
            I => \eeprom.n3567\
        );

    \I__2541\ : InMux
    port map (
            O => \N__16457\,
            I => \eeprom.n4223\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__16454\,
            I => \N__16450\
        );

    \I__2539\ : InMux
    port map (
            O => \N__16453\,
            I => \N__16446\
        );

    \I__2538\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16443\
        );

    \I__2537\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16440\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__16446\,
            I => \eeprom.n3499\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__16443\,
            I => \eeprom.n3499\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__16440\,
            I => \eeprom.n3499\
        );

    \I__2533\ : InMux
    port map (
            O => \N__16433\,
            I => \N__16430\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__16430\,
            I => \eeprom.n3566\
        );

    \I__2531\ : InMux
    port map (
            O => \N__16427\,
            I => \eeprom.n4224\
        );

    \I__2530\ : InMux
    port map (
            O => \N__16424\,
            I => \N__16421\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__16421\,
            I => \N__16417\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__16420\,
            I => \N__16414\
        );

    \I__2527\ : Span4Mux_h
    port map (
            O => \N__16417\,
            I => \N__16411\
        );

    \I__2526\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16408\
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__16411\,
            I => \eeprom.n3498\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__16408\,
            I => \eeprom.n3498\
        );

    \I__2523\ : InMux
    port map (
            O => \N__16403\,
            I => \N__16400\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__16400\,
            I => \N__16397\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__16397\,
            I => \eeprom.n3565\
        );

    \I__2520\ : InMux
    port map (
            O => \N__16394\,
            I => \eeprom.n4225\
        );

    \I__2519\ : InMux
    port map (
            O => \N__16391\,
            I => \N__16387\
        );

    \I__2518\ : InMux
    port map (
            O => \N__16390\,
            I => \N__16384\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__16387\,
            I => \N__16381\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__16384\,
            I => \N__16377\
        );

    \I__2515\ : Span4Mux_h
    port map (
            O => \N__16381\,
            I => \N__16374\
        );

    \I__2514\ : InMux
    port map (
            O => \N__16380\,
            I => \N__16371\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__16377\,
            I => \eeprom.n3497\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__16374\,
            I => \eeprom.n3497\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__16371\,
            I => \eeprom.n3497\
        );

    \I__2510\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16361\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__16361\,
            I => \eeprom.n3564\
        );

    \I__2508\ : InMux
    port map (
            O => \N__16358\,
            I => \eeprom.n4226\
        );

    \I__2507\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__16352\,
            I => \N__16348\
        );

    \I__2505\ : InMux
    port map (
            O => \N__16351\,
            I => \N__16345\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__16348\,
            I => \N__16340\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__16345\,
            I => \N__16340\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__16340\,
            I => \N__16337\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__16337\,
            I => \eeprom.n3496\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__16334\,
            I => \N__16331\
        );

    \I__2499\ : InMux
    port map (
            O => \N__16331\,
            I => \N__16325\
        );

    \I__2498\ : InMux
    port map (
            O => \N__16330\,
            I => \N__16314\
        );

    \I__2497\ : InMux
    port map (
            O => \N__16329\,
            I => \N__16314\
        );

    \I__2496\ : InMux
    port map (
            O => \N__16328\,
            I => \N__16311\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__16325\,
            I => \N__16308\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__16324\,
            I => \N__16305\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__16323\,
            I => \N__16302\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__16322\,
            I => \N__16294\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__16321\,
            I => \N__16291\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__16320\,
            I => \N__16286\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__16319\,
            I => \N__16280\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__16314\,
            I => \N__16274\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__16311\,
            I => \N__16269\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__16308\,
            I => \N__16269\
        );

    \I__2485\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16260\
        );

    \I__2484\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16260\
        );

    \I__2483\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16260\
        );

    \I__2482\ : InMux
    port map (
            O => \N__16300\,
            I => \N__16260\
        );

    \I__2481\ : InMux
    port map (
            O => \N__16299\,
            I => \N__16247\
        );

    \I__2480\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16247\
        );

    \I__2479\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16247\
        );

    \I__2478\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16247\
        );

    \I__2477\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16247\
        );

    \I__2476\ : InMux
    port map (
            O => \N__16290\,
            I => \N__16247\
        );

    \I__2475\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16236\
        );

    \I__2474\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16236\
        );

    \I__2473\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16236\
        );

    \I__2472\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16236\
        );

    \I__2471\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16236\
        );

    \I__2470\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16227\
        );

    \I__2469\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16227\
        );

    \I__2468\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16227\
        );

    \I__2467\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16227\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__16274\,
            I => \eeprom.n3529\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__16269\,
            I => \eeprom.n3529\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__16260\,
            I => \eeprom.n3529\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__16247\,
            I => \eeprom.n3529\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__16236\,
            I => \eeprom.n3529\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__16227\,
            I => \eeprom.n3529\
        );

    \I__2460\ : InMux
    port map (
            O => \N__16214\,
            I => \eeprom.n4227\
        );

    \I__2459\ : InMux
    port map (
            O => \N__16211\,
            I => \N__16208\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__16208\,
            I => \N__16205\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__16205\,
            I => \N__16202\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__16202\,
            I => \eeprom.n5355\
        );

    \I__2455\ : InMux
    port map (
            O => \N__16199\,
            I => \N__16196\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__16190\,
            I => \eeprom.n3382\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__2450\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16180\
        );

    \I__2449\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16177\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__16180\,
            I => \N__16172\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__16177\,
            I => \N__16172\
        );

    \I__2446\ : Span4Mux_v
    port map (
            O => \N__16172\,
            I => \N__16169\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__16169\,
            I => \eeprom.n3414\
        );

    \I__2444\ : CascadeMux
    port map (
            O => \N__16166\,
            I => \N__16162\
        );

    \I__2443\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16159\
        );

    \I__2442\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16156\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__16159\,
            I => \N__16152\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__16156\,
            I => \N__16149\
        );

    \I__2439\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16146\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__16152\,
            I => \N__16141\
        );

    \I__2437\ : Span4Mux_h
    port map (
            O => \N__16149\,
            I => \N__16141\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__16146\,
            I => \eeprom.n3417\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__16141\,
            I => \eeprom.n3417\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__16136\,
            I => \eeprom.n3414_cascade_\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__16133\,
            I => \eeprom.n5291_cascade_\
        );

    \I__2432\ : InMux
    port map (
            O => \N__16130\,
            I => \N__16125\
        );

    \I__2431\ : InMux
    port map (
            O => \N__16129\,
            I => \N__16122\
        );

    \I__2430\ : InMux
    port map (
            O => \N__16128\,
            I => \N__16119\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__16125\,
            I => \N__16116\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16113\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__16119\,
            I => \N__16110\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__16116\,
            I => \N__16105\
        );

    \I__2425\ : Span4Mux_h
    port map (
            O => \N__16113\,
            I => \N__16105\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__16110\,
            I => \eeprom.n3508\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__16105\,
            I => \eeprom.n3508\
        );

    \I__2422\ : InMux
    port map (
            O => \N__16100\,
            I => \N__16097\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__16097\,
            I => \eeprom.n3575\
        );

    \I__2420\ : InMux
    port map (
            O => \N__16094\,
            I => \eeprom.n4215\
        );

    \I__2419\ : InMux
    port map (
            O => \N__16091\,
            I => \N__16087\
        );

    \I__2418\ : InMux
    port map (
            O => \N__16090\,
            I => \N__16084\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__16087\,
            I => \N__16079\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__16084\,
            I => \N__16079\
        );

    \I__2415\ : Span4Mux_h
    port map (
            O => \N__16079\,
            I => \N__16076\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__16076\,
            I => \eeprom.n3507\
        );

    \I__2413\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16070\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__16070\,
            I => \eeprom.n3574\
        );

    \I__2411\ : InMux
    port map (
            O => \N__16067\,
            I => \eeprom.n4216\
        );

    \I__2410\ : InMux
    port map (
            O => \N__16064\,
            I => \N__16059\
        );

    \I__2409\ : InMux
    port map (
            O => \N__16063\,
            I => \N__16056\
        );

    \I__2408\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16053\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__16059\,
            I => \eeprom.n3506\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__16056\,
            I => \eeprom.n3506\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__16053\,
            I => \eeprom.n3506\
        );

    \I__2404\ : InMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__16043\,
            I => \N__16040\
        );

    \I__2402\ : Span4Mux_h
    port map (
            O => \N__16040\,
            I => \N__16037\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__16037\,
            I => \eeprom.n3573\
        );

    \I__2400\ : InMux
    port map (
            O => \N__16034\,
            I => \eeprom.n4217\
        );

    \I__2399\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16027\
        );

    \I__2398\ : InMux
    port map (
            O => \N__16030\,
            I => \N__16024\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__16027\,
            I => \N__16021\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__16024\,
            I => \N__16018\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__16021\,
            I => \eeprom.n3505\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__16018\,
            I => \eeprom.n3505\
        );

    \I__2393\ : InMux
    port map (
            O => \N__16013\,
            I => \N__16010\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__16010\,
            I => \eeprom.n3572\
        );

    \I__2391\ : InMux
    port map (
            O => \N__16007\,
            I => \eeprom.n4218\
        );

    \I__2390\ : InMux
    port map (
            O => \N__16004\,
            I => \N__16000\
        );

    \I__2389\ : InMux
    port map (
            O => \N__16003\,
            I => \N__15997\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__16000\,
            I => \N__15994\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__15997\,
            I => \N__15990\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__15994\,
            I => \N__15987\
        );

    \I__2385\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15984\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__15990\,
            I => \eeprom.n3504\
        );

    \I__2383\ : Odrv4
    port map (
            O => \N__15987\,
            I => \eeprom.n3504\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__15984\,
            I => \eeprom.n3504\
        );

    \I__2381\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15974\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__15974\,
            I => \eeprom.n3571\
        );

    \I__2379\ : InMux
    port map (
            O => \N__15971\,
            I => \eeprom.n4219\
        );

    \I__2378\ : InMux
    port map (
            O => \N__15968\,
            I => \N__15965\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__15965\,
            I => \N__15962\
        );

    \I__2376\ : Span4Mux_h
    port map (
            O => \N__15962\,
            I => \N__15957\
        );

    \I__2375\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15952\
        );

    \I__2374\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15952\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__15957\,
            I => \eeprom.n3503\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__15952\,
            I => \eeprom.n3503\
        );

    \I__2371\ : InMux
    port map (
            O => \N__15947\,
            I => \N__15944\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__15944\,
            I => \N__15941\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__15941\,
            I => \eeprom.n3570\
        );

    \I__2368\ : InMux
    port map (
            O => \N__15938\,
            I => \bfn_20_21_0_\
        );

    \I__2367\ : InMux
    port map (
            O => \N__15935\,
            I => \N__15932\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__15932\,
            I => \N__15929\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__15929\,
            I => \N__15926\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__15926\,
            I => \eeprom.n3569\
        );

    \I__2363\ : InMux
    port map (
            O => \N__15923\,
            I => \eeprom.n4221\
        );

    \I__2362\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15917\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__15917\,
            I => \N__15912\
        );

    \I__2360\ : InMux
    port map (
            O => \N__15916\,
            I => \N__15909\
        );

    \I__2359\ : InMux
    port map (
            O => \N__15915\,
            I => \N__15906\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__15912\,
            I => \N__15901\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__15909\,
            I => \N__15901\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__15906\,
            I => \N__15898\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__15901\,
            I => \eeprom.n3501\
        );

    \I__2354\ : Odrv12
    port map (
            O => \N__15898\,
            I => \eeprom.n3501\
        );

    \I__2353\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15890\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__15890\,
            I => \N__15887\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__15887\,
            I => \eeprom.n3568\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__15884\,
            I => \N__15881\
        );

    \I__2349\ : InMux
    port map (
            O => \N__15881\,
            I => \N__15877\
        );

    \I__2348\ : InMux
    port map (
            O => \N__15880\,
            I => \N__15874\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__15877\,
            I => \N__15871\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__15874\,
            I => \N__15867\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__15871\,
            I => \N__15864\
        );

    \I__2344\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15861\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__15867\,
            I => \eeprom.n3516\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__15864\,
            I => \eeprom.n3516\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__15861\,
            I => \eeprom.n3516\
        );

    \I__2340\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15851\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__15851\,
            I => \N__15848\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__15848\,
            I => \eeprom.n3583\
        );

    \I__2337\ : InMux
    port map (
            O => \N__15845\,
            I => \eeprom.n4207\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__15842\,
            I => \N__15838\
        );

    \I__2335\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15835\
        );

    \I__2334\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15832\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__15835\,
            I => \N__15828\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__15832\,
            I => \N__15825\
        );

    \I__2331\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15822\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__15828\,
            I => \eeprom.n3515\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__15825\,
            I => \eeprom.n3515\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__15822\,
            I => \eeprom.n3515\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__15815\,
            I => \N__15812\
        );

    \I__2326\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15809\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__15809\,
            I => \N__15806\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__15806\,
            I => \eeprom.n3582\
        );

    \I__2323\ : InMux
    port map (
            O => \N__15803\,
            I => \eeprom.n4208\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__15800\,
            I => \N__15797\
        );

    \I__2321\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15794\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__15794\,
            I => \N__15790\
        );

    \I__2319\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15787\
        );

    \I__2318\ : Span4Mux_h
    port map (
            O => \N__15790\,
            I => \N__15784\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__15787\,
            I => \eeprom.n3514\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__15784\,
            I => \eeprom.n3514\
        );

    \I__2315\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15776\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__2313\ : Span4Mux_v
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__15770\,
            I => \eeprom.n3581_adj_292\
        );

    \I__2311\ : InMux
    port map (
            O => \N__15767\,
            I => \eeprom.n4209\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__15764\,
            I => \N__15761\
        );

    \I__2309\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__15758\,
            I => \N__15754\
        );

    \I__2307\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15751\
        );

    \I__2306\ : Span4Mux_h
    port map (
            O => \N__15754\,
            I => \N__15748\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__15751\,
            I => \eeprom.n3513\
        );

    \I__2304\ : Odrv4
    port map (
            O => \N__15748\,
            I => \eeprom.n3513\
        );

    \I__2303\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15740\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__15737\,
            I => \eeprom.n3580\
        );

    \I__2300\ : InMux
    port map (
            O => \N__15734\,
            I => \eeprom.n4210\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__15731\,
            I => \N__15728\
        );

    \I__2298\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15724\
        );

    \I__2297\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15721\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__15724\,
            I => \N__15718\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__15721\,
            I => \eeprom.n3512\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__15718\,
            I => \eeprom.n3512\
        );

    \I__2293\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15710\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__15710\,
            I => \N__15707\
        );

    \I__2291\ : Span4Mux_h
    port map (
            O => \N__15707\,
            I => \N__15704\
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__15704\,
            I => \eeprom.n3579\
        );

    \I__2289\ : InMux
    port map (
            O => \N__15701\,
            I => \eeprom.n4211\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__2287\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__15692\,
            I => \N__15687\
        );

    \I__2285\ : InMux
    port map (
            O => \N__15691\,
            I => \N__15684\
        );

    \I__2284\ : InMux
    port map (
            O => \N__15690\,
            I => \N__15681\
        );

    \I__2283\ : Span4Mux_v
    port map (
            O => \N__15687\,
            I => \N__15678\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__15684\,
            I => \eeprom.n3511\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__15681\,
            I => \eeprom.n3511\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__15678\,
            I => \eeprom.n3511\
        );

    \I__2279\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15668\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__15668\,
            I => \eeprom.n3578\
        );

    \I__2277\ : InMux
    port map (
            O => \N__15665\,
            I => \bfn_20_20_0_\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__15662\,
            I => \N__15659\
        );

    \I__2275\ : InMux
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__15656\,
            I => \N__15651\
        );

    \I__2273\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15648\
        );

    \I__2272\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15645\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__15651\,
            I => \N__15642\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__15648\,
            I => \eeprom.n3510\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__15645\,
            I => \eeprom.n3510\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__15642\,
            I => \eeprom.n3510\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__15635\,
            I => \N__15632\
        );

    \I__2266\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15629\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__15629\,
            I => \eeprom.n3577\
        );

    \I__2264\ : InMux
    port map (
            O => \N__15626\,
            I => \eeprom.n4213\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__2262\ : InMux
    port map (
            O => \N__15620\,
            I => \N__15616\
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__15616\,
            I => \N__15610\
        );

    \I__2259\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15606\
        );

    \I__2258\ : Span4Mux_h
    port map (
            O => \N__15610\,
            I => \N__15603\
        );

    \I__2257\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15600\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__15606\,
            I => \eeprom.n3509\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__15603\,
            I => \eeprom.n3509\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__15600\,
            I => \eeprom.n3509\
        );

    \I__2253\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15590\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__15590\,
            I => \eeprom.n3576\
        );

    \I__2251\ : InMux
    port map (
            O => \N__15587\,
            I => \eeprom.n4214\
        );

    \I__2250\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15581\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__15581\,
            I => \eeprom.n5559\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__15578\,
            I => \N__15575\
        );

    \I__2247\ : InMux
    port map (
            O => \N__15575\,
            I => \N__15572\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__15572\,
            I => \eeprom.n3714\
        );

    \I__2245\ : InMux
    port map (
            O => \N__15569\,
            I => \eeprom.n4238\
        );

    \I__2244\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__15560\,
            I => \eeprom.n5562\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__2240\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15551\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__15548\,
            I => \eeprom.n3713\
        );

    \I__2237\ : InMux
    port map (
            O => \N__15545\,
            I => \eeprom.n4239\
        );

    \I__2236\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15539\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__15539\,
            I => \eeprom.n5565\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__15536\,
            I => \N__15533\
        );

    \I__2233\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15530\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__15530\,
            I => \eeprom.n3712\
        );

    \I__2231\ : InMux
    port map (
            O => \N__15527\,
            I => \eeprom.n4240\
        );

    \I__2230\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15521\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__15521\,
            I => \eeprom.n3711\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__2227\ : InMux
    port map (
            O => \N__15515\,
            I => \N__15512\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__15512\,
            I => \N__15509\
        );

    \I__2225\ : Span4Mux_h
    port map (
            O => \N__15509\,
            I => \N__15506\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__15506\,
            I => \eeprom.n5568\
        );

    \I__2223\ : InMux
    port map (
            O => \N__15503\,
            I => \eeprom.n4241\
        );

    \I__2222\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15494\
        );

    \I__2221\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15494\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__15494\,
            I => \eeprom.n3716\
        );

    \I__2219\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15488\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__15488\,
            I => \eeprom.n5553\
        );

    \I__2217\ : InMux
    port map (
            O => \N__15485\,
            I => \N__15482\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__15482\,
            I => \N__15479\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__15476\,
            I => \eeprom.n3586\
        );

    \I__2213\ : InMux
    port map (
            O => \N__15473\,
            I => \bfn_20_19_0_\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__15470\,
            I => \N__15466\
        );

    \I__2211\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15462\
        );

    \I__2210\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15459\
        );

    \I__2209\ : InMux
    port map (
            O => \N__15465\,
            I => \N__15456\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__15462\,
            I => \eeprom.n3518\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__15459\,
            I => \eeprom.n3518\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__15456\,
            I => \eeprom.n3518\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__15449\,
            I => \N__15446\
        );

    \I__2204\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15443\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__15443\,
            I => \eeprom.n3585_adj_296\
        );

    \I__2202\ : InMux
    port map (
            O => \N__15440\,
            I => \eeprom.n4205\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__15437\,
            I => \N__15433\
        );

    \I__2200\ : InMux
    port map (
            O => \N__15436\,
            I => \N__15430\
        );

    \I__2199\ : InMux
    port map (
            O => \N__15433\,
            I => \N__15427\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__15430\,
            I => \N__15423\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__15427\,
            I => \N__15420\
        );

    \I__2196\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15417\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__15423\,
            I => \eeprom.n3517\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__15420\,
            I => \eeprom.n3517\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__15417\,
            I => \eeprom.n3517\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__15410\,
            I => \N__15407\
        );

    \I__2191\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15404\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__15404\,
            I => \N__15401\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__15401\,
            I => \eeprom.n3584\
        );

    \I__2188\ : InMux
    port map (
            O => \N__15398\,
            I => \eeprom.n4206\
        );

    \I__2187\ : InMux
    port map (
            O => \N__15395\,
            I => \eeprom.n4229\
        );

    \I__2186\ : InMux
    port map (
            O => \N__15392\,
            I => \eeprom.n4230\
        );

    \I__2185\ : InMux
    port map (
            O => \N__15389\,
            I => \eeprom.n4231\
        );

    \I__2184\ : InMux
    port map (
            O => \N__15386\,
            I => \eeprom.n4232\
        );

    \I__2183\ : InMux
    port map (
            O => \N__15383\,
            I => \eeprom.n4233\
        );

    \I__2182\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15377\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__15377\,
            I => \eeprom.n5547\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__15374\,
            I => \N__15371\
        );

    \I__2179\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15368\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__15368\,
            I => \eeprom.n5362\
        );

    \I__2177\ : InMux
    port map (
            O => \N__15365\,
            I => \eeprom.n4234\
        );

    \I__2176\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__15359\,
            I => \eeprom.n5550\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__15356\,
            I => \N__15353\
        );

    \I__2173\ : InMux
    port map (
            O => \N__15353\,
            I => \N__15350\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__15350\,
            I => \eeprom.n3717\
        );

    \I__2171\ : InMux
    port map (
            O => \N__15347\,
            I => \bfn_20_18_0_\
        );

    \I__2170\ : InMux
    port map (
            O => \N__15344\,
            I => \eeprom.n4236\
        );

    \I__2169\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15338\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__15338\,
            I => \eeprom.n5556\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__15335\,
            I => \N__15332\
        );

    \I__2166\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15329\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__15329\,
            I => \eeprom.n3715\
        );

    \I__2164\ : InMux
    port map (
            O => \N__15326\,
            I => \eeprom.n4237\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__15323\,
            I => \N__15320\
        );

    \I__2162\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15316\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__15319\,
            I => \N__15313\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__15316\,
            I => \N__15309\
        );

    \I__2159\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15306\
        );

    \I__2158\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15303\
        );

    \I__2157\ : Span4Mux_h
    port map (
            O => \N__15309\,
            I => \N__15300\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__15306\,
            I => \N__15295\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15295\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__15300\,
            I => \eeprom.n3105\
        );

    \I__2153\ : Odrv12
    port map (
            O => \N__15295\,
            I => \eeprom.n3105\
        );

    \I__2152\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15287\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__15287\,
            I => \N__15284\
        );

    \I__2150\ : Sp12to4
    port map (
            O => \N__15284\,
            I => \N__15281\
        );

    \I__2149\ : Odrv12
    port map (
            O => \N__15281\,
            I => \eeprom.n3172\
        );

    \I__2148\ : InMux
    port map (
            O => \N__15278\,
            I => \eeprom.n4136\
        );

    \I__2147\ : InMux
    port map (
            O => \N__15275\,
            I => \N__15272\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__15272\,
            I => \N__15267\
        );

    \I__2145\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15264\
        );

    \I__2144\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15261\
        );

    \I__2143\ : Span4Mux_h
    port map (
            O => \N__15267\,
            I => \N__15258\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__15264\,
            I => \N__15255\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__15261\,
            I => \N__15252\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__15258\,
            I => \eeprom.n3104\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__15255\,
            I => \eeprom.n3104\
        );

    \I__2138\ : Odrv12
    port map (
            O => \N__15252\,
            I => \eeprom.n3104\
        );

    \I__2137\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__15242\,
            I => \N__15239\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__15236\,
            I => \eeprom.n3171\
        );

    \I__2133\ : InMux
    port map (
            O => \N__15233\,
            I => \eeprom.n4137\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__2131\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15222\
        );

    \I__2130\ : InMux
    port map (
            O => \N__15226\,
            I => \N__15219\
        );

    \I__2129\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15216\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__15222\,
            I => \N__15211\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__15219\,
            I => \N__15211\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__15216\,
            I => \eeprom.n3103\
        );

    \I__2125\ : Odrv12
    port map (
            O => \N__15211\,
            I => \eeprom.n3103\
        );

    \I__2124\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__15203\,
            I => \N__15200\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__15200\,
            I => \N__15197\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__15197\,
            I => \eeprom.n3170\
        );

    \I__2120\ : InMux
    port map (
            O => \N__15194\,
            I => \bfn_19_32_0_\
        );

    \I__2119\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15188\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__15188\,
            I => \N__15185\
        );

    \I__2117\ : Span4Mux_s2_v
    port map (
            O => \N__15185\,
            I => \N__15180\
        );

    \I__2116\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15175\
        );

    \I__2115\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15175\
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__15180\,
            I => \eeprom.n3102\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__15175\,
            I => \eeprom.n3102\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__2111\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15164\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__15164\,
            I => \N__15161\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__15161\,
            I => \N__15158\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__15158\,
            I => \eeprom.n3169\
        );

    \I__2107\ : InMux
    port map (
            O => \N__15155\,
            I => \eeprom.n4139\
        );

    \I__2106\ : InMux
    port map (
            O => \N__15152\,
            I => \N__15148\
        );

    \I__2105\ : InMux
    port map (
            O => \N__15151\,
            I => \N__15145\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__15148\,
            I => \N__15142\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__15145\,
            I => \N__15138\
        );

    \I__2102\ : Span4Mux_s3_v
    port map (
            O => \N__15142\,
            I => \N__15135\
        );

    \I__2101\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15132\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__15138\,
            I => \eeprom.n3101\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__15135\,
            I => \eeprom.n3101\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__15132\,
            I => \eeprom.n3101\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__15125\,
            I => \N__15122\
        );

    \I__2096\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15119\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__15119\,
            I => \N__15116\
        );

    \I__2094\ : Span4Mux_h
    port map (
            O => \N__15116\,
            I => \N__15113\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__15113\,
            I => \N__15110\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__15110\,
            I => \eeprom.n3168\
        );

    \I__2091\ : InMux
    port map (
            O => \N__15107\,
            I => \eeprom.n4140\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__2089\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15097\
        );

    \I__2088\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15094\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__15097\,
            I => \N__15091\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__15094\,
            I => \eeprom.n3100\
        );

    \I__2085\ : Odrv12
    port map (
            O => \N__15091\,
            I => \eeprom.n3100\
        );

    \I__2084\ : InMux
    port map (
            O => \N__15086\,
            I => \eeprom.n4141\
        );

    \I__2083\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15079\
        );

    \I__2082\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15076\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__15079\,
            I => \N__15073\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__15076\,
            I => \N__15070\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__15073\,
            I => \N__15067\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__15070\,
            I => \N__15064\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__15067\,
            I => \N__15061\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__15064\,
            I => \eeprom.n3199\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__15061\,
            I => \eeprom.n3199\
        );

    \I__2074\ : InMux
    port map (
            O => \N__15056\,
            I => \bfn_20_17_0_\
        );

    \I__2073\ : InMux
    port map (
            O => \N__15053\,
            I => \eeprom.n4228\
        );

    \I__2072\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15046\
        );

    \I__2071\ : InMux
    port map (
            O => \N__15049\,
            I => \N__15043\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__15046\,
            I => \N__15040\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__15043\,
            I => \eeprom.n3113\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__15040\,
            I => \eeprom.n3113\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__15035\,
            I => \N__15032\
        );

    \I__2066\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15029\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__15029\,
            I => \N__15026\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__15026\,
            I => \N__15023\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__15023\,
            I => \eeprom.n3180\
        );

    \I__2062\ : InMux
    port map (
            O => \N__15020\,
            I => \eeprom.n4128\
        );

    \I__2061\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15014\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__15014\,
            I => \N__15011\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__15011\,
            I => \N__15008\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__15008\,
            I => \eeprom.n3179\
        );

    \I__2057\ : InMux
    port map (
            O => \N__15005\,
            I => \eeprom.n4129\
        );

    \I__2056\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__14999\,
            I => \N__14994\
        );

    \I__2054\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14991\
        );

    \I__2053\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14988\
        );

    \I__2052\ : Span4Mux_s3_v
    port map (
            O => \N__14994\,
            I => \N__14985\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__14991\,
            I => \N__14980\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__14988\,
            I => \N__14980\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__14985\,
            I => \eeprom.n3111\
        );

    \I__2048\ : Odrv4
    port map (
            O => \N__14980\,
            I => \eeprom.n3111\
        );

    \I__2047\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14972\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__14966\,
            I => \eeprom.n3178\
        );

    \I__2043\ : InMux
    port map (
            O => \N__14963\,
            I => \bfn_19_31_0_\
        );

    \I__2042\ : InMux
    port map (
            O => \N__14960\,
            I => \eeprom.n4131\
        );

    \I__2041\ : InMux
    port map (
            O => \N__14957\,
            I => \eeprom.n4132\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__14954\,
            I => \N__14951\
        );

    \I__2039\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14947\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__14950\,
            I => \N__14944\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__14947\,
            I => \N__14941\
        );

    \I__2036\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14938\
        );

    \I__2035\ : Span4Mux_v
    port map (
            O => \N__14941\,
            I => \N__14935\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__14938\,
            I => \eeprom.n3108\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__14935\,
            I => \eeprom.n3108\
        );

    \I__2032\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14927\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__14924\,
            I => \N__14921\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__14921\,
            I => \eeprom.n3175\
        );

    \I__2028\ : InMux
    port map (
            O => \N__14918\,
            I => \eeprom.n4133\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__14915\,
            I => \N__14911\
        );

    \I__2026\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14907\
        );

    \I__2025\ : InMux
    port map (
            O => \N__14911\,
            I => \N__14902\
        );

    \I__2024\ : InMux
    port map (
            O => \N__14910\,
            I => \N__14902\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__14907\,
            I => \N__14899\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__14902\,
            I => \N__14896\
        );

    \I__2021\ : Odrv4
    port map (
            O => \N__14899\,
            I => \eeprom.n3107\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__14896\,
            I => \eeprom.n3107\
        );

    \I__2019\ : InMux
    port map (
            O => \N__14891\,
            I => \N__14888\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__14888\,
            I => \N__14885\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__14885\,
            I => \N__14882\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__14882\,
            I => \eeprom.n3174\
        );

    \I__2015\ : InMux
    port map (
            O => \N__14879\,
            I => \eeprom.n4134\
        );

    \I__2014\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14871\
        );

    \I__2013\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14866\
        );

    \I__2012\ : InMux
    port map (
            O => \N__14874\,
            I => \N__14866\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__14871\,
            I => \N__14863\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__14866\,
            I => \N__14860\
        );

    \I__2009\ : Odrv12
    port map (
            O => \N__14863\,
            I => \eeprom.n3106\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__14860\,
            I => \eeprom.n3106\
        );

    \I__2007\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__14852\,
            I => \N__14849\
        );

    \I__2005\ : Odrv12
    port map (
            O => \N__14849\,
            I => \eeprom.n3173\
        );

    \I__2004\ : InMux
    port map (
            O => \N__14846\,
            I => \eeprom.n4135\
        );

    \I__2003\ : InMux
    port map (
            O => \N__14843\,
            I => \N__14836\
        );

    \I__2002\ : InMux
    port map (
            O => \N__14842\,
            I => \N__14836\
        );

    \I__2001\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14833\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__14836\,
            I => \eeprom.n3012\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__14833\,
            I => \eeprom.n3012\
        );

    \I__1998\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14824\
        );

    \I__1997\ : InMux
    port map (
            O => \N__14827\,
            I => \N__14821\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__14824\,
            I => \N__14818\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__14821\,
            I => \N__14814\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__14818\,
            I => \N__14811\
        );

    \I__1993\ : InMux
    port map (
            O => \N__14817\,
            I => \N__14808\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__14814\,
            I => \eeprom.n3003\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__14811\,
            I => \eeprom.n3003\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__14808\,
            I => \eeprom.n3003\
        );

    \I__1989\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__14798\,
            I => \eeprom.n3086\
        );

    \I__1987\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14792\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__14792\,
            I => \N__14789\
        );

    \I__1985\ : Span4Mux_h
    port map (
            O => \N__14789\,
            I => \N__14786\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__14786\,
            I => \N__14783\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__14783\,
            I => \eeprom.n3186\
        );

    \I__1982\ : InMux
    port map (
            O => \N__14780\,
            I => \bfn_19_30_0_\
        );

    \I__1981\ : InMux
    port map (
            O => \N__14777\,
            I => \eeprom.n4123\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__14774\,
            I => \N__14770\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__14773\,
            I => \N__14767\
        );

    \I__1978\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14764\
        );

    \I__1977\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14760\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__14764\,
            I => \N__14757\
        );

    \I__1975\ : InMux
    port map (
            O => \N__14763\,
            I => \N__14754\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__14760\,
            I => \N__14751\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__14757\,
            I => \eeprom.n3117\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__14754\,
            I => \eeprom.n3117\
        );

    \I__1971\ : Odrv4
    port map (
            O => \N__14751\,
            I => \eeprom.n3117\
        );

    \I__1970\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14741\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__14741\,
            I => \N__14738\
        );

    \I__1968\ : Odrv12
    port map (
            O => \N__14738\,
            I => \eeprom.n3184\
        );

    \I__1967\ : InMux
    port map (
            O => \N__14735\,
            I => \eeprom.n4124\
        );

    \I__1966\ : InMux
    port map (
            O => \N__14732\,
            I => \eeprom.n4125\
        );

    \I__1965\ : InMux
    port map (
            O => \N__14729\,
            I => \eeprom.n4126\
        );

    \I__1964\ : InMux
    port map (
            O => \N__14726\,
            I => \eeprom.n4127\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__14723\,
            I => \N__14720\
        );

    \I__1962\ : InMux
    port map (
            O => \N__14720\,
            I => \N__14717\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__14717\,
            I => \N__14713\
        );

    \I__1960\ : InMux
    port map (
            O => \N__14716\,
            I => \N__14710\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__14713\,
            I => \eeprom.n3007\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__14710\,
            I => \eeprom.n3007\
        );

    \I__1957\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14702\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__14702\,
            I => \N__14699\
        );

    \I__1955\ : Span4Mux_h
    port map (
            O => \N__14699\,
            I => \N__14696\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__14696\,
            I => \eeprom.n3074\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__14693\,
            I => \eeprom.n3007_cascade_\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__14690\,
            I => \N__14686\
        );

    \I__1951\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14683\
        );

    \I__1950\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14680\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__14683\,
            I => \N__14677\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__14680\,
            I => \eeprom.n3006\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__14677\,
            I => \eeprom.n3006\
        );

    \I__1946\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14669\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__14669\,
            I => \eeprom.n21_adj_336\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__14666\,
            I => \eeprom.n3006_cascade_\
        );

    \I__1943\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__14660\,
            I => \N__14657\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__14657\,
            I => \eeprom.n18_adj_335\
        );

    \I__1940\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__14651\,
            I => \eeprom.n24_adj_340\
        );

    \I__1938\ : CascadeMux
    port map (
            O => \N__14648\,
            I => \N__14645\
        );

    \I__1937\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14640\
        );

    \I__1936\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14637\
        );

    \I__1935\ : InMux
    port map (
            O => \N__14643\,
            I => \N__14634\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__14640\,
            I => \N__14631\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__14637\,
            I => \N__14626\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__14634\,
            I => \N__14626\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__14631\,
            I => \eeprom.n3008\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__14626\,
            I => \eeprom.n3008\
        );

    \I__1929\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14617\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__14620\,
            I => \N__14614\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__14617\,
            I => \N__14611\
        );

    \I__1926\ : InMux
    port map (
            O => \N__14614\,
            I => \N__14608\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__14611\,
            I => \eeprom.n3005\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__14608\,
            I => \eeprom.n3005\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \eeprom.n3005_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__14600\,
            I => \N__14597\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__14594\,
            I => \N__14591\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__14591\,
            I => \eeprom.n3072\
        );

    \I__1918\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14585\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__14585\,
            I => \eeprom.n3082\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__14582\,
            I => \N__14577\
        );

    \I__1915\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14572\
        );

    \I__1914\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14572\
        );

    \I__1913\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14569\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__14572\,
            I => \eeprom.n3010\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__14569\,
            I => \eeprom.n3010\
        );

    \I__1910\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14561\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__14561\,
            I => \N__14557\
        );

    \I__1908\ : InMux
    port map (
            O => \N__14560\,
            I => \N__14554\
        );

    \I__1907\ : Span12Mux_s6_v
    port map (
            O => \N__14557\,
            I => \N__14551\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__14554\,
            I => \eeprom.n3002\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__14551\,
            I => \eeprom.n3002\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__14546\,
            I => \eeprom.n3002_cascade_\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__14543\,
            I => \N__14540\
        );

    \I__1902\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14537\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__14537\,
            I => \N__14534\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__14534\,
            I => \N__14531\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__14531\,
            I => \eeprom.n20_adj_337\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__14528\,
            I => \N__14525\
        );

    \I__1897\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14522\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__14522\,
            I => \N__14519\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__14516\,
            I => \eeprom.n3078\
        );

    \I__1893\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14509\
        );

    \I__1892\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14505\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__14509\,
            I => \N__14502\
        );

    \I__1890\ : InMux
    port map (
            O => \N__14508\,
            I => \N__14499\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__14505\,
            I => \eeprom.n3016\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__14502\,
            I => \eeprom.n3016\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__14499\,
            I => \eeprom.n3016\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__14492\,
            I => \N__14488\
        );

    \I__1885\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14484\
        );

    \I__1884\ : InMux
    port map (
            O => \N__14488\,
            I => \N__14481\
        );

    \I__1883\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14478\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__14484\,
            I => \N__14475\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__14481\,
            I => \eeprom.n3018\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__14478\,
            I => \eeprom.n3018\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__14475\,
            I => \eeprom.n3018\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__14468\,
            I => \eeprom.n2914_cascade_\
        );

    \I__1877\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14459\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__14459\,
            I => \eeprom.n3073\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__1873\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14449\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__14452\,
            I => \N__14446\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__14449\,
            I => \N__14443\
        );

    \I__1870\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14439\
        );

    \I__1869\ : Span4Mux_h
    port map (
            O => \N__14443\,
            I => \N__14436\
        );

    \I__1868\ : InMux
    port map (
            O => \N__14442\,
            I => \N__14433\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__14439\,
            I => \eeprom.n3014\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__14436\,
            I => \eeprom.n3014\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__14433\,
            I => \eeprom.n3014\
        );

    \I__1864\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14423\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__14423\,
            I => \N__14419\
        );

    \I__1862\ : InMux
    port map (
            O => \N__14422\,
            I => \N__14416\
        );

    \I__1861\ : Span4Mux_h
    port map (
            O => \N__14419\,
            I => \N__14413\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__14416\,
            I => \eeprom.n3205\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__14413\,
            I => \eeprom.n3205\
        );

    \I__1858\ : InMux
    port map (
            O => \N__14408\,
            I => \N__14405\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__14405\,
            I => \N__14402\
        );

    \I__1856\ : Span4Mux_h
    port map (
            O => \N__14402\,
            I => \N__14399\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__14399\,
            I => \eeprom.n3272\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__14396\,
            I => \eeprom.n3205_cascade_\
        );

    \I__1853\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14389\
        );

    \I__1852\ : InMux
    port map (
            O => \N__14392\,
            I => \N__14386\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__14386\,
            I => \eeprom.n3204\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__14383\,
            I => \eeprom.n3204\
        );

    \I__1848\ : InMux
    port map (
            O => \N__14378\,
            I => \N__14375\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__14375\,
            I => \N__14372\
        );

    \I__1846\ : Span4Mux_h
    port map (
            O => \N__14372\,
            I => \N__14369\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__14369\,
            I => \eeprom.n3271\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__14366\,
            I => \N__14363\
        );

    \I__1843\ : InMux
    port map (
            O => \N__14363\,
            I => \N__14360\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__14360\,
            I => \N__14355\
        );

    \I__1841\ : InMux
    port map (
            O => \N__14359\,
            I => \N__14350\
        );

    \I__1840\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14350\
        );

    \I__1839\ : Span4Mux_h
    port map (
            O => \N__14355\,
            I => \N__14347\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__14350\,
            I => \eeprom.n3207\
        );

    \I__1837\ : Odrv4
    port map (
            O => \N__14347\,
            I => \eeprom.n3207\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__14342\,
            I => \N__14339\
        );

    \I__1835\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14336\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__14336\,
            I => \N__14332\
        );

    \I__1833\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14329\
        );

    \I__1832\ : Span4Mux_v
    port map (
            O => \N__14332\,
            I => \N__14326\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__14329\,
            I => \eeprom.n3017\
        );

    \I__1830\ : Odrv4
    port map (
            O => \N__14326\,
            I => \eeprom.n3017\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__14321\,
            I => \eeprom.n3017_cascade_\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__14318\,
            I => \eeprom.n5147_cascade_\
        );

    \I__1827\ : InMux
    port map (
            O => \N__14315\,
            I => \N__14311\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__14314\,
            I => \N__14308\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__14311\,
            I => \N__14305\
        );

    \I__1824\ : InMux
    port map (
            O => \N__14308\,
            I => \N__14301\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__14305\,
            I => \N__14298\
        );

    \I__1822\ : InMux
    port map (
            O => \N__14304\,
            I => \N__14295\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__14301\,
            I => \eeprom.n3009\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__14298\,
            I => \eeprom.n3009\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__14295\,
            I => \eeprom.n3009\
        );

    \I__1818\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14284\
        );

    \I__1817\ : InMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__14284\,
            I => \N__14278\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__14281\,
            I => \eeprom.n3206\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__14278\,
            I => \eeprom.n3206\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__14273\,
            I => \eeprom.n20_adj_301_cascade_\
        );

    \I__1812\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14267\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__14267\,
            I => \eeprom.n16_adj_303\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__14264\,
            I => \N__14261\
        );

    \I__1809\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14256\
        );

    \I__1808\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14253\
        );

    \I__1807\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14250\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__14256\,
            I => \N__14245\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__14253\,
            I => \N__14245\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__14250\,
            I => \eeprom.n3212\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__14245\,
            I => \eeprom.n3212\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__14240\,
            I => \eeprom.n28_adj_305_cascade_\
        );

    \I__1801\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14234\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__14234\,
            I => \eeprom.n24_adj_304\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__14231\,
            I => \eeprom.n3232_cascade_\
        );

    \I__1798\ : InMux
    port map (
            O => \N__14228\,
            I => \N__14225\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__14222\,
            I => \N__14219\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__14219\,
            I => \eeprom.n3274\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__14216\,
            I => \N__14213\
        );

    \I__1793\ : InMux
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__14210\,
            I => \N__14206\
        );

    \I__1791\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14203\
        );

    \I__1790\ : Span4Mux_v
    port map (
            O => \N__14206\,
            I => \N__14200\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__14203\,
            I => \eeprom.n3306\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__14200\,
            I => \eeprom.n3306\
        );

    \I__1787\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14191\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__14194\,
            I => \N__14188\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__14191\,
            I => \N__14184\
        );

    \I__1784\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14181\
        );

    \I__1783\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14178\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__14184\,
            I => \eeprom.n3305\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__14181\,
            I => \eeprom.n3305\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__14178\,
            I => \eeprom.n3305\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__14171\,
            I => \eeprom.n3306_cascade_\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__14168\,
            I => \N__14165\
        );

    \I__1777\ : InMux
    port map (
            O => \N__14165\,
            I => \N__14161\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14154\
        );

    \I__1774\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14151\
        );

    \I__1773\ : InMux
    port map (
            O => \N__14157\,
            I => \N__14148\
        );

    \I__1772\ : Odrv4
    port map (
            O => \N__14154\,
            I => \eeprom.n3308\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__14151\,
            I => \eeprom.n3308\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__14148\,
            I => \eeprom.n3308\
        );

    \I__1769\ : InMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__14138\,
            I => \eeprom.n27\
        );

    \I__1767\ : InMux
    port map (
            O => \N__14135\,
            I => \N__14132\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__14132\,
            I => \N__14129\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__14129\,
            I => \eeprom.n5309\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__14126\,
            I => \eeprom.n18_adj_260_cascade_\
        );

    \I__1763\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14120\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__14120\,
            I => \eeprom.n24\
        );

    \I__1761\ : InMux
    port map (
            O => \N__14117\,
            I => \N__14114\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__14114\,
            I => \eeprom.n22\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__14111\,
            I => \eeprom.n26_adj_262_cascade_\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__14108\,
            I => \eeprom.n3133_cascade_\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__14105\,
            I => \N__14102\
        );

    \I__1756\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14099\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__14099\,
            I => \N__14096\
        );

    \I__1754\ : Span4Mux_h
    port map (
            O => \N__14096\,
            I => \N__14093\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__14093\,
            I => \eeprom.n3373\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__1751\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14084\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__14084\,
            I => \N__14081\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__14081\,
            I => \N__14078\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__14078\,
            I => \eeprom.n3369\
        );

    \I__1747\ : InMux
    port map (
            O => \N__14075\,
            I => \N__14071\
        );

    \I__1746\ : InMux
    port map (
            O => \N__14074\,
            I => \N__14068\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__14068\,
            I => \N__14062\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__14065\,
            I => \eeprom.n3401\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__14062\,
            I => \eeprom.n3401\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__14057\,
            I => \N__14053\
        );

    \I__1740\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14049\
        );

    \I__1739\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14046\
        );

    \I__1738\ : InMux
    port map (
            O => \N__14052\,
            I => \N__14043\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__14049\,
            I => \eeprom.n3400\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__14046\,
            I => \eeprom.n3400\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__14043\,
            I => \eeprom.n3400\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__14036\,
            I => \N__14032\
        );

    \I__1733\ : InMux
    port map (
            O => \N__14035\,
            I => \N__14028\
        );

    \I__1732\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14025\
        );

    \I__1731\ : InMux
    port map (
            O => \N__14031\,
            I => \N__14022\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__14028\,
            I => \eeprom.n3399\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__14025\,
            I => \eeprom.n3399\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__14022\,
            I => \eeprom.n3399\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__14015\,
            I => \eeprom.n3401_cascade_\
        );

    \I__1726\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__14009\,
            I => \eeprom.n27_adj_263\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__14006\,
            I => \N__14003\
        );

    \I__1723\ : InMux
    port map (
            O => \N__14003\,
            I => \N__13998\
        );

    \I__1722\ : InMux
    port map (
            O => \N__14002\,
            I => \N__13993\
        );

    \I__1721\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13993\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__13998\,
            I => \eeprom.n3402\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__13993\,
            I => \eeprom.n3402\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__1717\ : InMux
    port map (
            O => \N__13985\,
            I => \N__13982\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__13979\,
            I => \eeprom.n3469\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__13976\,
            I => \N__13972\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__1712\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13965\
        );

    \I__1711\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13962\
        );

    \I__1710\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13959\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__13965\,
            I => \eeprom.n3307\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__13962\,
            I => \eeprom.n3307\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__13959\,
            I => \eeprom.n3307\
        );

    \I__1706\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13947\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__13951\,
            I => \N__13944\
        );

    \I__1704\ : InMux
    port map (
            O => \N__13950\,
            I => \N__13941\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__13947\,
            I => \N__13938\
        );

    \I__1702\ : InMux
    port map (
            O => \N__13944\,
            I => \N__13935\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__13941\,
            I => \N__13932\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__13938\,
            I => \eeprom.n3311\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__13935\,
            I => \eeprom.n3311\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__13932\,
            I => \eeprom.n3311\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__13925\,
            I => \N__13920\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__13924\,
            I => \N__13917\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__13923\,
            I => \N__13914\
        );

    \I__1694\ : InMux
    port map (
            O => \N__13920\,
            I => \N__13911\
        );

    \I__1693\ : InMux
    port map (
            O => \N__13917\,
            I => \N__13908\
        );

    \I__1692\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13905\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__13911\,
            I => \eeprom.n3312\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__13908\,
            I => \eeprom.n3312\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__13905\,
            I => \eeprom.n3312\
        );

    \I__1688\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13894\
        );

    \I__1687\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13891\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__13894\,
            I => \N__13887\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13884\
        );

    \I__1684\ : InMux
    port map (
            O => \N__13890\,
            I => \N__13881\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__13887\,
            I => \N__13876\
        );

    \I__1682\ : Span4Mux_h
    port map (
            O => \N__13884\,
            I => \N__13876\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__13881\,
            I => \eeprom.n3309\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__13876\,
            I => \eeprom.n3309\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \eeprom.n28_cascade_\
        );

    \I__1678\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13865\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__13865\,
            I => \eeprom.n25\
        );

    \I__1676\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13859\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__13859\,
            I => \N__13856\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__13856\,
            I => \N__13853\
        );

    \I__1673\ : Odrv4
    port map (
            O => \N__13853\,
            I => \eeprom.n3385\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__13850\,
            I => \eeprom.n3331_cascade_\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__13847\,
            I => \N__13844\
        );

    \I__1670\ : InMux
    port map (
            O => \N__13844\,
            I => \N__13841\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__1668\ : Span4Mux_v
    port map (
            O => \N__13838\,
            I => \N__13835\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__13835\,
            I => \eeprom.n3281\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__13832\,
            I => \N__13829\
        );

    \I__1665\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13826\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__13826\,
            I => \N__13823\
        );

    \I__1663\ : Odrv4
    port map (
            O => \N__13823\,
            I => \eeprom.n3485\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__13820\,
            I => \N__13815\
        );

    \I__1661\ : InMux
    port map (
            O => \N__13819\,
            I => \N__13812\
        );

    \I__1660\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13809\
        );

    \I__1659\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13806\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__13812\,
            I => \eeprom.n3398\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__13809\,
            I => \eeprom.n3398\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__13806\,
            I => \eeprom.n3398\
        );

    \I__1655\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13795\
        );

    \I__1654\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13792\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__13795\,
            I => \N__13789\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__13792\,
            I => \N__13784\
        );

    \I__1651\ : Span4Mux_h
    port map (
            O => \N__13789\,
            I => \N__13784\
        );

    \I__1650\ : Odrv4
    port map (
            O => \N__13784\,
            I => \eeprom.n3397\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__13781\,
            I => \N__13776\
        );

    \I__1648\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13773\
        );

    \I__1647\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13770\
        );

    \I__1646\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13767\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__13773\,
            I => \eeprom.n3408\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__13770\,
            I => \eeprom.n3408\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__13767\,
            I => \eeprom.n3408\
        );

    \I__1642\ : InMux
    port map (
            O => \N__13760\,
            I => \N__13756\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__13759\,
            I => \N__13752\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__13756\,
            I => \N__13749\
        );

    \I__1639\ : InMux
    port map (
            O => \N__13755\,
            I => \N__13746\
        );

    \I__1638\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13743\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__13749\,
            I => \eeprom.n3411\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__13746\,
            I => \eeprom.n3411\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__13743\,
            I => \eeprom.n3411\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__13736\,
            I => \eeprom.n18_cascade_\
        );

    \I__1633\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13730\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__13730\,
            I => \eeprom.n29\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__13727\,
            I => \eeprom.n30_cascade_\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__13724\,
            I => \eeprom.n3430_cascade_\
        );

    \I__1629\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13718\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__13718\,
            I => \N__13715\
        );

    \I__1627\ : Span4Mux_h
    port map (
            O => \N__13715\,
            I => \N__13712\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__13712\,
            I => \eeprom.n3467\
        );

    \I__1625\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13706\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__13706\,
            I => \N__13703\
        );

    \I__1623\ : Span4Mux_h
    port map (
            O => \N__13703\,
            I => \N__13700\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__13700\,
            I => \eeprom.n3466\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__13697\,
            I => \eeprom.n3498_cascade_\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__13694\,
            I => \N__13691\
        );

    \I__1619\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13688\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__13688\,
            I => \N__13685\
        );

    \I__1617\ : Odrv4
    port map (
            O => \N__13685\,
            I => \eeprom.n28_adj_267\
        );

    \I__1616\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13679\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__13679\,
            I => \N__13676\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__13676\,
            I => \eeprom.n3476\
        );

    \I__1613\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13670\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__13670\,
            I => \N__13667\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__13667\,
            I => \N__13664\
        );

    \I__1610\ : Odrv4
    port map (
            O => \N__13664\,
            I => \eeprom.n3486\
        );

    \I__1609\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13658\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__13658\,
            I => \N__13655\
        );

    \I__1607\ : Span4Mux_h
    port map (
            O => \N__13655\,
            I => \N__13652\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__13652\,
            I => \eeprom.n3468\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__13649\,
            I => \eeprom.n3608_cascade_\
        );

    \I__1604\ : InMux
    port map (
            O => \N__13646\,
            I => \N__13643\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__13640\,
            I => \eeprom.n3480\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__13637\,
            I => \eeprom.n3512_cascade_\
        );

    \I__1600\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13631\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__13631\,
            I => \eeprom.n5175\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__13628\,
            I => \eeprom.n5177_cascade_\
        );

    \I__1597\ : InMux
    port map (
            O => \N__13625\,
            I => \N__13622\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__13622\,
            I => \N__13619\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__13619\,
            I => \eeprom.n31_adj_341\
        );

    \I__1594\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13613\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__13613\,
            I => \N__13610\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__13610\,
            I => \eeprom.n3598\
        );

    \I__1591\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13604\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__13604\,
            I => \N__13601\
        );

    \I__1589\ : Odrv12
    port map (
            O => \N__13601\,
            I => \eeprom.n3483\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__13598\,
            I => \eeprom.n5031_cascade_\
        );

    \I__1587\ : InMux
    port map (
            O => \N__13595\,
            I => \N__13592\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__13592\,
            I => \eeprom.n5161\
        );

    \I__1585\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13586\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__13586\,
            I => \eeprom.n29_adj_274\
        );

    \I__1583\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13576\
        );

    \I__1581\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13573\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__13576\,
            I => \eeprom.n3612\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__13573\,
            I => \eeprom.n3612\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__13568\,
            I => \N__13564\
        );

    \I__1577\ : InMux
    port map (
            O => \N__13567\,
            I => \N__13561\
        );

    \I__1576\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13558\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__13561\,
            I => \N__13552\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__13558\,
            I => \N__13552\
        );

    \I__1573\ : InMux
    port map (
            O => \N__13557\,
            I => \N__13549\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__13552\,
            I => \eeprom.n3617\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__13549\,
            I => \eeprom.n3617\
        );

    \I__1570\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13541\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__13541\,
            I => \N__13538\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__13538\,
            I => \eeprom.n3596\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__13535\,
            I => \eeprom.n3609_cascade_\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__13532\,
            I => \eeprom.n5021_cascade_\
        );

    \I__1565\ : InMux
    port map (
            O => \N__13529\,
            I => \N__13526\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__13526\,
            I => \eeprom.n5023\
        );

    \I__1563\ : InMux
    port map (
            O => \N__13523\,
            I => \N__13520\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__13520\,
            I => \N__13517\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__13517\,
            I => \N__13514\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__13514\,
            I => \eeprom.n3474\
        );

    \I__1559\ : InMux
    port map (
            O => \N__13511\,
            I => \N__13506\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__13510\,
            I => \N__13503\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__13509\,
            I => \N__13500\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__13506\,
            I => \N__13497\
        );

    \I__1555\ : InMux
    port map (
            O => \N__13503\,
            I => \N__13494\
        );

    \I__1554\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13491\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__13497\,
            I => \eeprom.n3407\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__13494\,
            I => \eeprom.n3407\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__13491\,
            I => \eeprom.n3407\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__13484\,
            I => \eeprom.n5019_cascade_\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__13481\,
            I => \eeprom.n28_adj_342_cascade_\
        );

    \I__1548\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13474\
        );

    \I__1547\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13471\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__13474\,
            I => \N__13468\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__13471\,
            I => \eeprom.n3615\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__13468\,
            I => \eeprom.n3615\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__13463\,
            I => \eeprom.n3628_cascade_\
        );

    \I__1542\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13457\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__13457\,
            I => \eeprom.n1204\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__13454\,
            I => \eeprom.n3714_cascade_\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__13451\,
            I => \N__13447\
        );

    \I__1538\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13444\
        );

    \I__1537\ : InMux
    port map (
            O => \N__13447\,
            I => \N__13441\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__13444\,
            I => \eeprom.n1201\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__13441\,
            I => \eeprom.n1201\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__13436\,
            I => \N__13431\
        );

    \I__1533\ : InMux
    port map (
            O => \N__13435\,
            I => \N__13421\
        );

    \I__1532\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13421\
        );

    \I__1531\ : InMux
    port map (
            O => \N__13431\,
            I => \N__13416\
        );

    \I__1530\ : InMux
    port map (
            O => \N__13430\,
            I => \N__13416\
        );

    \I__1529\ : InMux
    port map (
            O => \N__13429\,
            I => \N__13407\
        );

    \I__1528\ : InMux
    port map (
            O => \N__13428\,
            I => \N__13407\
        );

    \I__1527\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13407\
        );

    \I__1526\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13407\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__13421\,
            I => \eeprom.n3628\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__13416\,
            I => \eeprom.n3628\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__13407\,
            I => \eeprom.n3628\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__13400\,
            I => \eeprom.n5025_cascade_\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__13397\,
            I => \eeprom.n5027_cascade_\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__13394\,
            I => \eeprom.n5029_cascade_\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__13391\,
            I => \eeprom.n3712_cascade_\
        );

    \I__1518\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13385\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__13385\,
            I => \eeprom.n1207\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__13382\,
            I => \N__13379\
        );

    \I__1515\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13375\
        );

    \I__1514\ : InMux
    port map (
            O => \N__13378\,
            I => \N__13372\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__13375\,
            I => \eeprom.n3618\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__13372\,
            I => \eeprom.n3618\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__13367\,
            I => \eeprom.n3717_cascade_\
        );

    \I__1510\ : InMux
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__13361\,
            I => \eeprom.n1208\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__13358\,
            I => \eeprom.n5362_cascade_\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__13355\,
            I => \N__13352\
        );

    \I__1506\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13349\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__13349\,
            I => \eeprom.n1206\
        );

    \I__1504\ : InMux
    port map (
            O => \N__13346\,
            I => \N__13343\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__13343\,
            I => \eeprom.n1205\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__13340\,
            I => \N__13336\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__13339\,
            I => \N__13333\
        );

    \I__1500\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13330\
        );

    \I__1499\ : InMux
    port map (
            O => \N__13333\,
            I => \N__13326\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__13330\,
            I => \N__13323\
        );

    \I__1497\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13320\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__13326\,
            I => \eeprom.n3616\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__13323\,
            I => \eeprom.n3616\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__13320\,
            I => \eeprom.n3616\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__13313\,
            I => \eeprom.n3715_cascade_\
        );

    \I__1492\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__13307\,
            I => \eeprom.n5017\
        );

    \I__1490\ : InMux
    port map (
            O => \N__13304\,
            I => \eeprom.n4116\
        );

    \I__1489\ : InMux
    port map (
            O => \N__13301\,
            I => \eeprom.n4117\
        );

    \I__1488\ : InMux
    port map (
            O => \N__13298\,
            I => \eeprom.n4118\
        );

    \I__1487\ : InMux
    port map (
            O => \N__13295\,
            I => \eeprom.n4119\
        );

    \I__1486\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13289\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__13289\,
            I => \N__13286\
        );

    \I__1484\ : Span4Mux_h
    port map (
            O => \N__13286\,
            I => \N__13283\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__13283\,
            I => \eeprom.n3070\
        );

    \I__1482\ : InMux
    port map (
            O => \N__13280\,
            I => \bfn_18_31_0_\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__13277\,
            I => \N__13274\
        );

    \I__1480\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13271\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__1478\ : Span4Mux_h
    port map (
            O => \N__13268\,
            I => \N__13265\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__13265\,
            I => \eeprom.n3069\
        );

    \I__1476\ : InMux
    port map (
            O => \N__13262\,
            I => \eeprom.n4121\
        );

    \I__1475\ : InMux
    port map (
            O => \N__13259\,
            I => \eeprom.n4122\
        );

    \I__1474\ : InMux
    port map (
            O => \N__13256\,
            I => \N__13253\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__13253\,
            I => \eeprom.n3071\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__13250\,
            I => \N__13247\
        );

    \I__1471\ : InMux
    port map (
            O => \N__13247\,
            I => \N__13242\
        );

    \I__1470\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13239\
        );

    \I__1469\ : InMux
    port map (
            O => \N__13245\,
            I => \N__13236\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__13242\,
            I => \N__13231\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__13239\,
            I => \N__13231\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__13236\,
            I => \eeprom.n3004\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__13231\,
            I => \eeprom.n3004\
        );

    \I__1464\ : InMux
    port map (
            O => \N__13226\,
            I => \N__13222\
        );

    \I__1463\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13219\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__13222\,
            I => \N__13215\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__13219\,
            I => \N__13212\
        );

    \I__1460\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13209\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__13215\,
            I => \eeprom.n3613\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__13212\,
            I => \eeprom.n3613\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__13209\,
            I => \eeprom.n3613\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__1455\ : InMux
    port map (
            O => \N__13199\,
            I => \N__13196\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__13196\,
            I => \eeprom.n1202\
        );

    \I__1453\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__13190\,
            I => \eeprom.n3083\
        );

    \I__1451\ : InMux
    port map (
            O => \N__13187\,
            I => \eeprom.n4107\
        );

    \I__1450\ : InMux
    port map (
            O => \N__13184\,
            I => \eeprom.n4108\
        );

    \I__1449\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13178\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__13178\,
            I => \N__13175\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__13175\,
            I => \eeprom.n3081\
        );

    \I__1446\ : InMux
    port map (
            O => \N__13172\,
            I => \eeprom.n4109\
        );

    \I__1445\ : InMux
    port map (
            O => \N__13169\,
            I => \eeprom.n4110\
        );

    \I__1444\ : InMux
    port map (
            O => \N__13166\,
            I => \N__13163\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__13163\,
            I => \eeprom.n3079\
        );

    \I__1442\ : InMux
    port map (
            O => \N__13160\,
            I => \eeprom.n4111\
        );

    \I__1441\ : InMux
    port map (
            O => \N__13157\,
            I => \bfn_18_30_0_\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__13154\,
            I => \N__13151\
        );

    \I__1439\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13148\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__13148\,
            I => \N__13145\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__13145\,
            I => \eeprom.n3077\
        );

    \I__1436\ : InMux
    port map (
            O => \N__13142\,
            I => \eeprom.n4113\
        );

    \I__1435\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__13136\,
            I => \N__13133\
        );

    \I__1433\ : Odrv12
    port map (
            O => \N__13133\,
            I => \eeprom.n3076\
        );

    \I__1432\ : InMux
    port map (
            O => \N__13130\,
            I => \eeprom.n4114\
        );

    \I__1431\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13124\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__13124\,
            I => \N__13121\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__13121\,
            I => \eeprom.n3075\
        );

    \I__1428\ : InMux
    port map (
            O => \N__13118\,
            I => \eeprom.n4115\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__13115\,
            I => \eeprom.n3034_cascade_\
        );

    \I__1426\ : InMux
    port map (
            O => \N__13112\,
            I => \bfn_18_29_0_\
        );

    \I__1425\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13106\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__13106\,
            I => \eeprom.n3085\
        );

    \I__1423\ : InMux
    port map (
            O => \N__13103\,
            I => \eeprom.n4105\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__13100\,
            I => \N__13097\
        );

    \I__1421\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13094\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__13094\,
            I => \N__13091\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__13091\,
            I => \eeprom.n3084\
        );

    \I__1418\ : InMux
    port map (
            O => \N__13088\,
            I => \eeprom.n4106\
        );

    \I__1417\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13082\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__13082\,
            I => \N__13079\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__13079\,
            I => \eeprom.n3270\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__13076\,
            I => \eeprom.n3203_cascade_\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__13073\,
            I => \eeprom.n3113_cascade_\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__13070\,
            I => \eeprom.n5305_cascade_\
        );

    \I__1411\ : InMux
    port map (
            O => \N__13067\,
            I => \N__13064\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__13064\,
            I => \N__13061\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__13061\,
            I => \eeprom.n3273\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__13058\,
            I => \eeprom.n3206_cascade_\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__13055\,
            I => \eeprom.n3108_cascade_\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__13052\,
            I => \N__13049\
        );

    \I__1405\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13045\
        );

    \I__1404\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13042\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__13045\,
            I => \N__13039\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__13042\,
            I => \N__13036\
        );

    \I__1401\ : Span4Mux_v
    port map (
            O => \N__13039\,
            I => \N__13030\
        );

    \I__1400\ : Span4Mux_h
    port map (
            O => \N__13036\,
            I => \N__13030\
        );

    \I__1399\ : InMux
    port map (
            O => \N__13035\,
            I => \N__13027\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__13030\,
            I => \eeprom.n3202\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__13027\,
            I => \eeprom.n3202\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__13022\,
            I => \N__13018\
        );

    \I__1395\ : InMux
    port map (
            O => \N__13021\,
            I => \N__13015\
        );

    \I__1394\ : InMux
    port map (
            O => \N__13018\,
            I => \N__13012\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__13015\,
            I => \N__13008\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__13012\,
            I => \N__13005\
        );

    \I__1391\ : InMux
    port map (
            O => \N__13011\,
            I => \N__13002\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__13008\,
            I => \eeprom.n3201\
        );

    \I__1389\ : Odrv4
    port map (
            O => \N__13005\,
            I => \eeprom.n3201\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__13002\,
            I => \eeprom.n3201\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__12995\,
            I => \N__12992\
        );

    \I__1386\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12989\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__12989\,
            I => \N__12985\
        );

    \I__1384\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12982\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__12985\,
            I => \eeprom.n3203\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__12982\,
            I => \eeprom.n3203\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__1380\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12970\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__12973\,
            I => \N__12967\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__12970\,
            I => \N__12964\
        );

    \I__1377\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12961\
        );

    \I__1376\ : Span4Mux_v
    port map (
            O => \N__12964\,
            I => \N__12958\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__12961\,
            I => \eeprom.n3200\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__12958\,
            I => \eeprom.n3200\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__12953\,
            I => \eeprom.n3200_cascade_\
        );

    \I__1372\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12947\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__12947\,
            I => \N__12944\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__12944\,
            I => \N__12941\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__12941\,
            I => \eeprom.n3286\
        );

    \I__1368\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12935\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__12935\,
            I => \N__12932\
        );

    \I__1366\ : Span4Mux_h
    port map (
            O => \N__12932\,
            I => \N__12929\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__12929\,
            I => \eeprom.n3280\
        );

    \I__1364\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12923\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__12923\,
            I => \N__12920\
        );

    \I__1362\ : Span4Mux_h
    port map (
            O => \N__12920\,
            I => \N__12917\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__12917\,
            I => \eeprom.n3275\
        );

    \I__1360\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12911\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__12908\,
            I => \N__12905\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__12905\,
            I => \eeprom.n3276\
        );

    \I__1356\ : InMux
    port map (
            O => \N__12902\,
            I => \N__12899\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__12899\,
            I => \N__12896\
        );

    \I__1354\ : Span4Mux_h
    port map (
            O => \N__12896\,
            I => \N__12893\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__12893\,
            I => \eeprom.n3279\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__12890\,
            I => \eeprom.n3204_cascade_\
        );

    \I__1351\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__12884\,
            I => \N__12881\
        );

    \I__1349\ : Span4Mux_v
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__12878\,
            I => \eeprom.n3267\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__12875\,
            I => \eeprom.n3299_cascade_\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__12872\,
            I => \N__12868\
        );

    \I__1345\ : InMux
    port map (
            O => \N__12871\,
            I => \N__12865\
        );

    \I__1344\ : InMux
    port map (
            O => \N__12868\,
            I => \N__12862\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__12865\,
            I => \N__12859\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__12862\,
            I => \N__12854\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__12859\,
            I => \N__12854\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__12854\,
            I => \eeprom.n3298\
        );

    \I__1339\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__12848\,
            I => \eeprom.n3379\
        );

    \I__1337\ : InMux
    port map (
            O => \N__12845\,
            I => \N__12841\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__12844\,
            I => \N__12838\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__12841\,
            I => \N__12835\
        );

    \I__1334\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12832\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__12835\,
            I => \N__12829\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__12832\,
            I => \eeprom.n3299\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__12829\,
            I => \eeprom.n3299\
        );

    \I__1330\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12821\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__12821\,
            I => \N__12818\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__12818\,
            I => \eeprom.n3366\
        );

    \I__1327\ : InMux
    port map (
            O => \N__12815\,
            I => \N__12812\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__12812\,
            I => \N__12809\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__12809\,
            I => \N__12806\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__12806\,
            I => \eeprom.n3269\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__1322\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12797\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__12797\,
            I => \N__12793\
        );

    \I__1320\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12790\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__12793\,
            I => \eeprom.n3301\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__12790\,
            I => \eeprom.n3301\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__12785\,
            I => \eeprom.n3301_cascade_\
        );

    \I__1316\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__12779\,
            I => \N__12776\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__12776\,
            I => \eeprom.n3368\
        );

    \I__1313\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__12767\,
            I => \eeprom.n3374\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__12764\,
            I => \N__12761\
        );

    \I__1309\ : InMux
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__12758\,
            I => \N__12754\
        );

    \I__1307\ : CascadeMux
    port map (
            O => \N__12757\,
            I => \N__12751\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__12754\,
            I => \N__12747\
        );

    \I__1305\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12744\
        );

    \I__1304\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12741\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__12747\,
            I => \eeprom.n3406\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__12744\,
            I => \eeprom.n3406\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__12741\,
            I => \eeprom.n3406\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__12734\,
            I => \N__12731\
        );

    \I__1299\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__1297\ : Odrv4
    port map (
            O => \N__12725\,
            I => \eeprom.n3370\
        );

    \I__1296\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__12719\,
            I => \N__12716\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__12713\,
            I => \eeprom.n3268\
        );

    \I__1292\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12707\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__12707\,
            I => \N__12702\
        );

    \I__1290\ : InMux
    port map (
            O => \N__12706\,
            I => \N__12697\
        );

    \I__1289\ : InMux
    port map (
            O => \N__12705\,
            I => \N__12697\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__12702\,
            I => \eeprom.n3300\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__12697\,
            I => \eeprom.n3300\
        );

    \I__1286\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12689\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__12689\,
            I => \N__12686\
        );

    \I__1284\ : Span4Mux_h
    port map (
            O => \N__12686\,
            I => \N__12683\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__12683\,
            I => \eeprom.n3376\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__12680\,
            I => \N__12677\
        );

    \I__1281\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__12674\,
            I => \N__12671\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__12668\,
            I => \eeprom.n3380\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__12665\,
            I => \N__12661\
        );

    \I__1276\ : InMux
    port map (
            O => \N__12664\,
            I => \N__12658\
        );

    \I__1275\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12655\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__12658\,
            I => \eeprom.n3412\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__12655\,
            I => \eeprom.n3412\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__12650\,
            I => \eeprom.n3412_cascade_\
        );

    \I__1271\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12644\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__12644\,
            I => \eeprom.n3479\
        );

    \I__1269\ : InMux
    port map (
            O => \N__12641\,
            I => \N__12638\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__12638\,
            I => \N__12635\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__12635\,
            I => \eeprom.n3375\
        );

    \I__1266\ : InMux
    port map (
            O => \N__12632\,
            I => \N__12629\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__12629\,
            I => \N__12626\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__12626\,
            I => \eeprom.n3378\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__12623\,
            I => \N__12619\
        );

    \I__1262\ : InMux
    port map (
            O => \N__12622\,
            I => \N__12616\
        );

    \I__1261\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12613\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__12616\,
            I => \eeprom.n3410\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__12613\,
            I => \eeprom.n3410\
        );

    \I__1258\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12605\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__12605\,
            I => \eeprom.n3477\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__12602\,
            I => \eeprom.n3410_cascade_\
        );

    \I__1255\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12596\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__12596\,
            I => \eeprom.n3465\
        );

    \I__1253\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12590\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__12590\,
            I => \N__12587\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__12587\,
            I => \N__12584\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__12584\,
            I => \eeprom.n3367\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__12581\,
            I => \eeprom.n3505_cascade_\
        );

    \I__1248\ : InMux
    port map (
            O => \N__12578\,
            I => \N__12575\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__12575\,
            I => \eeprom.n30_adj_273\
        );

    \I__1246\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12569\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__12569\,
            I => \eeprom.n3478\
        );

    \I__1244\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__12563\,
            I => \eeprom.n3472\
        );

    \I__1242\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12557\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__12557\,
            I => \eeprom.n3484\
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__12554\,
            I => \N__12551\
        );

    \I__1239\ : InMux
    port map (
            O => \N__12551\,
            I => \N__12548\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__12548\,
            I => \eeprom.n3475\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__12545\,
            I => \eeprom.n3507_cascade_\
        );

    \I__1236\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12539\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__12539\,
            I => \eeprom.n31\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__12536\,
            I => \N__12533\
        );

    \I__1233\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__12530\,
            I => \eeprom.n3482\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__12527\,
            I => \eeprom.n3514_cascade_\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__12524\,
            I => \eeprom.n5323_cascade_\
        );

    \I__1229\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12518\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__12518\,
            I => \eeprom.n5321\
        );

    \I__1227\ : InMux
    port map (
            O => \N__12515\,
            I => \N__12512\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__12512\,
            I => \eeprom.n4753\
        );

    \I__1225\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__12506\,
            I => \eeprom.n3605\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__1222\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12497\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__12497\,
            I => \N__12494\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__12494\,
            I => \N__12491\
        );

    \I__1219\ : Odrv4
    port map (
            O => \N__12491\,
            I => \eeprom.n3471\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__12488\,
            I => \eeprom.n32_cascade_\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__12485\,
            I => \eeprom.n3529_cascade_\
        );

    \I__1216\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12479\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__12479\,
            I => \eeprom.n3481\
        );

    \I__1214\ : CascadeMux
    port map (
            O => \N__12476\,
            I => \eeprom.n3513_cascade_\
        );

    \I__1213\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__12470\,
            I => \N__12467\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__12467\,
            I => \eeprom.n3473\
        );

    \I__1210\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12458\
        );

    \I__1209\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12458\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__12458\,
            I => \N__12454\
        );

    \I__1207\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12451\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__12454\,
            I => blink_counter_24
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__12451\,
            I => blink_counter_24
        );

    \I__1204\ : InMux
    port map (
            O => \N__12446\,
            I => \N__12439\
        );

    \I__1203\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12439\
        );

    \I__1202\ : InMux
    port map (
            O => \N__12444\,
            I => \N__12436\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__12439\,
            I => blink_counter_22
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__12436\,
            I => blink_counter_22
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__12431\,
            I => \N__12427\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__12430\,
            I => \N__12424\
        );

    \I__1197\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12418\
        );

    \I__1196\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12418\
        );

    \I__1195\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12415\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__12418\,
            I => blink_counter_23
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__12415\,
            I => blink_counter_23
        );

    \I__1192\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12403\
        );

    \I__1191\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12403\
        );

    \I__1190\ : InMux
    port map (
            O => \N__12408\,
            I => \N__12400\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__12403\,
            I => blink_counter_21
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__12400\,
            I => blink_counter_21
        );

    \I__1187\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__12389\,
            I => \N__12386\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__12386\,
            I => n5420
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__12383\,
            I => \N__12380\
        );

    \I__1182\ : InMux
    port map (
            O => \N__12380\,
            I => \N__12377\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__12377\,
            I => \eeprom.n1203\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__12374\,
            I => \eeprom.n3713_cascade_\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__12371\,
            I => \eeprom.n3618_cascade_\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__12368\,
            I => \eeprom.n3615_cascade_\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__12365\,
            I => \eeprom.n5221_cascade_\
        );

    \I__1176\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12359\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__12359\,
            I => \eeprom.n5225\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__12356\,
            I => \N__12353\
        );

    \I__1173\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12349\
        );

    \I__1172\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12345\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__12349\,
            I => \N__12342\
        );

    \I__1170\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12339\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__12345\,
            I => \eeprom.n3614\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__12342\,
            I => \eeprom.n3614\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__12339\,
            I => \eeprom.n3614\
        );

    \I__1166\ : InMux
    port map (
            O => \N__12332\,
            I => \eeprom.n3966\
        );

    \I__1165\ : InMux
    port map (
            O => \N__12329\,
            I => \eeprom.n3967\
        );

    \I__1164\ : InMux
    port map (
            O => \N__12326\,
            I => \eeprom.n3968\
        );

    \I__1163\ : InMux
    port map (
            O => \N__12323\,
            I => \eeprom.n3969\
        );

    \I__1162\ : InMux
    port map (
            O => \N__12320\,
            I => \eeprom.n3970\
        );

    \I__1161\ : InMux
    port map (
            O => \N__12317\,
            I => \eeprom.n3971\
        );

    \I__1160\ : InMux
    port map (
            O => \N__12314\,
            I => \eeprom.n3972\
        );

    \I__1159\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12308\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__12308\,
            I => \N__12305\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__12305\,
            I => \N__12302\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__12302\,
            I => n5421
        );

    \I__1155\ : InMux
    port map (
            O => \N__12299\,
            I => \eeprom.n4155\
        );

    \I__1154\ : InMux
    port map (
            O => \N__12296\,
            I => \eeprom.n4156\
        );

    \I__1153\ : InMux
    port map (
            O => \N__12293\,
            I => \bfn_17_29_0_\
        );

    \I__1152\ : InMux
    port map (
            O => \N__12290\,
            I => \eeprom.n4158\
        );

    \I__1151\ : InMux
    port map (
            O => \N__12287\,
            I => \eeprom.n4159\
        );

    \I__1150\ : InMux
    port map (
            O => \N__12284\,
            I => \eeprom.n4160\
        );

    \I__1149\ : InMux
    port map (
            O => \N__12281\,
            I => \eeprom.n4161\
        );

    \I__1148\ : InMux
    port map (
            O => \N__12278\,
            I => \bfn_18_17_0_\
        );

    \I__1147\ : InMux
    port map (
            O => \N__12275\,
            I => \eeprom.n4146\
        );

    \I__1146\ : InMux
    port map (
            O => \N__12272\,
            I => \eeprom.n4147\
        );

    \I__1145\ : InMux
    port map (
            O => \N__12269\,
            I => \eeprom.n4148\
        );

    \I__1144\ : InMux
    port map (
            O => \N__12266\,
            I => \bfn_17_28_0_\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__12263\,
            I => \N__12260\
        );

    \I__1142\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12257\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__12257\,
            I => \N__12254\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__12254\,
            I => \eeprom.n3277\
        );

    \I__1139\ : InMux
    port map (
            O => \N__12251\,
            I => \eeprom.n4150\
        );

    \I__1138\ : InMux
    port map (
            O => \N__12248\,
            I => \eeprom.n4151\
        );

    \I__1137\ : InMux
    port map (
            O => \N__12245\,
            I => \eeprom.n4152\
        );

    \I__1136\ : InMux
    port map (
            O => \N__12242\,
            I => \eeprom.n4153\
        );

    \I__1135\ : InMux
    port map (
            O => \N__12239\,
            I => \eeprom.n4154\
        );

    \I__1134\ : InMux
    port map (
            O => \N__12236\,
            I => \eeprom.n4179\
        );

    \I__1133\ : InMux
    port map (
            O => \N__12233\,
            I => \eeprom.n4180\
        );

    \I__1132\ : InMux
    port map (
            O => \N__12230\,
            I => \eeprom.n4181\
        );

    \I__1131\ : InMux
    port map (
            O => \N__12227\,
            I => \eeprom.n4182\
        );

    \I__1130\ : InMux
    port map (
            O => \N__12224\,
            I => \bfn_17_27_0_\
        );

    \I__1129\ : InMux
    port map (
            O => \N__12221\,
            I => \eeprom.n4142\
        );

    \I__1128\ : InMux
    port map (
            O => \N__12218\,
            I => \eeprom.n4143\
        );

    \I__1127\ : InMux
    port map (
            O => \N__12215\,
            I => \eeprom.n4144\
        );

    \I__1126\ : InMux
    port map (
            O => \N__12212\,
            I => \eeprom.n4145\
        );

    \I__1125\ : InMux
    port map (
            O => \N__12209\,
            I => \eeprom.n4170\
        );

    \I__1124\ : InMux
    port map (
            O => \N__12206\,
            I => \eeprom.n4171\
        );

    \I__1123\ : InMux
    port map (
            O => \N__12203\,
            I => \eeprom.n4172\
        );

    \I__1122\ : InMux
    port map (
            O => \N__12200\,
            I => \eeprom.n4173\
        );

    \I__1121\ : InMux
    port map (
            O => \N__12197\,
            I => \eeprom.n4174\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__12194\,
            I => \N__12191\
        );

    \I__1119\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12188\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__12188\,
            I => \N__12185\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__12185\,
            I => \eeprom.n3372\
        );

    \I__1116\ : InMux
    port map (
            O => \N__12182\,
            I => \eeprom.n4175\
        );

    \I__1115\ : InMux
    port map (
            O => \N__12179\,
            I => \eeprom.n4176\
        );

    \I__1114\ : InMux
    port map (
            O => \N__12176\,
            I => \bfn_17_26_0_\
        );

    \I__1113\ : InMux
    port map (
            O => \N__12173\,
            I => \eeprom.n4178\
        );

    \I__1112\ : InMux
    port map (
            O => \N__12170\,
            I => \bfn_17_24_0_\
        );

    \I__1111\ : InMux
    port map (
            O => \N__12167\,
            I => \eeprom.n4162\
        );

    \I__1110\ : InMux
    port map (
            O => \N__12164\,
            I => \eeprom.n4163\
        );

    \I__1109\ : InMux
    port map (
            O => \N__12161\,
            I => \eeprom.n4164\
        );

    \I__1108\ : InMux
    port map (
            O => \N__12158\,
            I => \eeprom.n4165\
        );

    \I__1107\ : InMux
    port map (
            O => \N__12155\,
            I => \eeprom.n4166\
        );

    \I__1106\ : InMux
    port map (
            O => \N__12152\,
            I => \eeprom.n4167\
        );

    \I__1105\ : InMux
    port map (
            O => \N__12149\,
            I => \eeprom.n4168\
        );

    \I__1104\ : InMux
    port map (
            O => \N__12146\,
            I => \bfn_17_25_0_\
        );

    \I__1103\ : InMux
    port map (
            O => \N__12143\,
            I => \eeprom.n4197\
        );

    \I__1102\ : InMux
    port map (
            O => \N__12140\,
            I => \bfn_17_23_0_\
        );

    \I__1101\ : InMux
    port map (
            O => \N__12137\,
            I => \eeprom.n4199\
        );

    \I__1100\ : InMux
    port map (
            O => \N__12134\,
            I => \eeprom.n4200\
        );

    \I__1099\ : InMux
    port map (
            O => \N__12131\,
            I => \eeprom.n4201\
        );

    \I__1098\ : InMux
    port map (
            O => \N__12128\,
            I => \eeprom.n4202\
        );

    \I__1097\ : InMux
    port map (
            O => \N__12125\,
            I => \eeprom.n4203\
        );

    \I__1096\ : InMux
    port map (
            O => \N__12122\,
            I => \eeprom.n4204\
        );

    \I__1095\ : InMux
    port map (
            O => \N__12119\,
            I => \eeprom.n4188\
        );

    \I__1094\ : InMux
    port map (
            O => \N__12116\,
            I => \eeprom.n4189\
        );

    \I__1093\ : InMux
    port map (
            O => \N__12113\,
            I => \bfn_17_22_0_\
        );

    \I__1092\ : InMux
    port map (
            O => \N__12110\,
            I => \eeprom.n4191\
        );

    \I__1091\ : InMux
    port map (
            O => \N__12107\,
            I => \eeprom.n4192\
        );

    \I__1090\ : InMux
    port map (
            O => \N__12104\,
            I => \eeprom.n4193\
        );

    \I__1089\ : InMux
    port map (
            O => \N__12101\,
            I => \eeprom.n4194\
        );

    \I__1088\ : InMux
    port map (
            O => \N__12098\,
            I => \eeprom.n4195\
        );

    \I__1087\ : InMux
    port map (
            O => \N__12095\,
            I => \eeprom.n4196\
        );

    \I__1086\ : InMux
    port map (
            O => \N__12092\,
            I => n3928
        );

    \I__1085\ : InMux
    port map (
            O => \N__12089\,
            I => \bfn_17_20_0_\
        );

    \I__1084\ : InMux
    port map (
            O => \N__12086\,
            I => n3930
        );

    \I__1083\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12080\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__12080\,
            I => \N__12077\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__12077\,
            I => \N__12073\
        );

    \I__1080\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12070\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__12073\,
            I => blink_counter_25
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__12070\,
            I => blink_counter_25
        );

    \I__1077\ : InMux
    port map (
            O => \N__12065\,
            I => \bfn_17_21_0_\
        );

    \I__1076\ : InMux
    port map (
            O => \N__12062\,
            I => \eeprom.n4183\
        );

    \I__1075\ : InMux
    port map (
            O => \N__12059\,
            I => \eeprom.n4184\
        );

    \I__1074\ : InMux
    port map (
            O => \N__12056\,
            I => \eeprom.n4185\
        );

    \I__1073\ : InMux
    port map (
            O => \N__12053\,
            I => \eeprom.n4186\
        );

    \I__1072\ : InMux
    port map (
            O => \N__12050\,
            I => \eeprom.n4187\
        );

    \I__1071\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12044\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__12044\,
            I => n12
        );

    \I__1069\ : InMux
    port map (
            O => \N__12041\,
            I => n3919
        );

    \I__1068\ : InMux
    port map (
            O => \N__12038\,
            I => \N__12035\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__12035\,
            I => n11_adj_364
        );

    \I__1066\ : InMux
    port map (
            O => \N__12032\,
            I => n3920
        );

    \I__1065\ : InMux
    port map (
            O => \N__12029\,
            I => \N__12026\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__12026\,
            I => n10_adj_363
        );

    \I__1063\ : InMux
    port map (
            O => \N__12023\,
            I => \bfn_17_19_0_\
        );

    \I__1062\ : InMux
    port map (
            O => \N__12020\,
            I => \N__12017\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__12017\,
            I => n9
        );

    \I__1060\ : InMux
    port map (
            O => \N__12014\,
            I => n3922
        );

    \I__1059\ : InMux
    port map (
            O => \N__12011\,
            I => \N__12008\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__12008\,
            I => n8_adj_362
        );

    \I__1057\ : InMux
    port map (
            O => \N__12005\,
            I => n3923
        );

    \I__1056\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11999\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__11999\,
            I => n7
        );

    \I__1054\ : InMux
    port map (
            O => \N__11996\,
            I => n3924
        );

    \I__1053\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11990\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__11990\,
            I => n6
        );

    \I__1051\ : InMux
    port map (
            O => \N__11987\,
            I => n3925
        );

    \I__1050\ : InMux
    port map (
            O => \N__11984\,
            I => n3926
        );

    \I__1049\ : InMux
    port map (
            O => \N__11981\,
            I => n3927
        );

    \I__1048\ : InMux
    port map (
            O => \N__11978\,
            I => \N__11975\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__11975\,
            I => n20
        );

    \I__1046\ : InMux
    port map (
            O => \N__11972\,
            I => n3911
        );

    \I__1045\ : InMux
    port map (
            O => \N__11969\,
            I => \N__11966\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__11966\,
            I => n19
        );

    \I__1043\ : InMux
    port map (
            O => \N__11963\,
            I => n3912
        );

    \I__1042\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__11957\,
            I => n18
        );

    \I__1040\ : InMux
    port map (
            O => \N__11954\,
            I => \bfn_17_18_0_\
        );

    \I__1039\ : InMux
    port map (
            O => \N__11951\,
            I => \N__11948\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__11948\,
            I => n17
        );

    \I__1037\ : InMux
    port map (
            O => \N__11945\,
            I => n3914
        );

    \I__1036\ : InMux
    port map (
            O => \N__11942\,
            I => \N__11939\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__11939\,
            I => n16
        );

    \I__1034\ : InMux
    port map (
            O => \N__11936\,
            I => n3915
        );

    \I__1033\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11930\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__11930\,
            I => n15
        );

    \I__1031\ : InMux
    port map (
            O => \N__11927\,
            I => n3916
        );

    \I__1030\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11921\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__11921\,
            I => n14
        );

    \I__1028\ : InMux
    port map (
            O => \N__11918\,
            I => n3917
        );

    \I__1027\ : InMux
    port map (
            O => \N__11915\,
            I => \N__11912\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__11912\,
            I => n13
        );

    \I__1025\ : InMux
    port map (
            O => \N__11909\,
            I => n3918
        );

    \I__1024\ : IoInMux
    port map (
            O => \N__11906\,
            I => \N__11903\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__11903\,
            I => \N__11900\
        );

    \I__1022\ : Span4Mux_s2_v
    port map (
            O => \N__11900\,
            I => \N__11897\
        );

    \I__1021\ : Sp12to4
    port map (
            O => \N__11897\,
            I => \N__11894\
        );

    \I__1020\ : Span12Mux_h
    port map (
            O => \N__11894\,
            I => \N__11891\
        );

    \I__1019\ : Odrv12
    port map (
            O => \N__11891\,
            I => \LED_c\
        );

    \I__1018\ : InMux
    port map (
            O => \N__11888\,
            I => \N__11885\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__11885\,
            I => n26
        );

    \I__1016\ : InMux
    port map (
            O => \N__11882\,
            I => \bfn_17_17_0_\
        );

    \I__1015\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__11876\,
            I => n25
        );

    \I__1013\ : InMux
    port map (
            O => \N__11873\,
            I => n3906
        );

    \I__1012\ : InMux
    port map (
            O => \N__11870\,
            I => \N__11867\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__11867\,
            I => n24
        );

    \I__1010\ : InMux
    port map (
            O => \N__11864\,
            I => n3907
        );

    \I__1009\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11858\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__11858\,
            I => n23
        );

    \I__1007\ : InMux
    port map (
            O => \N__11855\,
            I => n3908
        );

    \I__1006\ : InMux
    port map (
            O => \N__11852\,
            I => \N__11849\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__11849\,
            I => n22
        );

    \I__1004\ : InMux
    port map (
            O => \N__11846\,
            I => n3909
        );

    \I__1003\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11840\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__11840\,
            I => n21
        );

    \I__1001\ : InMux
    port map (
            O => \N__11837\,
            I => n3910
        );

    \I__1000\ : IoInMux
    port map (
            O => \N__11834\,
            I => \N__11831\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__11831\,
            I => \N__11828\
        );

    \I__998\ : IoSpan4Mux
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__997\ : IoSpan4Mux
    port map (
            O => \N__11825\,
            I => \N__11822\
        );

    \I__996\ : IoSpan4Mux
    port map (
            O => \N__11822\,
            I => \N__11819\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__11819\,
            I => \CLK_pad_gb_input\
        );

    \INVeeprom.i2c.write_enable_132C\ : INV
    port map (
            O => \INVeeprom.i2c.write_enable_132C_net\,
            I => \N__29683\
        );

    \INVeeprom.i2c.sda_out_133C\ : INV
    port map (
            O => \INVeeprom.i2c.sda_out_133C_net\,
            I => \N__29656\
        );

    \INVeeprom.i2c.i2c_scl_enable_124C\ : INV
    port map (
            O => \INVeeprom.i2c.i2c_scl_enable_124C_net\,
            I => \N__29696\
        );

    \IN_MUX_bfv_27_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_27_23_0_\
        );

    \IN_MUX_bfv_27_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4249\,
            carryinitout => \bfn_27_24_0_\
        );

    \IN_MUX_bfv_27_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4257\,
            carryinitout => \bfn_27_25_0_\
        );

    \IN_MUX_bfv_27_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4265\,
            carryinitout => \bfn_27_26_0_\
        );

    \IN_MUX_bfv_20_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_17_0_\
        );

    \IN_MUX_bfv_20_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4235\,
            carryinitout => \bfn_20_18_0_\
        );

    \IN_MUX_bfv_20_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_19_0_\
        );

    \IN_MUX_bfv_20_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4212\,
            carryinitout => \bfn_20_20_0_\
        );

    \IN_MUX_bfv_20_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4220\,
            carryinitout => \bfn_20_21_0_\
        );

    \IN_MUX_bfv_17_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_21_0_\
        );

    \IN_MUX_bfv_17_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4190\,
            carryinitout => \bfn_17_22_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4198\,
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_17_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4169\,
            carryinitout => \bfn_17_25_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4177\,
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_17_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_27_0_\
        );

    \IN_MUX_bfv_17_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4149\,
            carryinitout => \bfn_17_28_0_\
        );

    \IN_MUX_bfv_17_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4157\,
            carryinitout => \bfn_17_29_0_\
        );

    \IN_MUX_bfv_19_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_19_30_0_\
        );

    \IN_MUX_bfv_19_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4130\,
            carryinitout => \bfn_19_31_0_\
        );

    \IN_MUX_bfv_19_32_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4138\,
            carryinitout => \bfn_19_32_0_\
        );

    \IN_MUX_bfv_18_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_29_0_\
        );

    \IN_MUX_bfv_18_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4112\,
            carryinitout => \bfn_18_30_0_\
        );

    \IN_MUX_bfv_18_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4120\,
            carryinitout => \bfn_18_31_0_\
        );

    \IN_MUX_bfv_20_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_29_0_\
        );

    \IN_MUX_bfv_20_30_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4095\,
            carryinitout => \bfn_20_30_0_\
        );

    \IN_MUX_bfv_20_31_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4103\,
            carryinitout => \bfn_20_31_0_\
        );

    \IN_MUX_bfv_21_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_27_0_\
        );

    \IN_MUX_bfv_21_28_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4079\,
            carryinitout => \bfn_21_28_0_\
        );

    \IN_MUX_bfv_21_29_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4087\,
            carryinitout => \bfn_21_29_0_\
        );

    \IN_MUX_bfv_22_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_25_0_\
        );

    \IN_MUX_bfv_22_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4064\,
            carryinitout => \bfn_22_26_0_\
        );

    \IN_MUX_bfv_21_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_23_0_\
        );

    \IN_MUX_bfv_21_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4050\,
            carryinitout => \bfn_21_24_0_\
        );

    \IN_MUX_bfv_24_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_23_0_\
        );

    \IN_MUX_bfv_24_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4037\,
            carryinitout => \bfn_24_24_0_\
        );

    \IN_MUX_bfv_22_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_22_0_\
        );

    \IN_MUX_bfv_22_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4025\,
            carryinitout => \bfn_22_23_0_\
        );

    \IN_MUX_bfv_21_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_20_0_\
        );

    \IN_MUX_bfv_21_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4014\,
            carryinitout => \bfn_21_21_0_\
        );

    \IN_MUX_bfv_22_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_17_0_\
        );

    \IN_MUX_bfv_22_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n4004\,
            carryinitout => \bfn_22_18_0_\
        );

    \IN_MUX_bfv_24_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_17_0_\
        );

    \IN_MUX_bfv_24_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3995\,
            carryinitout => \bfn_24_18_0_\
        );

    \IN_MUX_bfv_23_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_23_18_0_\
        );

    \IN_MUX_bfv_23_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3987\,
            carryinitout => \bfn_23_19_0_\
        );

    \IN_MUX_bfv_24_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_24_20_0_\
        );

    \IN_MUX_bfv_27_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_27_17_0_\
        );

    \IN_MUX_bfv_30_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_30_20_0_\
        );

    \IN_MUX_bfv_26_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_26_21_0_\
        );

    \IN_MUX_bfv_26_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3938\,
            carryinitout => \bfn_26_22_0_\
        );

    \IN_MUX_bfv_26_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3946\,
            carryinitout => \bfn_26_23_0_\
        );

    \IN_MUX_bfv_26_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \eeprom.n3954\,
            carryinitout => \bfn_26_24_0_\
        );

    \IN_MUX_bfv_18_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_17_0_\
        );

    \IN_MUX_bfv_28_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_28_21_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3913,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3921,
            carryinitout => \bfn_17_19_0_\
        );

    \IN_MUX_bfv_17_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n3929,
            carryinitout => \bfn_17_20_0_\
        );

    \CLK_pad_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11834\,
            GLOBALBUFFEROUTPUT => \CLK_N\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i4592_3_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__12083\,
            in1 => \N__12395\,
            in2 => \_gnd_net_\,
            in3 => \N__12311\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i0_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11888\,
            in2 => \_gnd_net_\,
            in3 => \N__11882\,
            lcout => n26,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => n3906,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i1_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11879\,
            in2 => \_gnd_net_\,
            in3 => \N__11873\,
            lcout => n25,
            ltout => OPEN,
            carryin => n3906,
            carryout => n3907,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i2_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11870\,
            in2 => \_gnd_net_\,
            in3 => \N__11864\,
            lcout => n24,
            ltout => OPEN,
            carryin => n3907,
            carryout => n3908,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i3_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11861\,
            in2 => \_gnd_net_\,
            in3 => \N__11855\,
            lcout => n23,
            ltout => OPEN,
            carryin => n3908,
            carryout => n3909,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i4_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11852\,
            in2 => \_gnd_net_\,
            in3 => \N__11846\,
            lcout => n22,
            ltout => OPEN,
            carryin => n3909,
            carryout => n3910,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i5_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11843\,
            in2 => \_gnd_net_\,
            in3 => \N__11837\,
            lcout => n21,
            ltout => OPEN,
            carryin => n3910,
            carryout => n3911,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i6_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11978\,
            in2 => \_gnd_net_\,
            in3 => \N__11972\,
            lcout => n20,
            ltout => OPEN,
            carryin => n3911,
            carryout => n3912,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i7_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11969\,
            in2 => \_gnd_net_\,
            in3 => \N__11963\,
            lcout => n19,
            ltout => OPEN,
            carryin => n3912,
            carryout => n3913,
            clk => \N__29856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i8_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11960\,
            in2 => \_gnd_net_\,
            in3 => \N__11954\,
            lcout => n18,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => n3914,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i9_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11951\,
            in2 => \_gnd_net_\,
            in3 => \N__11945\,
            lcout => n17,
            ltout => OPEN,
            carryin => n3914,
            carryout => n3915,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i10_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11942\,
            in2 => \_gnd_net_\,
            in3 => \N__11936\,
            lcout => n16,
            ltout => OPEN,
            carryin => n3915,
            carryout => n3916,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i11_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11933\,
            in2 => \_gnd_net_\,
            in3 => \N__11927\,
            lcout => n15,
            ltout => OPEN,
            carryin => n3916,
            carryout => n3917,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i12_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11924\,
            in2 => \_gnd_net_\,
            in3 => \N__11918\,
            lcout => n14,
            ltout => OPEN,
            carryin => n3917,
            carryout => n3918,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i13_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11915\,
            in2 => \_gnd_net_\,
            in3 => \N__11909\,
            lcout => n13,
            ltout => OPEN,
            carryin => n3918,
            carryout => n3919,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i14_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12047\,
            in2 => \_gnd_net_\,
            in3 => \N__12041\,
            lcout => n12,
            ltout => OPEN,
            carryin => n3919,
            carryout => n3920,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i15_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12038\,
            in2 => \_gnd_net_\,
            in3 => \N__12032\,
            lcout => n11_adj_364,
            ltout => OPEN,
            carryin => n3920,
            carryout => n3921,
            clk => \N__29857\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i16_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12029\,
            in2 => \_gnd_net_\,
            in3 => \N__12023\,
            lcout => n10_adj_363,
            ltout => OPEN,
            carryin => \bfn_17_19_0_\,
            carryout => n3922,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i17_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12020\,
            in2 => \_gnd_net_\,
            in3 => \N__12014\,
            lcout => n9,
            ltout => OPEN,
            carryin => n3922,
            carryout => n3923,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i18_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12011\,
            in2 => \_gnd_net_\,
            in3 => \N__12005\,
            lcout => n8_adj_362,
            ltout => OPEN,
            carryin => n3923,
            carryout => n3924,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i19_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12002\,
            in2 => \_gnd_net_\,
            in3 => \N__11996\,
            lcout => n7,
            ltout => OPEN,
            carryin => n3924,
            carryout => n3925,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i20_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11993\,
            in2 => \_gnd_net_\,
            in3 => \N__11987\,
            lcout => n6,
            ltout => OPEN,
            carryin => n3925,
            carryout => n3926,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i21_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12408\,
            in2 => \_gnd_net_\,
            in3 => \N__11984\,
            lcout => blink_counter_21,
            ltout => OPEN,
            carryin => n3926,
            carryout => n3927,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i22_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12444\,
            in2 => \_gnd_net_\,
            in3 => \N__11981\,
            lcout => blink_counter_22,
            ltout => OPEN,
            carryin => n3927,
            carryout => n3928,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i23_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12423\,
            in2 => \_gnd_net_\,
            in3 => \N__12092\,
            lcout => blink_counter_23,
            ltout => OPEN,
            carryin => n3928,
            carryout => n3929,
            clk => \N__29858\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i24_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12457\,
            in2 => \_gnd_net_\,
            in3 => \N__12089\,
            lcout => blink_counter_24,
            ltout => OPEN,
            carryin => \bfn_17_20_0_\,
            carryout => n3930,
            clk => \N__29859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \blink_counter_227__i25_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12076\,
            in2 => \_gnd_net_\,
            in3 => \N__12086\,
            lcout => blink_counter_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29859\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_2_lut_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23421\,
            in2 => \_gnd_net_\,
            in3 => \N__12065\,
            lcout => \eeprom.n3486\,
            ltout => OPEN,
            carryin => \bfn_17_21_0_\,
            carryout => \eeprom.n4183\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_3_lut_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28538\,
            in2 => \N__16664\,
            in3 => \N__12062\,
            lcout => \eeprom.n3485\,
            ltout => OPEN,
            carryin => \eeprom.n4183\,
            carryout => \eeprom.n4184\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_4_lut_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16166\,
            in3 => \N__12059\,
            lcout => \eeprom.n3484\,
            ltout => OPEN,
            carryin => \eeprom.n4184\,
            carryout => \eeprom.n4185\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_5_lut_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16625\,
            in3 => \N__12056\,
            lcout => \eeprom.n3483\,
            ltout => OPEN,
            carryin => \eeprom.n4185\,
            carryout => \eeprom.n4186\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_6_lut_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17228\,
            in3 => \N__12053\,
            lcout => \eeprom.n3482\,
            ltout => OPEN,
            carryin => \eeprom.n4186\,
            carryout => \eeprom.n4187\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_7_lut_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16183\,
            in2 => \_gnd_net_\,
            in3 => \N__12050\,
            lcout => \eeprom.n3481\,
            ltout => OPEN,
            carryin => \eeprom.n4187\,
            carryout => \eeprom.n4188\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_8_lut_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16511\,
            in3 => \N__12119\,
            lcout => \eeprom.n3480\,
            ltout => OPEN,
            carryin => \eeprom.n4188\,
            carryout => \eeprom.n4189\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_9_lut_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28539\,
            in2 => \N__12665\,
            in3 => \N__12116\,
            lcout => \eeprom.n3479\,
            ltout => OPEN,
            carryin => \eeprom.n4189\,
            carryout => \eeprom.n4190\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_10_lut_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28764\,
            in2 => \N__13759\,
            in3 => \N__12113\,
            lcout => \eeprom.n3478\,
            ltout => OPEN,
            carryin => \bfn_17_22_0_\,
            carryout => \eeprom.n4191\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_11_lut_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28768\,
            in2 => \N__12623\,
            in3 => \N__12110\,
            lcout => \eeprom.n3477\,
            ltout => OPEN,
            carryin => \eeprom.n4191\,
            carryout => \eeprom.n4192\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_12_lut_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28765\,
            in2 => \N__17033\,
            in3 => \N__12107\,
            lcout => \eeprom.n3476\,
            ltout => OPEN,
            carryin => \eeprom.n4192\,
            carryout => \eeprom.n4193\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_13_lut_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28769\,
            in2 => \N__13781\,
            in3 => \N__12104\,
            lcout => \eeprom.n3475\,
            ltout => OPEN,
            carryin => \eeprom.n4193\,
            carryout => \eeprom.n4194\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_14_lut_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28766\,
            in2 => \N__13510\,
            in3 => \N__12101\,
            lcout => \eeprom.n3474\,
            ltout => OPEN,
            carryin => \eeprom.n4194\,
            carryout => \eeprom.n4195\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_15_lut_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28770\,
            in2 => \N__12757\,
            in3 => \N__12098\,
            lcout => \eeprom.n3473\,
            ltout => OPEN,
            carryin => \eeprom.n4195\,
            carryout => \eeprom.n4196\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_16_lut_LC_17_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28767\,
            in2 => \N__16751\,
            in3 => \N__12095\,
            lcout => \eeprom.n3472\,
            ltout => OPEN,
            carryin => \eeprom.n4196\,
            carryout => \eeprom.n4197\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_17_lut_LC_17_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28771\,
            in2 => \N__16710\,
            in3 => \N__12143\,
            lcout => \eeprom.n3471\,
            ltout => OPEN,
            carryin => \eeprom.n4197\,
            carryout => \eeprom.n4198\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_18_lut_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28772\,
            in2 => \N__19262\,
            in3 => \N__12140\,
            lcout => \eeprom.n3470\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \eeprom.n4199\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_19_lut_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28777\,
            in2 => \N__14006\,
            in3 => \N__12137\,
            lcout => \eeprom.n3469\,
            ltout => OPEN,
            carryin => \eeprom.n4199\,
            carryout => \eeprom.n4200\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_20_lut_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14074\,
            in2 => \N__28874\,
            in3 => \N__12134\,
            lcout => \eeprom.n3468\,
            ltout => OPEN,
            carryin => \eeprom.n4200\,
            carryout => \eeprom.n4201\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_21_lut_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28781\,
            in2 => \N__14057\,
            in3 => \N__12131\,
            lcout => \eeprom.n3467\,
            ltout => OPEN,
            carryin => \eeprom.n4201\,
            carryout => \eeprom.n4202\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_22_lut_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28773\,
            in2 => \N__14036\,
            in3 => \N__12128\,
            lcout => \eeprom.n3466\,
            ltout => OPEN,
            carryin => \eeprom.n4202\,
            carryout => \eeprom.n4203\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_23_lut_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13818\,
            in2 => \N__28873\,
            in3 => \N__12125\,
            lcout => \eeprom.n3465\,
            ltout => OPEN,
            carryin => \eeprom.n4203\,
            carryout => \eeprom.n4204\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2290_24_lut_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28782\,
            in1 => \N__13798\,
            in2 => \N__19223\,
            in3 => \N__12122\,
            lcout => \eeprom.n3496\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2232_3_lut_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14195\,
            in2 => \N__12194\,
            in3 => \N__17155\,
            lcout => \eeprom.n3404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_2_lut_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22659\,
            in2 => \_gnd_net_\,
            in3 => \N__12170\,
            lcout => \eeprom.n3386\,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => \eeprom.n4162\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_3_lut_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28783\,
            in2 => \N__16880\,
            in3 => \N__12167\,
            lcout => \eeprom.n3385\,
            ltout => OPEN,
            carryin => \eeprom.n4162\,
            carryout => \eeprom.n4163\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_4_lut_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16951\,
            in2 => \_gnd_net_\,
            in3 => \N__12164\,
            lcout => \eeprom.n3384\,
            ltout => OPEN,
            carryin => \eeprom.n4163\,
            carryout => \eeprom.n4164\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_5_lut_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16910\,
            in3 => \N__12161\,
            lcout => \eeprom.n3383\,
            ltout => OPEN,
            carryin => \eeprom.n4164\,
            carryout => \eeprom.n4165\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_6_lut_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17660\,
            in3 => \N__12158\,
            lcout => \eeprom.n3382\,
            ltout => OPEN,
            carryin => \eeprom.n4165\,
            carryout => \eeprom.n4166\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_7_lut_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16934\,
            in3 => \N__12155\,
            lcout => \eeprom.n3381\,
            ltout => OPEN,
            carryin => \eeprom.n4166\,
            carryout => \eeprom.n4167\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_8_lut_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16583\,
            in3 => \N__12152\,
            lcout => \eeprom.n3380\,
            ltout => OPEN,
            carryin => \eeprom.n4167\,
            carryout => \eeprom.n4168\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_9_lut_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28784\,
            in2 => \N__13923\,
            in3 => \N__12149\,
            lcout => \eeprom.n3379\,
            ltout => OPEN,
            carryin => \eeprom.n4168\,
            carryout => \eeprom.n4169\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_10_lut_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28875\,
            in2 => \N__13951\,
            in3 => \N__12146\,
            lcout => \eeprom.n3378\,
            ltout => OPEN,
            carryin => \bfn_17_25_0_\,
            carryout => \eeprom.n4170\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_11_lut_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28878\,
            in2 => \N__17180\,
            in3 => \N__12209\,
            lcout => \eeprom.n3377\,
            ltout => OPEN,
            carryin => \eeprom.n4170\,
            carryout => \eeprom.n4171\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_12_lut_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13890\,
            in2 => \N__28928\,
            in3 => \N__12206\,
            lcout => \eeprom.n3376\,
            ltout => OPEN,
            carryin => \eeprom.n4171\,
            carryout => \eeprom.n4172\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_13_lut_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28882\,
            in2 => \N__14164\,
            in3 => \N__12203\,
            lcout => \eeprom.n3375\,
            ltout => OPEN,
            carryin => \eeprom.n4172\,
            carryout => \eeprom.n4173\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_14_lut_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28876\,
            in2 => \N__13975\,
            in3 => \N__12200\,
            lcout => \eeprom.n3374\,
            ltout => OPEN,
            carryin => \eeprom.n4173\,
            carryout => \eeprom.n4174\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_15_lut_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28883\,
            in2 => \N__14216\,
            in3 => \N__12197\,
            lcout => \eeprom.n3373\,
            ltout => OPEN,
            carryin => \eeprom.n4174\,
            carryout => \eeprom.n4175\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_16_lut_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28877\,
            in2 => \N__14194\,
            in3 => \N__12182\,
            lcout => \eeprom.n3372\,
            ltout => OPEN,
            carryin => \eeprom.n4175\,
            carryout => \eeprom.n4176\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_17_lut_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28884\,
            in2 => \N__16820\,
            in3 => \N__12179\,
            lcout => \eeprom.n3371\,
            ltout => OPEN,
            carryin => \eeprom.n4176\,
            carryout => \eeprom.n4177\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_18_lut_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28365\,
            in2 => \N__16847\,
            in3 => \N__12176\,
            lcout => \eeprom.n3370\,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => \eeprom.n4178\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_19_lut_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28885\,
            in2 => \N__16785\,
            in3 => \N__12173\,
            lcout => \eeprom.n3369\,
            ltout => OPEN,
            carryin => \eeprom.n4178\,
            carryout => \eeprom.n4179\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_20_lut_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28366\,
            in2 => \N__12803\,
            in3 => \N__12236\,
            lcout => \eeprom.n3368\,
            ltout => OPEN,
            carryin => \eeprom.n4179\,
            carryout => \eeprom.n4180\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_21_lut_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12710\,
            in2 => \N__28543\,
            in3 => \N__12233\,
            lcout => \eeprom.n3367\,
            ltout => OPEN,
            carryin => \eeprom.n4180\,
            carryout => \eeprom.n4181\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_22_lut_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12845\,
            in2 => \N__28929\,
            in3 => \N__12230\,
            lcout => \eeprom.n3366\,
            ltout => OPEN,
            carryin => \eeprom.n4181\,
            carryout => \eeprom.n4182\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2223_23_lut_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__28370\,
            in1 => \N__17159\,
            in2 => \N__12872\,
            in3 => \N__12227\,
            lcout => \eeprom.n3397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2169_3_lut_LC_17_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18186\,
            in2 => \N__12263\,
            in3 => \N__17782\,
            lcout => \eeprom.n3309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_2_lut_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24231\,
            in2 => \_gnd_net_\,
            in3 => \N__12224\,
            lcout => \eeprom.n3286\,
            ltout => OPEN,
            carryin => \bfn_17_27_0_\,
            carryout => \eeprom.n4142\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_3_lut_LC_17_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28371\,
            in2 => \N__16989\,
            in3 => \N__12221\,
            lcout => \eeprom.n3285\,
            ltout => OPEN,
            carryin => \eeprom.n4142\,
            carryout => \eeprom.n4143\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_4_lut_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17327\,
            in3 => \N__12218\,
            lcout => \eeprom.n3284\,
            ltout => OPEN,
            carryin => \eeprom.n4143\,
            carryout => \eeprom.n4144\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_5_lut_LC_17_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17495\,
            in3 => \N__12215\,
            lcout => \eeprom.n3283\,
            ltout => OPEN,
            carryin => \eeprom.n4144\,
            carryout => \eeprom.n4145\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_6_lut_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17402\,
            in3 => \N__12212\,
            lcout => \eeprom.n3282\,
            ltout => OPEN,
            carryin => \eeprom.n4145\,
            carryout => \eeprom.n4146\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_7_lut_LC_17_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17513\,
            in2 => \_gnd_net_\,
            in3 => \N__12275\,
            lcout => \eeprom.n3281\,
            ltout => OPEN,
            carryin => \eeprom.n4146\,
            carryout => \eeprom.n4147\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_8_lut_LC_17_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17584\,
            in2 => \_gnd_net_\,
            in3 => \N__12272\,
            lcout => \eeprom.n3280\,
            ltout => OPEN,
            carryin => \eeprom.n4147\,
            carryout => \eeprom.n4148\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_9_lut_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14259\,
            in2 => \N__28544\,
            in3 => \N__12269\,
            lcout => \eeprom.n3279\,
            ltout => OPEN,
            carryin => \eeprom.n4148\,
            carryout => \eeprom.n4149\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_10_lut_LC_17_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18224\,
            in2 => \N__28930\,
            in3 => \N__12266\,
            lcout => \eeprom.n3278\,
            ltout => OPEN,
            carryin => \bfn_17_28_0_\,
            carryout => \eeprom.n4150\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_11_lut_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28892\,
            in2 => \N__18194\,
            in3 => \N__12251\,
            lcout => \eeprom.n3277\,
            ltout => OPEN,
            carryin => \eeprom.n4150\,
            carryout => \eeprom.n4151\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_12_lut_LC_17_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28375\,
            in2 => \N__17836\,
            in3 => \N__12248\,
            lcout => \eeprom.n3276\,
            ltout => OPEN,
            carryin => \eeprom.n4151\,
            carryout => \eeprom.n4152\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_13_lut_LC_17_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17251\,
            in2 => \N__28545\,
            in3 => \N__12245\,
            lcout => \eeprom.n3275\,
            ltout => OPEN,
            carryin => \eeprom.n4152\,
            carryout => \eeprom.n4153\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_14_lut_LC_17_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28379\,
            in2 => \N__14366\,
            in3 => \N__12242\,
            lcout => \eeprom.n3274\,
            ltout => OPEN,
            carryin => \eeprom.n4153\,
            carryout => \eeprom.n4154\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_15_lut_LC_17_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14288\,
            in2 => \N__28546\,
            in3 => \N__12239\,
            lcout => \eeprom.n3273\,
            ltout => OPEN,
            carryin => \eeprom.n4154\,
            carryout => \eeprom.n4155\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_16_lut_LC_17_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14426\,
            in2 => \N__28931\,
            in3 => \N__12299\,
            lcout => \eeprom.n3272\,
            ltout => OPEN,
            carryin => \eeprom.n4155\,
            carryout => \eeprom.n4156\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_17_lut_LC_17_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14393\,
            in2 => \N__28547\,
            in3 => \N__12296\,
            lcout => \eeprom.n3271\,
            ltout => OPEN,
            carryin => \eeprom.n4156\,
            carryout => \eeprom.n4157\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_18_lut_LC_17_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28386\,
            in2 => \N__12995\,
            in3 => \N__12293\,
            lcout => \eeprom.n3270\,
            ltout => OPEN,
            carryin => \bfn_17_29_0_\,
            carryout => \eeprom.n4158\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_19_lut_LC_17_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13048\,
            in2 => \N__28548\,
            in3 => \N__12290\,
            lcout => \eeprom.n3269\,
            ltout => OPEN,
            carryin => \eeprom.n4158\,
            carryout => \eeprom.n4159\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_20_lut_LC_17_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28390\,
            in2 => \N__13022\,
            in3 => \N__12287\,
            lcout => \eeprom.n3268\,
            ltout => OPEN,
            carryin => \eeprom.n4159\,
            carryout => \eeprom.n4160\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_21_lut_LC_17_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28391\,
            in2 => \N__12977\,
            in3 => \N__12284\,
            lcout => \eeprom.n3267\,
            ltout => OPEN,
            carryin => \eeprom.n4160\,
            carryout => \eeprom.n4161\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2156_22_lut_LC_17_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28392\,
            in1 => \N__15082\,
            in2 => \N__17786\,
            in3 => \N__12281\,
            lcout => \eeprom.n3298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1960_3_lut_LC_17_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19748\,
            in2 => \N__18824\,
            in3 => \N__18779\,
            lcout => \eeprom.n3004\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_2_lut_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21577\,
            in2 => \_gnd_net_\,
            in3 => \N__12278\,
            lcout => \eeprom.n1208\,
            ltout => OPEN,
            carryin => \bfn_18_17_0_\,
            carryout => \eeprom.n3966\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_3_lut_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13378\,
            in2 => \N__28537\,
            in3 => \N__12332\,
            lcout => \eeprom.n1207\,
            ltout => OPEN,
            carryin => \eeprom.n3966\,
            carryout => \eeprom.n3967\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_4_lut_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13568\,
            in3 => \N__12329\,
            lcout => \eeprom.n1206\,
            ltout => OPEN,
            carryin => \eeprom.n3967\,
            carryout => \eeprom.n3968\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_5_lut_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13340\,
            in3 => \N__12326\,
            lcout => \eeprom.n1205\,
            ltout => OPEN,
            carryin => \eeprom.n3968\,
            carryout => \eeprom.n3969\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_6_lut_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13478\,
            in2 => \_gnd_net_\,
            in3 => \N__12323\,
            lcout => \eeprom.n1204\,
            ltout => OPEN,
            carryin => \eeprom.n3969\,
            carryout => \eeprom.n3970\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_7_lut_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12356\,
            in3 => \N__12320\,
            lcout => \eeprom.n1203\,
            ltout => OPEN,
            carryin => \eeprom.n3970\,
            carryout => \eeprom.n3971\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_8_lut_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13225\,
            in2 => \_gnd_net_\,
            in3 => \N__12317\,
            lcout => \eeprom.n1202\,
            ltout => OPEN,
            carryin => \eeprom.n3971\,
            carryout => \eeprom.n3972\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_823_9_lut_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__28356\,
            in1 => \N__13583\,
            in2 => \_gnd_net_\,
            in3 => \N__12314\,
            lcout => \eeprom.n1201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4591_4_lut_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010110000"
        )
    port map (
            in0 => \N__12464\,
            in1 => \N__12446\,
            in2 => \N__12431\,
            in3 => \N__12410\,
            lcout => n5421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4738_1_lut_2_lut_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13451\,
            in3 => \N__13435\,
            lcout => \eeprom.n5568\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4590_4_lut_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101000000"
        )
    port map (
            in0 => \N__12463\,
            in1 => \N__12445\,
            in2 => \N__12430\,
            in3 => \N__12409\,
            lcout => n5420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2445_3_lut_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12352\,
            in2 => \N__12383\,
            in3 => \N__13434\,
            lcout => \eeprom.n3713\,
            ltout => \eeprom.n3713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4732_1_lut_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12374\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2382_3_lut_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15485\,
            in1 => \N__29459\,
            in2 => \_gnd_net_\,
            in3 => \N__16328\,
            lcout => \eeprom.n3618\,
            ltout => \eeprom.n3618_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_100_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__21576\,
            in1 => \N__12509\,
            in2 => \N__12371\,
            in3 => \N__12362\,
            lcout => \eeprom.n5017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2379_3_lut_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15854\,
            in2 => \N__16323\,
            in3 => \N__15880\,
            lcout => \eeprom.n3615\,
            ltout => \eeprom.n3615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_89_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12368\,
            in3 => \N__13218\,
            lcout => OPEN,
            ltout => \eeprom.n5221_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_99_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12348\,
            in1 => \N__13557\,
            in2 => \N__12365\,
            in3 => \N__13329\,
            lcout => \eeprom.n5225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2378_3_lut_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15841\,
            in2 => \N__15815\,
            in3 => \N__16300\,
            lcout => \eeprom.n3614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2369_3_lut_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__16064\,
            in1 => \_gnd_net_\,
            in2 => \N__16324\,
            in3 => \N__16046\,
            lcout => \eeprom.n3605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2380_3_lut_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15436\,
            in2 => \N__15410\,
            in3 => \N__16301\,
            lcout => \eeprom.n3616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2299_3_lut_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16715\,
            in2 => \N__12503\,
            in3 => \N__19221\,
            lcout => \eeprom.n3503\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i14_3_lut_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__16129\,
            in1 => \_gnd_net_\,
            in2 => \N__13694\,
            in3 => \N__16062\,
            lcout => OPEN,
            ltout => \eeprom.n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i17_4_lut_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12542\,
            in1 => \N__12578\,
            in2 => \N__12488\,
            in3 => \N__13589\,
            lcout => \eeprom.n3529\,
            ltout => \eeprom.n3529_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2377_3_lut_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15793\,
            in2 => \N__12485\,
            in3 => \N__15779\,
            lcout => \eeprom.n3613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2309_3_lut_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__12482\,
            in1 => \_gnd_net_\,
            in2 => \N__16187\,
            in3 => \N__19194\,
            lcout => \eeprom.n3513\,
            ltout => \eeprom.n3513_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_19_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12476\,
            in3 => \N__15831\,
            lcout => \eeprom.n5321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2301_3_lut_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12473\,
            in2 => \N__12764\,
            in3 => \N__19195\,
            lcout => \eeprom.n3505\,
            ltout => \eeprom.n3505_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_22_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15727\,
            in1 => \N__15993\,
            in2 => \N__12581\,
            in3 => \N__12515\,
            lcout => \eeprom.n30_adj_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4682_3_lut_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12572\,
            in2 => \N__19206\,
            in3 => \N__13760\,
            lcout => \eeprom.n3510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2300_3_lut_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12566\,
            in2 => \N__16750\,
            in3 => \N__19172\,
            lcout => \eeprom.n3504\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2312_3_lut_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16165\,
            in2 => \N__19205\,
            in3 => \N__12560\,
            lcout => \eeprom.n3516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2303_3_lut_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13780\,
            in2 => \N__12554\,
            in3 => \N__19173\,
            lcout => \eeprom.n3507\,
            ltout => \eeprom.n3507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_adj_23_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15690\,
            in1 => \N__15609\,
            in2 => \N__12545\,
            in3 => \N__15654\,
            lcout => \eeprom.n31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2310_3_lut_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17227\,
            in2 => \N__12536\,
            in3 => \N__19168\,
            lcout => \eeprom.n3514\,
            ltout => \eeprom.n3514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_20_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__15870\,
            in1 => \_gnd_net_\,
            in2 => \N__12527\,
            in3 => \N__15426\,
            lcout => OPEN,
            ltout => \eeprom.n5323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_21_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__29457\,
            in1 => \N__15465\,
            in2 => \N__12524\,
            in3 => \N__12521\,
            lcout => \eeprom.n4753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12664\,
            in1 => \N__12750\,
            in2 => \N__13509\,
            in3 => \N__12622\,
            lcout => \eeprom.n29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2236_3_lut_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13898\,
            in2 => \N__17157\,
            in3 => \N__12692\,
            lcout => \eeprom.n3408\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2240_3_lut_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16582\,
            in2 => \N__12680\,
            in3 => \N__17132\,
            lcout => \eeprom.n3412\,
            ltout => \eeprom.n3412_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2307_3_lut_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19188\,
            in1 => \_gnd_net_\,
            in2 => \N__12650\,
            in3 => \N__12647\,
            lcout => \eeprom.n3511\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2235_3_lut_LC_18_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__12641\,
            in1 => \_gnd_net_\,
            in2 => \N__14168\,
            in3 => \N__17136\,
            lcout => \eeprom.n3407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2238_3_lut_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12632\,
            in1 => \_gnd_net_\,
            in2 => \N__17156\,
            in3 => \N__13952\,
            lcout => \eeprom.n3410\,
            ltout => \eeprom.n3410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2305_3_lut_LC_18_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12608\,
            in2 => \N__12602\,
            in3 => \N__19189\,
            lcout => \eeprom.n3509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2293_3_lut_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__13819\,
            in1 => \_gnd_net_\,
            in2 => \N__19215\,
            in3 => \N__12599\,
            lcout => \eeprom.n3497\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2227_3_lut_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12706\,
            in2 => \N__17158\,
            in3 => \N__12593\,
            lcout => \eeprom.n3399\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2159_3_lut_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12887\,
            in2 => \N__12973\,
            in3 => \N__17764\,
            lcout => \eeprom.n3299\,
            ltout => \eeprom.n3299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_LC_18_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12796\,
            in1 => \N__12705\,
            in2 => \N__12875\,
            in3 => \N__12871\,
            lcout => \eeprom.n25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4681_3_lut_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12851\,
            in2 => \N__13925\,
            in3 => \N__17140\,
            lcout => \eeprom.n3411\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2226_3_lut_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17146\,
            in1 => \_gnd_net_\,
            in2 => \N__12844\,
            in3 => \N__12824\,
            lcout => \eeprom.n3398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2161_3_lut_LC_18_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__12815\,
            in1 => \_gnd_net_\,
            in2 => \N__13052\,
            in3 => \N__17763\,
            lcout => \eeprom.n3301\,
            ltout => \eeprom.n3301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2228_3_lut_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17145\,
            in1 => \_gnd_net_\,
            in2 => \N__12785\,
            in3 => \N__12782\,
            lcout => \eeprom.n3400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2234_3_lut_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12773\,
            in2 => \N__13976\,
            in3 => \N__17141\,
            lcout => \eeprom.n3406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2230_3_lut_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16840\,
            in2 => \N__12734\,
            in3 => \N__17149\,
            lcout => \eeprom.n3402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2160_3_lut_LC_18_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12722\,
            in2 => \N__17775\,
            in3 => \N__13021\,
            lcout => \eeprom.n3300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2092_3_lut_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15151\,
            in2 => \N__15125\,
            in3 => \N__17947\,
            lcout => \eeprom.n3200\,
            ltout => \eeprom.n3200_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_38_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12953\,
            in3 => \N__15083\,
            lcout => \eeprom.n16_adj_303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2178_3_lut_LC_18_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12950\,
            in1 => \N__24235\,
            in2 => \_gnd_net_\,
            in3 => \N__17744\,
            lcout => \eeprom.n3318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2172_rep_14_3_lut_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12938\,
            in2 => \N__17774\,
            in3 => \N__17585\,
            lcout => \eeprom.n3312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2167_3_lut_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__17252\,
            in1 => \_gnd_net_\,
            in2 => \N__17776\,
            in3 => \N__12926\,
            lcout => \eeprom.n3307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2168_3_lut_LC_18_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17837\,
            in2 => \N__17777\,
            in3 => \N__12914\,
            lcout => \eeprom.n3308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2171_3_lut_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12902\,
            in2 => \N__14264\,
            in3 => \N__17758\,
            lcout => \eeprom.n3311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2096_3_lut_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15290\,
            in2 => \N__15323\,
            in3 => \N__17946\,
            lcout => \eeprom.n3204\,
            ltout => \eeprom.n3204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_adj_39_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12988\,
            in1 => \N__13035\,
            in2 => \N__12890\,
            in3 => \N__13011\,
            lcout => \eeprom.n24_adj_304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2098_3_lut_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17945\,
            in2 => \N__14915\,
            in3 => \N__14891\,
            lcout => \eeprom.n3206\,
            ltout => \eeprom.n3206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2165_3_lut_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13067\,
            in2 => \N__13058\,
            in3 => \N__17754\,
            lcout => \eeprom.n3305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2032_3_lut_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13139\,
            in2 => \N__14314\,
            in3 => \N__18146\,
            lcout => \eeprom.n3108\,
            ltout => \eeprom.n3108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17292\,
            in1 => \N__14997\,
            in2 => \N__13055\,
            in3 => \N__14910\,
            lcout => \eeprom.n24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i8_4_lut_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15183\,
            in1 => \N__15141\,
            in2 => \N__15104\,
            in3 => \N__15226\,
            lcout => \eeprom.n22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2094_3_lut_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17933\,
            in2 => \N__15230\,
            in3 => \N__15206\,
            lcout => \eeprom.n3202\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2093_3_lut_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17934\,
            in1 => \_gnd_net_\,
            in2 => \N__15170\,
            in3 => \N__15184\,
            lcout => \eeprom.n3201\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2110_3_lut_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14795\,
            in1 => \N__22407\,
            in2 => \_gnd_net_\,
            in3 => \N__17926\,
            lcout => \eeprom.n3218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2095_3_lut_LC_18_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15245\,
            in2 => \N__17953\,
            in3 => \N__15275\,
            lcout => \eeprom.n3203\,
            ltout => \eeprom.n3203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2162_3_lut_LC_18_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13085\,
            in2 => \N__13076\,
            in3 => \N__17772\,
            lcout => \eeprom.n3302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2102_3_lut_LC_18_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14998\,
            in2 => \N__17952\,
            in3 => \N__14975\,
            lcout => \eeprom.n3210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2025_3_lut_LC_18_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14560\,
            in2 => \N__13277\,
            in3 => \N__18124\,
            lcout => \eeprom.n3101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2104_3_lut_LC_18_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15049\,
            in2 => \N__15035\,
            in3 => \N__17954\,
            lcout => \eeprom.n3212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2040_3_lut_LC_18_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14335\,
            in2 => \N__13100\,
            in3 => \N__18119\,
            lcout => \eeprom.n3116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2037_3_lut_LC_18_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13181\,
            in2 => \N__14452\,
            in3 => \N__18120\,
            lcout => \eeprom.n3113\,
            ltout => \eeprom.n3113_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_13_LC_18_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13073\,
            in3 => \N__17529\,
            lcout => OPEN,
            ltout => \eeprom.n5305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_14_LC_18_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14763\,
            in1 => \N__17616\,
            in2 => \N__13070\,
            in3 => \N__17433\,
            lcout => \eeprom.n5309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2026_3_lut_LC_18_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13292\,
            in2 => \N__18142\,
            in3 => \N__14827\,
            lcout => \eeprom.n3102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2033_3_lut_LC_18_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14581\,
            in2 => \N__13154\,
            in3 => \N__18101\,
            lcout => \eeprom.n3109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2035_3_lut_LC_18_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14843\,
            in2 => \N__18133\,
            in3 => \N__13166\,
            lcout => \eeprom.n3111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2041_3_lut_LC_18_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13109\,
            in2 => \N__14492\,
            in3 => \N__18100\,
            lcout => \eeprom.n3117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2031_3_lut_LC_18_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13127\,
            in2 => \N__18134\,
            in3 => \N__14644\,
            lcout => \eeprom.n3107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i8_4_lut_adj_79_LC_18_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14716\,
            in1 => \N__14817\,
            in2 => \N__14620\,
            in3 => \N__13246\,
            lcout => \eeprom.n21_adj_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_88_LC_18_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14842\,
            in1 => \N__14580\,
            in2 => \N__14543\,
            in3 => \N__14654\,
            lcout => \eeprom.n3034\,
            ltout => \eeprom.n3034_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2039_3_lut_LC_18_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13193\,
            in2 => \N__13115\,
            in3 => \N__14512\,
            lcout => \eeprom.n3115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_2_lut_LC_18_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24196\,
            in2 => \_gnd_net_\,
            in3 => \N__13112\,
            lcout => \eeprom.n3086\,
            ltout => OPEN,
            carryin => \bfn_18_29_0_\,
            carryout => \eeprom.n4105\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_3_lut_LC_18_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14491\,
            in2 => \N__28560\,
            in3 => \N__13103\,
            lcout => \eeprom.n3085\,
            ltout => OPEN,
            carryin => \eeprom.n4105\,
            carryout => \eeprom.n4106\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_4_lut_LC_18_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14342\,
            in3 => \N__13088\,
            lcout => \eeprom.n3084\,
            ltout => OPEN,
            carryin => \eeprom.n4106\,
            carryout => \eeprom.n4107\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_5_lut_LC_18_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14513\,
            in2 => \_gnd_net_\,
            in3 => \N__13187\,
            lcout => \eeprom.n3083\,
            ltout => OPEN,
            carryin => \eeprom.n4107\,
            carryout => \eeprom.n4108\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_6_lut_LC_18_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18281\,
            in3 => \N__13184\,
            lcout => \eeprom.n3082\,
            ltout => OPEN,
            carryin => \eeprom.n4108\,
            carryout => \eeprom.n4109\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_7_lut_LC_18_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14456\,
            in3 => \N__13172\,
            lcout => \eeprom.n3081\,
            ltout => OPEN,
            carryin => \eeprom.n4109\,
            carryout => \eeprom.n4110\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_8_lut_LC_18_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18260\,
            in3 => \N__13169\,
            lcout => \eeprom.n3080\,
            ltout => OPEN,
            carryin => \eeprom.n4110\,
            carryout => \eeprom.n4111\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_9_lut_LC_18_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14841\,
            in2 => \N__28561\,
            in3 => \N__13160\,
            lcout => \eeprom.n3079\,
            ltout => OPEN,
            carryin => \eeprom.n4111\,
            carryout => \eeprom.n4112\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_10_lut_LC_18_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28896\,
            in2 => \N__18017\,
            in3 => \N__13157\,
            lcout => \eeprom.n3078\,
            ltout => OPEN,
            carryin => \bfn_18_30_0_\,
            carryout => \eeprom.n4113\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_11_lut_LC_18_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28904\,
            in2 => \N__14582\,
            in3 => \N__13142\,
            lcout => \eeprom.n3077\,
            ltout => OPEN,
            carryin => \eeprom.n4113\,
            carryout => \eeprom.n4114\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_12_lut_LC_18_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14315\,
            in2 => \N__28934\,
            in3 => \N__13130\,
            lcout => \eeprom.n3076\,
            ltout => OPEN,
            carryin => \eeprom.n4114\,
            carryout => \eeprom.n4115\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_13_lut_LC_18_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28908\,
            in2 => \N__14648\,
            in3 => \N__13118\,
            lcout => \eeprom.n3075\,
            ltout => OPEN,
            carryin => \eeprom.n4115\,
            carryout => \eeprom.n4116\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_14_lut_LC_18_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28897\,
            in2 => \N__14723\,
            in3 => \N__13304\,
            lcout => \eeprom.n3074\,
            ltout => OPEN,
            carryin => \eeprom.n4116\,
            carryout => \eeprom.n4117\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_15_lut_LC_18_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14689\,
            in2 => \N__28932\,
            in3 => \N__13301\,
            lcout => \eeprom.n3073\,
            ltout => OPEN,
            carryin => \eeprom.n4117\,
            carryout => \eeprom.n4118\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_16_lut_LC_18_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14621\,
            in2 => \N__28935\,
            in3 => \N__13298\,
            lcout => \eeprom.n3072\,
            ltout => OPEN,
            carryin => \eeprom.n4118\,
            carryout => \eeprom.n4119\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_17_lut_LC_18_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13245\,
            in2 => \N__28933\,
            in3 => \N__13295\,
            lcout => \eeprom.n3071\,
            ltout => OPEN,
            carryin => \eeprom.n4119\,
            carryout => \eeprom.n4120\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_18_lut_LC_18_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14828\,
            in2 => \N__28936\,
            in3 => \N__13280\,
            lcout => \eeprom.n3070\,
            ltout => OPEN,
            carryin => \bfn_18_31_0_\,
            carryout => \eeprom.n4121\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_19_lut_LC_18_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14564\,
            in2 => \N__28937\,
            in3 => \N__13262\,
            lcout => \eeprom.n3069\,
            ltout => OPEN,
            carryin => \eeprom.n4121\,
            carryout => \eeprom.n4122\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2022_20_lut_LC_18_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28915\,
            in1 => \N__18673\,
            in2 => \N__18145\,
            in3 => \N__13259\,
            lcout => \eeprom.n3100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2027_3_lut_LC_18_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13256\,
            in2 => \N__13250\,
            in3 => \N__18138\,
            lcout => \eeprom.n3103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2444_3_lut_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13226\,
            in2 => \N__13202\,
            in3 => \N__13429\,
            lcout => \eeprom.n3712\,
            ltout => \eeprom.n3712_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4735_1_lut_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13391\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5565\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2449_3_lut_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13388\,
            in2 => \N__13382\,
            in3 => \N__13428\,
            lcout => \eeprom.n3717\,
            ltout => \eeprom.n3717_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4720_1_lut_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13367\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2450_rep_4_3_lut_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__13364\,
            in1 => \N__21578\,
            in2 => \_gnd_net_\,
            in3 => \N__13426\,
            lcout => \eeprom.n5362\,
            ltout => \eeprom.n5362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4717_1_lut_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13358\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5547\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2448_3_lut_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13567\,
            in2 => \N__13355\,
            in3 => \N__13427\,
            lcout => \eeprom.n3716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2447_3_lut_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13346\,
            in2 => \N__13339\,
            in3 => \N__13430\,
            lcout => \eeprom.n3715\,
            ltout => \eeprom.n3715_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4726_1_lut_LC_19_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13313\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5556\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_101_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__16329\,
            in1 => \N__15935\,
            in2 => \N__19088\,
            in3 => \N__13310\,
            lcout => OPEN,
            ltout => \eeprom.n5019_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_103_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__16424\,
            in1 => \N__16403\,
            in2 => \N__13484\,
            in3 => \N__16330\,
            lcout => OPEN,
            ltout => \eeprom.n28_adj_342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_104_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13544\,
            in1 => \N__16211\,
            in2 => \N__13481\,
            in3 => \N__13595\,
            lcout => \eeprom.n3628\,
            ltout => \eeprom.n3628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2446_3_lut_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110101"
        )
    port map (
            in0 => \N__13477\,
            in1 => \_gnd_net_\,
            in2 => \N__13463\,
            in3 => \N__13460\,
            lcout => \eeprom.n3714\,
            ltout => \eeprom.n3714_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4729_1_lut_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13454\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5559\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4741_2_lut_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__13450\,
            in1 => \_gnd_net_\,
            in2 => \N__13436\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n3711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_93_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__15977\,
            in1 => \N__16003\,
            in2 => \N__16321\,
            in3 => \N__13529\,
            lcout => OPEN,
            ltout => \eeprom.n5025_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_94_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__15961\,
            in1 => \N__15947\,
            in2 => \N__13400\,
            in3 => \N__16297\,
            lcout => OPEN,
            ltout => \eeprom.n5027_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_95_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__16298\,
            in1 => \N__15893\,
            in2 => \N__13397\,
            in3 => \N__15920\,
            lcout => OPEN,
            ltout => \eeprom.n5029_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_98_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111100"
        )
    port map (
            in0 => \N__16466\,
            in1 => \N__16486\,
            in2 => \N__13394\,
            in3 => \N__16299\,
            lcout => OPEN,
            ltout => \eeprom.n5031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_102_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13579\,
            in1 => \N__13616\,
            in2 => \N__13598\,
            in3 => \N__13625\,
            lcout => \eeprom.n5161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_24_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15960\,
            in1 => \N__15915\,
            in2 => \N__16487\,
            in3 => \N__19084\,
            lcout => \eeprom.n29_adj_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2376_3_lut_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__15757\,
            in1 => \N__15743\,
            in2 => \N__16322\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n3612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2381_3_lut_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15469\,
            in2 => \N__15449\,
            in3 => \N__16290\,
            lcout => \eeprom.n3617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2360_3_lut_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__16364\,
            in1 => \_gnd_net_\,
            in2 => \N__16319\,
            in3 => \N__16390\,
            lcout => \eeprom.n3596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2373_3_lut_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15655\,
            in2 => \N__15635\,
            in3 => \N__16277\,
            lcout => OPEN,
            ltout => \eeprom.n3609_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_91_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__16278\,
            in1 => \N__16130\,
            in2 => \N__13535\,
            in3 => \N__16100\,
            lcout => OPEN,
            ltout => \eeprom.n5021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_92_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__16091\,
            in1 => \N__16073\,
            in2 => \N__13532\,
            in3 => \N__16279\,
            lcout => \eeprom.n5023\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2302_3_lut_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13523\,
            in2 => \N__19220\,
            in3 => \N__13511\,
            lcout => \eeprom.n3506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2314_rep_5_3_lut_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13673\,
            in1 => \N__23426\,
            in2 => \_gnd_net_\,
            in3 => \N__19196\,
            lcout => \eeprom.n3518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2296_3_lut_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14075\,
            in1 => \_gnd_net_\,
            in2 => \N__19219\,
            in3 => \N__13661\,
            lcout => \eeprom.n3500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2372_3_lut_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__15593\,
            in1 => \_gnd_net_\,
            in2 => \N__15619\,
            in3 => \N__16283\,
            lcout => OPEN,
            ltout => \eeprom.n3608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_90_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111000"
        )
    port map (
            in0 => \N__16284\,
            in1 => \N__15671\,
            in2 => \N__13649\,
            in3 => \N__15691\,
            lcout => \eeprom.n5175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2308_3_lut_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13646\,
            in2 => \N__19204\,
            in3 => \N__16510\,
            lcout => \eeprom.n3512\,
            ltout => \eeprom.n3512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_96_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011000"
        )
    port map (
            in0 => \N__16285\,
            in1 => \N__15713\,
            in2 => \N__13637\,
            in3 => \N__13634\,
            lcout => OPEN,
            ltout => \eeprom.n5177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_97_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111010"
        )
    port map (
            in0 => \N__16031\,
            in1 => \N__16013\,
            in2 => \N__13628\,
            in3 => \N__16289\,
            lcout => \eeprom.n31_adj_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2362_3_lut_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16433\,
            in2 => \N__16320\,
            in3 => \N__16453\,
            lcout => \eeprom.n3598\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2311_3_lut_LC_19_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13607\,
            in2 => \N__19203\,
            in3 => \N__16618\,
            lcout => \eeprom.n3515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2313_3_lut_LC_19_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16657\,
            in2 => \N__13832\,
            in3 => \N__19161\,
            lcout => \eeprom.n3517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13820\,
            in3 => \N__13799\,
            lcout => OPEN,
            ltout => \eeprom.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_LC_19_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13779\,
            in1 => \N__13755\,
            in2 => \N__13736\,
            in3 => \N__17022\,
            lcout => OPEN,
            ltout => \eeprom.n30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i16_4_lut_LC_19_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13733\,
            in1 => \N__14012\,
            in2 => \N__13727\,
            in3 => \N__16682\,
            lcout => \eeprom.n3430\,
            ltout => \eeprom.n3430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2295_3_lut_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14056\,
            in2 => \N__13724\,
            in3 => \N__13721\,
            lcout => \eeprom.n3499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2294_3_lut_LC_19_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14035\,
            in2 => \N__19222\,
            in3 => \N__13709\,
            lcout => \eeprom.n3498\,
            ltout => \eeprom.n3498_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_18_LC_19_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16351\,
            in1 => \N__16380\,
            in2 => \N__13697\,
            in3 => \N__16449\,
            lcout => \eeprom.n28_adj_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2304_3_lut_LC_19_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__19214\,
            in1 => \_gnd_net_\,
            in2 => \N__17029\,
            in3 => \N__13682\,
            lcout => \eeprom.n3508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2233_3_lut_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14209\,
            in2 => \N__14105\,
            in3 => \N__17147\,
            lcout => \eeprom.n3405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2229_3_lut_LC_19_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__17148\,
            in1 => \_gnd_net_\,
            in2 => \N__14090\,
            in3 => \N__16790\,
            lcout => \eeprom.n3401\,
            ltout => \eeprom.n3401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_17_LC_19_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14052\,
            in1 => \N__14031\,
            in2 => \N__14015\,
            in3 => \N__14001\,
            lcout => \eeprom.n27_adj_263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2297_3_lut_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__14002\,
            in1 => \_gnd_net_\,
            in2 => \N__13988\,
            in3 => \N__19190\,
            lcout => \eeprom.n3501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_111_LC_19_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13968\,
            in1 => \N__13950\,
            in2 => \N__13924\,
            in3 => \N__13897\,
            lcout => OPEN,
            ltout => \eeprom.n28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i15_4_lut_LC_19_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14141\,
            in1 => \N__16757\,
            in2 => \N__13871\,
            in3 => \N__13868\,
            lcout => \eeprom.n3331\,
            ltout => \eeprom.n3331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2245_3_lut_LC_19_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13862\,
            in2 => \N__13850\,
            in3 => \N__16878\,
            lcout => \eeprom.n3417\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2173_3_lut_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17509\,
            in2 => \N__13847\,
            in3 => \N__17736\,
            lcout => \eeprom.n3313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_36_LC_19_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__24236\,
            in1 => \N__14358\,
            in2 => \N__17456\,
            in3 => \N__16990\,
            lcout => OPEN,
            ltout => \eeprom.n20_adj_301_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_adj_40_LC_19_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14422\,
            in1 => \N__14287\,
            in2 => \N__14273\,
            in3 => \N__18167\,
            lcout => OPEN,
            ltout => \eeprom.n28_adj_305_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i14_4_lut_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14270\,
            in1 => \N__14260\,
            in2 => \N__14240\,
            in3 => \N__14237\,
            lcout => \eeprom.n3232\,
            ltout => \eeprom.n3232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2166_3_lut_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14359\,
            in1 => \_gnd_net_\,
            in2 => \N__14231\,
            in3 => \N__14228\,
            lcout => \eeprom.n3306\,
            ltout => \eeprom.n3306_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_113_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14187\,
            in1 => \N__17170\,
            in2 => \N__14171\,
            in3 => \N__14157\,
            lcout => \eeprom.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4_4_lut_LC_19_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__22412\,
            in1 => \N__14874\,
            in2 => \N__17359\,
            in3 => \N__14135\,
            lcout => OPEN,
            ltout => \eeprom.n18_adj_260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i12_4_lut_adj_15_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15312\,
            in1 => \N__15270\,
            in2 => \N__14126\,
            in3 => \N__14123\,
            lcout => OPEN,
            ltout => \eeprom.n26_adj_262_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i13_4_lut_adj_16_LC_19_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14117\,
            in1 => \N__17983\,
            in2 => \N__14111\,
            in3 => \N__18033\,
            lcout => \eeprom.n3133\,
            ltout => \eeprom.n3133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2103_3_lut_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__18034\,
            in1 => \_gnd_net_\,
            in2 => \N__14108\,
            in3 => \N__15017\,
            lcout => \eeprom.n3211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2097_3_lut_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14855\,
            in2 => \N__17956\,
            in3 => \N__14875\,
            lcout => \eeprom.n3205\,
            ltout => \eeprom.n3205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2164_3_lut_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14408\,
            in2 => \N__14396\,
            in3 => \N__17762\,
            lcout => \eeprom.n3304\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2163_3_lut_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14392\,
            in2 => \N__17778\,
            in3 => \N__14378\,
            lcout => \eeprom.n3303\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2099_3_lut_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14930\,
            in2 => \N__14950\,
            in3 => \N__17941\,
            lcout => \eeprom.n3207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1973_3_lut_LC_19_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18380\,
            in2 => \N__19478\,
            in3 => \N__18740\,
            lcout => \eeprom.n3017\,
            ltout => \eeprom.n3017_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_77_LC_19_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14508\,
            in1 => \N__14442\,
            in2 => \N__14321\,
            in3 => \N__18236\,
            lcout => OPEN,
            ltout => \eeprom.n5147_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_78_LC_19_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__24189\,
            in1 => \N__14487\,
            in2 => \N__14318\,
            in3 => \N__14304\,
            lcout => \eeprom.n18_adj_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2108_3_lut_LC_19_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14744\,
            in2 => \N__14774\,
            in3 => \N__17922\,
            lcout => \eeprom.n3216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1965_3_lut_LC_19_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18476\,
            in2 => \N__18494\,
            in3 => \N__18741\,
            lcout => \eeprom.n3009\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1958_3_lut_LC_19_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18800\,
            in2 => \N__18774\,
            in3 => \N__19718\,
            lcout => \eeprom.n3002\,
            ltout => \eeprom.n3002_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_3_lut_LC_19_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18013\,
            in2 => \N__14546\,
            in3 => \N__18674\,
            lcout => \eeprom.n20_adj_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2034_3_lut_LC_19_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18009\,
            in2 => \N__14528\,
            in3 => \N__18128\,
            lcout => \eeprom.n3110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1972_3_lut_LC_19_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__18364\,
            in1 => \_gnd_net_\,
            in2 => \N__18350\,
            in3 => \N__18745\,
            lcout => \eeprom.n3016\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1974_3_lut_LC_19_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__18395\,
            in1 => \N__22466\,
            in2 => \N__18775\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n3018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1902_3_lut_LC_19_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20858\,
            in2 => \N__19379\,
            in3 => \N__19670\,
            lcout => \eeprom.n2914\,
            ltout => \eeprom.n2914_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_34_LC_19_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18327\,
            in1 => \N__18363\,
            in2 => \N__14468\,
            in3 => \N__18401\,
            lcout => \eeprom.n5301\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2029_3_lut_LC_19_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__14465\,
            in1 => \_gnd_net_\,
            in2 => \N__14690\,
            in3 => \N__18129\,
            lcout => \eeprom.n3105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1970_3_lut_LC_19_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18593\,
            in2 => \N__18617\,
            in3 => \N__18746\,
            lcout => \eeprom.n3014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1963_3_lut_LC_19_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18884\,
            in2 => \N__18776\,
            in3 => \N__18427\,
            lcout => \eeprom.n3007\,
            ltout => \eeprom.n3007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2030_3_lut_LC_19_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14705\,
            in2 => \N__14693\,
            in3 => \N__18109\,
            lcout => \eeprom.n3106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1962_3_lut_LC_19_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18872\,
            in2 => \N__18778\,
            in3 => \N__19589\,
            lcout => \eeprom.n3006\,
            ltout => \eeprom.n3006_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_85_LC_19_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14672\,
            in1 => \N__14643\,
            in2 => \N__14666\,
            in3 => \N__14663\,
            lcout => \eeprom.n24_adj_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1964_3_lut_LC_19_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18440\,
            in2 => \N__18777\,
            in3 => \N__18461\,
            lcout => \eeprom.n3008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1961_3_lut_LC_19_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18753\,
            in2 => \N__18860\,
            in3 => \N__18836\,
            lcout => \eeprom.n3005\,
            ltout => \eeprom.n3005_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2028_3_lut_LC_19_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18110\,
            in1 => \_gnd_net_\,
            in2 => \N__14603\,
            in3 => \N__14600\,
            lcout => \eeprom.n3104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2038_3_lut_LC_19_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18277\,
            in1 => \N__14588\,
            in2 => \_gnd_net_\,
            in3 => \N__18108\,
            lcout => \eeprom.n3114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1966_3_lut_LC_19_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18503\,
            in2 => \N__18784\,
            in3 => \N__19448\,
            lcout => \eeprom.n3010\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1968_3_lut_LC_19_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18545\,
            in2 => \N__18533\,
            in3 => \N__18770\,
            lcout => \eeprom.n3012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1959_3_lut_LC_19_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18809\,
            in2 => \N__18783\,
            in3 => \N__19775\,
            lcout => \eeprom.n3003\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2042_3_lut_LC_19_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__14801\,
            in1 => \N__24197\,
            in2 => \N__18143\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n3118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_2_lut_LC_19_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22411\,
            in2 => \_gnd_net_\,
            in3 => \N__14780\,
            lcout => \eeprom.n3186\,
            ltout => OPEN,
            carryin => \bfn_19_30_0_\,
            carryout => \eeprom.n4123\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_3_lut_LC_19_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28562\,
            in2 => \N__17352\,
            in3 => \N__14777\,
            lcout => \eeprom.n3185\,
            ltout => OPEN,
            carryin => \eeprom.n4123\,
            carryout => \eeprom.n4124\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_4_lut_LC_19_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14773\,
            in3 => \N__14735\,
            lcout => \eeprom.n3184\,
            ltout => OPEN,
            carryin => \eeprom.n4124\,
            carryout => \eeprom.n4125\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_5_lut_LC_19_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17446\,
            in3 => \N__14732\,
            lcout => \eeprom.n3183\,
            ltout => OPEN,
            carryin => \eeprom.n4125\,
            carryout => \eeprom.n4126\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_6_lut_LC_19_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17542\,
            in3 => \N__14729\,
            lcout => \eeprom.n3182\,
            ltout => OPEN,
            carryin => \eeprom.n4126\,
            carryout => \eeprom.n4127\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_7_lut_LC_19_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17629\,
            in3 => \N__14726\,
            lcout => \eeprom.n3181\,
            ltout => OPEN,
            carryin => \eeprom.n4127\,
            carryout => \eeprom.n4128\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_8_lut_LC_19_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15050\,
            in2 => \_gnd_net_\,
            in3 => \N__15020\,
            lcout => \eeprom.n3180\,
            ltout => OPEN,
            carryin => \eeprom.n4128\,
            carryout => \eeprom.n4129\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_9_lut_LC_19_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28563\,
            in2 => \N__18041\,
            in3 => \N__15005\,
            lcout => \eeprom.n3179\,
            ltout => OPEN,
            carryin => \eeprom.n4129\,
            carryout => \eeprom.n4130\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_10_lut_LC_19_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15002\,
            in2 => \N__28710\,
            in3 => \N__14963\,
            lcout => \eeprom.n3178\,
            ltout => OPEN,
            carryin => \bfn_19_31_0_\,
            carryout => \eeprom.n4131\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_11_lut_LC_19_31_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17984\,
            in2 => \N__28713\,
            in3 => \N__14960\,
            lcout => \eeprom.n3177\,
            ltout => OPEN,
            carryin => \eeprom.n4131\,
            carryout => \eeprom.n4132\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_12_lut_LC_19_31_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17299\,
            in2 => \N__28711\,
            in3 => \N__14957\,
            lcout => \eeprom.n3176\,
            ltout => OPEN,
            carryin => \eeprom.n4132\,
            carryout => \eeprom.n4133\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_13_lut_LC_19_31_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28576\,
            in2 => \N__14954\,
            in3 => \N__14918\,
            lcout => \eeprom.n3175\,
            ltout => OPEN,
            carryin => \eeprom.n4133\,
            carryout => \eeprom.n4134\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_14_lut_LC_19_31_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14914\,
            in2 => \N__28712\,
            in3 => \N__14879\,
            lcout => \eeprom.n3174\,
            ltout => OPEN,
            carryin => \eeprom.n4134\,
            carryout => \eeprom.n4135\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_15_lut_LC_19_31_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14876\,
            in2 => \N__28714\,
            in3 => \N__14846\,
            lcout => \eeprom.n3173\,
            ltout => OPEN,
            carryin => \eeprom.n4135\,
            carryout => \eeprom.n4136\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_16_lut_LC_19_31_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28586\,
            in2 => \N__15319\,
            in3 => \N__15278\,
            lcout => \eeprom.n3172\,
            ltout => OPEN,
            carryin => \eeprom.n4136\,
            carryout => \eeprom.n4137\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_17_lut_LC_19_31_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15271\,
            in2 => \N__28715\,
            in3 => \N__15233\,
            lcout => \eeprom.n3171\,
            ltout => OPEN,
            carryin => \eeprom.n4137\,
            carryout => \eeprom.n4138\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_18_lut_LC_19_32_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15225\,
            in2 => \N__28708\,
            in3 => \N__15194\,
            lcout => \eeprom.n3170\,
            ltout => OPEN,
            carryin => \bfn_19_32_0_\,
            carryout => \eeprom.n4139\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_19_lut_LC_19_32_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15191\,
            in2 => \N__28716\,
            in3 => \N__15155\,
            lcout => \eeprom.n3169\,
            ltout => OPEN,
            carryin => \eeprom.n4139\,
            carryout => \eeprom.n4140\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_20_lut_LC_19_32_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15152\,
            in2 => \N__28709\,
            in3 => \N__15107\,
            lcout => \eeprom.n3168\,
            ltout => OPEN,
            carryin => \eeprom.n4140\,
            carryout => \eeprom.n4141\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2089_21_lut_LC_19_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28593\,
            in1 => \N__15100\,
            in2 => \N__17957\,
            in3 => \N__15086\,
            lcout => \eeprom.n3199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_2_lut_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__25496\,
            in1 => \N__26708\,
            in2 => \N__25379\,
            in3 => \N__15056\,
            lcout => \eeprom.enable_N_60_0\,
            ltout => OPEN,
            carryin => \bfn_20_17_0_\,
            carryout => \eeprom.n4228\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_3_lut_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25667\,
            in1 => \N__23066\,
            in2 => \N__26737\,
            in3 => \N__15053\,
            lcout => \eeprom.enable_N_60_1\,
            ltout => OPEN,
            carryin => \eeprom.n4228\,
            carryout => \eeprom.n4229\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_4_lut_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__24812\,
            in1 => \N__26712\,
            in2 => \N__21974\,
            in3 => \N__15395\,
            lcout => \eeprom.enable_N_60_2\,
            ltout => OPEN,
            carryin => \eeprom.n4229\,
            carryout => \eeprom.n4230\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_5_lut_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25772\,
            in1 => \N__25319\,
            in2 => \N__26738\,
            in3 => \N__15392\,
            lcout => \eeprom.enable_N_60_3\,
            ltout => OPEN,
            carryin => \eeprom.n4230\,
            carryout => \eeprom.n4231\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_6_lut_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__24767\,
            in1 => \N__26716\,
            in2 => \N__21593\,
            in3 => \N__15389\,
            lcout => \eeprom.enable_N_60_4\,
            ltout => OPEN,
            carryin => \eeprom.n4231\,
            carryout => \eeprom.n4232\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_7_lut_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25361\,
            in1 => \N__19001\,
            in2 => \N__26739\,
            in3 => \N__15386\,
            lcout => \eeprom.enable_N_60_5\,
            ltout => OPEN,
            carryin => \eeprom.n4232\,
            carryout => \eeprom.n4233\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_8_lut_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__29408\,
            in1 => \N__26720\,
            in2 => \N__29369\,
            in3 => \N__15383\,
            lcout => \eeprom.enable_N_60_6\,
            ltout => OPEN,
            carryin => \eeprom.n4233\,
            carryout => \eeprom.n4234\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_9_lut_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__15380\,
            in1 => \N__26740\,
            in2 => \N__15374\,
            in3 => \N__15365\,
            lcout => \eeprom.enable_N_60_7\,
            ltout => OPEN,
            carryin => \eeprom.n4234\,
            carryout => \eeprom.n4235\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_10_lut_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__15362\,
            in1 => \N__26731\,
            in2 => \N__15356\,
            in3 => \N__15347\,
            lcout => \eeprom.enable_N_60_8\,
            ltout => OPEN,
            carryin => \bfn_20_18_0_\,
            carryout => \eeprom.n4236\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_11_lut_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__15491\,
            in1 => \N__15500\,
            in2 => \N__26744\,
            in3 => \N__15344\,
            lcout => \eeprom.enable_N_60_9\,
            ltout => OPEN,
            carryin => \eeprom.n4236\,
            carryout => \eeprom.n4237\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_12_lut_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__15341\,
            in1 => \N__26735\,
            in2 => \N__15335\,
            in3 => \N__15326\,
            lcout => \eeprom.enable_N_60_10\,
            ltout => OPEN,
            carryin => \eeprom.n4237\,
            carryout => \eeprom.n4238\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_13_lut_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__15584\,
            in1 => \N__26741\,
            in2 => \N__15578\,
            in3 => \N__15569\,
            lcout => \eeprom.enable_N_60_11\,
            ltout => OPEN,
            carryin => \eeprom.n4238\,
            carryout => \eeprom.n4239\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_14_lut_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__15566\,
            in1 => \N__26736\,
            in2 => \N__15557\,
            in3 => \N__15545\,
            lcout => \eeprom.enable_N_60_12\,
            ltout => OPEN,
            carryin => \eeprom.n4239\,
            carryout => \eeprom.n4240\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_15_lut_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__15542\,
            in1 => \N__26742\,
            in2 => \N__15536\,
            in3 => \N__15527\,
            lcout => \eeprom.enable_N_60_13\,
            ltout => OPEN,
            carryin => \eeprom.n4240\,
            carryout => \eeprom.n4241\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2473_16_lut_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__26743\,
            in1 => \N__15524\,
            in2 => \N__15518\,
            in3 => \N__15503\,
            lcout => \eeprom.enable_N_60_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4723_1_lut_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15499\,
            lcout => \eeprom.n5553\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_2_lut_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29458\,
            in2 => \_gnd_net_\,
            in3 => \N__15473\,
            lcout => \eeprom.n3586\,
            ltout => OPEN,
            carryin => \bfn_20_19_0_\,
            carryout => \eeprom.n4205\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_3_lut_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28504\,
            in2 => \N__15470\,
            in3 => \N__15440\,
            lcout => \eeprom.n3585_adj_296\,
            ltout => OPEN,
            carryin => \eeprom.n4205\,
            carryout => \eeprom.n4206\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_4_lut_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15437\,
            in3 => \N__15398\,
            lcout => \eeprom.n3584\,
            ltout => OPEN,
            carryin => \eeprom.n4206\,
            carryout => \eeprom.n4207\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_5_lut_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15884\,
            in3 => \N__15845\,
            lcout => \eeprom.n3583\,
            ltout => OPEN,
            carryin => \eeprom.n4207\,
            carryout => \eeprom.n4208\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_6_lut_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15842\,
            in3 => \N__15803\,
            lcout => \eeprom.n3582\,
            ltout => OPEN,
            carryin => \eeprom.n4208\,
            carryout => \eeprom.n4209\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_7_lut_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15800\,
            in3 => \N__15767\,
            lcout => \eeprom.n3581_adj_292\,
            ltout => OPEN,
            carryin => \eeprom.n4209\,
            carryout => \eeprom.n4210\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_8_lut_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15764\,
            in3 => \N__15734\,
            lcout => \eeprom.n3580\,
            ltout => OPEN,
            carryin => \eeprom.n4210\,
            carryout => \eeprom.n4211\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_9_lut_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28505\,
            in2 => \N__15731\,
            in3 => \N__15701\,
            lcout => \eeprom.n3579\,
            ltout => OPEN,
            carryin => \eeprom.n4211\,
            carryout => \eeprom.n4212\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_10_lut_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28633\,
            in2 => \N__15698\,
            in3 => \N__15665\,
            lcout => \eeprom.n3578\,
            ltout => OPEN,
            carryin => \bfn_20_20_0_\,
            carryout => \eeprom.n4213\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_11_lut_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28644\,
            in2 => \N__15662\,
            in3 => \N__15626\,
            lcout => \eeprom.n3577\,
            ltout => OPEN,
            carryin => \eeprom.n4213\,
            carryout => \eeprom.n4214\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_12_lut_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28634\,
            in2 => \N__15623\,
            in3 => \N__15587\,
            lcout => \eeprom.n3576\,
            ltout => OPEN,
            carryin => \eeprom.n4214\,
            carryout => \eeprom.n4215\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_13_lut_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16128\,
            in2 => \N__28759\,
            in3 => \N__16094\,
            lcout => \eeprom.n3575\,
            ltout => OPEN,
            carryin => \eeprom.n4215\,
            carryout => \eeprom.n4216\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_14_lut_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16090\,
            in2 => \N__28762\,
            in3 => \N__16067\,
            lcout => \eeprom.n3574\,
            ltout => OPEN,
            carryin => \eeprom.n4216\,
            carryout => \eeprom.n4217\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_15_lut_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16063\,
            in2 => \N__28760\,
            in3 => \N__16034\,
            lcout => \eeprom.n3573\,
            ltout => OPEN,
            carryin => \eeprom.n4217\,
            carryout => \eeprom.n4218\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_16_lut_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16030\,
            in2 => \N__28763\,
            in3 => \N__16007\,
            lcout => \eeprom.n3572\,
            ltout => OPEN,
            carryin => \eeprom.n4218\,
            carryout => \eeprom.n4219\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_17_lut_LC_20_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16004\,
            in2 => \N__28761\,
            in3 => \N__15971\,
            lcout => \eeprom.n3571\,
            ltout => OPEN,
            carryin => \eeprom.n4219\,
            carryout => \eeprom.n4220\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_18_lut_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15968\,
            in2 => \N__28554\,
            in3 => \N__15938\,
            lcout => \eeprom.n3570\,
            ltout => OPEN,
            carryin => \bfn_20_21_0_\,
            carryout => \eeprom.n4221\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_19_lut_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19074\,
            in2 => \N__28557\,
            in3 => \N__15923\,
            lcout => \eeprom.n3569\,
            ltout => OPEN,
            carryin => \eeprom.n4221\,
            carryout => \eeprom.n4222\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_20_lut_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15916\,
            in2 => \N__28555\,
            in3 => \N__16490\,
            lcout => \eeprom.n3568\,
            ltout => OPEN,
            carryin => \eeprom.n4222\,
            carryout => \eeprom.n4223\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_21_lut_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16485\,
            in2 => \N__28558\,
            in3 => \N__16457\,
            lcout => \eeprom.n3567\,
            ltout => OPEN,
            carryin => \eeprom.n4223\,
            carryout => \eeprom.n4224\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_22_lut_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28428\,
            in2 => \N__16454\,
            in3 => \N__16427\,
            lcout => \eeprom.n3566\,
            ltout => OPEN,
            carryin => \eeprom.n4224\,
            carryout => \eeprom.n4225\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_23_lut_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28418\,
            in2 => \N__16420\,
            in3 => \N__16394\,
            lcout => \eeprom.n3565\,
            ltout => OPEN,
            carryin => \eeprom.n4225\,
            carryout => \eeprom.n4226\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_24_lut_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16391\,
            in2 => \N__28556\,
            in3 => \N__16358\,
            lcout => \eeprom.n3564\,
            ltout => OPEN,
            carryin => \eeprom.n4226\,
            carryout => \eeprom.n4227\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_2357_25_lut_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28429\,
            in1 => \N__16355\,
            in2 => \N__16334\,
            in3 => \N__16214\,
            lcout => \eeprom.n5355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2242_3_lut_LC_20_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16199\,
            in2 => \N__17151\,
            in3 => \N__17659\,
            lcout => \eeprom.n3414\,
            ltout => \eeprom.n3414_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_LC_20_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16155\,
            in2 => \N__16136\,
            in3 => \N__16617\,
            lcout => OPEN,
            ltout => \eeprom.n5291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__16656\,
            in1 => \N__23422\,
            in2 => \N__16133\,
            in3 => \N__17201\,
            lcout => OPEN,
            ltout => \eeprom.n4824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16737\,
            in1 => \N__19254\,
            in2 => \N__16718\,
            in3 => \N__16714\,
            lcout => \eeprom.n28_adj_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2246_3_lut_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22670\,
            in1 => \N__16676\,
            in2 => \_gnd_net_\,
            in3 => \N__17115\,
            lcout => \eeprom.n3418\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2244_3_lut_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16637\,
            in2 => \N__17150\,
            in3 => \N__16952\,
            lcout => \eeprom.n3416\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2243_3_lut_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16906\,
            in2 => \N__16598\,
            in3 => \N__17119\,
            lcout => \eeprom.n3415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_108_LC_20_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17655\,
            in3 => \N__16572\,
            lcout => \eeprom.n5313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2231_3_lut_LC_20_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16819\,
            in2 => \N__16556\,
            in3 => \N__17125\,
            lcout => \eeprom.n3403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2174_3_lut_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17398\,
            in2 => \N__16541\,
            in3 => \N__17740\,
            lcout => \eeprom.n3314\,
            ltout => \eeprom.n3314_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2241_3_lut_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16526\,
            in2 => \N__16514\,
            in3 => \N__17123\,
            lcout => \eeprom.n3413\,
            ltout => \eeprom.n3413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_12_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17231\,
            in3 => \N__17217\,
            lcout => \eeprom.n5289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2170_3_lut_LC_20_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17195\,
            in2 => \N__17773\,
            in3 => \N__18223\,
            lcout => \eeprom.n3310\,
            ltout => \eeprom.n3310_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2237_3_lut_LC_20_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__17124\,
            in1 => \_gnd_net_\,
            in2 => \N__17048\,
            in3 => \N__17045\,
            lcout => \eeprom.n3409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2176_3_lut_LC_20_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__17006\,
            in1 => \N__17320\,
            in2 => \N__17771\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n3316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2177_3_lut_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16994\,
            in1 => \N__17735\,
            in2 => \_gnd_net_\,
            in3 => \N__16964\,
            lcout => \eeprom.n3317\,
            ltout => \eeprom.n3317_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_109_LC_20_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16924\,
            in2 => \N__16913\,
            in3 => \N__16905\,
            lcout => OPEN,
            ltout => \eeprom.n5315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_110_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__22666\,
            in1 => \N__16879\,
            in2 => \N__16856\,
            in3 => \N__16853\,
            lcout => OPEN,
            ltout => \eeprom.n4820_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_112_LC_20_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16836\,
            in1 => \N__16809\,
            in2 => \N__16793\,
            in3 => \N__16789\,
            lcout => \eeprom.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2175_3_lut_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17491\,
            in2 => \N__17801\,
            in3 => \N__17731\,
            lcout => \eeprom.n3315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2105_3_lut_LC_20_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17630\,
            in2 => \N__17600\,
            in3 => \N__17920\,
            lcout => \eeprom.n3213\,
            ltout => \eeprom.n3213_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_31_LC_20_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17561\,
            in3 => \N__17388\,
            lcout => \eeprom.n5205\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2106_3_lut_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17558\,
            in2 => \N__17546\,
            in3 => \N__17919\,
            lcout => \eeprom.n3214\,
            ltout => \eeprom.n3214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_32_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17484\,
            in1 => \N__17319\,
            in2 => \N__17465\,
            in3 => \N__17462\,
            lcout => \eeprom.n5209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2107_3_lut_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17447\,
            in2 => \N__17417\,
            in3 => \N__17915\,
            lcout => \eeprom.n3215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2109_3_lut_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__17372\,
            in1 => \_gnd_net_\,
            in2 => \N__17948\,
            in3 => \N__17360\,
            lcout => \eeprom.n3217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2100_3_lut_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17300\,
            in2 => \N__17267\,
            in3 => \N__17921\,
            lcout => \eeprom.n3208\,
            ltout => \eeprom.n3208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_37_LC_20_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18216\,
            in1 => \N__17820\,
            in2 => \N__18197\,
            in3 => \N__18193\,
            lcout => \eeprom.n26_adj_302\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1969_3_lut_LC_20_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18574\,
            in2 => \N__18560\,
            in3 => \N__18723\,
            lcout => \eeprom.n3013\,
            ltout => \eeprom.n3013_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2036_3_lut_LC_20_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__18161\,
            in1 => \_gnd_net_\,
            in2 => \N__18149\,
            in3 => \N__18144\,
            lcout => \eeprom.n3112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_2_lut_LC_20_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19434\,
            in2 => \_gnd_net_\,
            in3 => \N__19317\,
            lcout => \eeprom.n18_adj_330\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1967_3_lut_LC_20_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__19318\,
            in1 => \_gnd_net_\,
            in2 => \N__18760\,
            in3 => \N__18518\,
            lcout => \eeprom.n3011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_LC_20_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__22465\,
            in1 => \N__18849\,
            in2 => \N__19474\,
            in3 => \N__17990\,
            lcout => \eeprom.n15_adj_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2101_3_lut_LC_20_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17979\,
            in2 => \N__17955\,
            in3 => \N__17849\,
            lcout => \eeprom.n3209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1904_3_lut_LC_20_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20960\,
            in2 => \N__19400\,
            in3 => \N__19643\,
            lcout => \eeprom.n2916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1898_3_lut_LC_20_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19535\,
            in2 => \N__19672\,
            in3 => \N__21365\,
            lcout => \eeprom.n2910\,
            ltout => \eeprom.n2910_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_67_LC_20_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19588\,
            in1 => \N__19790\,
            in2 => \N__18302\,
            in3 => \N__18299\,
            lcout => OPEN,
            ltout => \eeprom.n22_adj_331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i11_4_lut_adj_68_LC_20_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18426\,
            in1 => \N__18459\,
            in2 => \N__18293\,
            in3 => \N__18290\,
            lcout => \eeprom.n2935\,
            ltout => \eeprom.n2935_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1971_3_lut_LC_20_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__18311\,
            in1 => \_gnd_net_\,
            in2 => \N__18284\,
            in3 => \N__18331\,
            lcout => \eeprom.n3015\,
            ltout => \eeprom.n3015_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_76_LC_20_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18250\,
            in2 => \N__18239\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1894_3_lut_LC_20_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21163\,
            in2 => \N__19499\,
            in3 => \N__19644\,
            lcout => \eeprom.n2906\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1896_3_lut_LC_20_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19514\,
            in2 => \N__19673\,
            in3 => \N__21275\,
            lcout => \eeprom.n2908\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_LC_20_28_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21273\,
            in1 => \N__21210\,
            in2 => \N__21109\,
            in3 => \N__21074\,
            lcout => OPEN,
            ltout => \eeprom.n18_adj_290_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_adj_29_LC_20_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21364\,
            in1 => \N__21024\,
            in2 => \N__18230\,
            in3 => \N__21401\,
            lcout => OPEN,
            ltout => \eeprom.n20_adj_291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i10_4_lut_adj_30_LC_20_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19298\,
            in1 => \N__21310\,
            in2 => \N__18227\,
            in3 => \N__21159\,
            lcout => \eeprom.n2836\,
            ltout => \eeprom.n2836_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1903_3_lut_LC_20_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__19388\,
            in1 => \_gnd_net_\,
            in2 => \N__18407\,
            in3 => \N__20900\,
            lcout => \eeprom.n2915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1897_3_lut_LC_20_28_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21311\,
            in2 => \N__19526\,
            in3 => \N__19642\,
            lcout => \eeprom.n2909\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1905_3_lut_LC_20_28_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__20990\,
            in1 => \N__19409\,
            in2 => \N__19671\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1901_3_lut_LC_20_28_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__19364\,
            in1 => \_gnd_net_\,
            in2 => \N__20819\,
            in3 => \N__19638\,
            lcout => \eeprom.n2913\,
            ltout => \eeprom.n2913_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_33_LC_20_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18404\,
            in3 => \N__18609\,
            lcout => \eeprom.n5297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_2_lut_LC_20_29_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22464\,
            in2 => \_gnd_net_\,
            in3 => \N__18383\,
            lcout => \eeprom.n2986\,
            ltout => OPEN,
            carryin => \bfn_20_29_0_\,
            carryout => \eeprom.n4088\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_3_lut_LC_20_29_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19473\,
            in2 => \N__28559\,
            in3 => \N__18371\,
            lcout => \eeprom.n2985\,
            ltout => OPEN,
            carryin => \eeprom.n4088\,
            carryout => \eeprom.n4089\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_4_lut_LC_20_29_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18368\,
            in3 => \N__18338\,
            lcout => \eeprom.n2984\,
            ltout => OPEN,
            carryin => \eeprom.n4089\,
            carryout => \eeprom.n4090\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_5_lut_LC_20_29_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18335\,
            in3 => \N__18620\,
            lcout => \eeprom.n2983\,
            ltout => OPEN,
            carryin => \eeprom.n4090\,
            carryout => \eeprom.n4091\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_6_lut_LC_20_29_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18616\,
            in3 => \N__18581\,
            lcout => \eeprom.n2982\,
            ltout => OPEN,
            carryin => \eeprom.n4091\,
            carryout => \eeprom.n4092\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_7_lut_LC_20_29_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18578\,
            in3 => \N__18548\,
            lcout => \eeprom.n2981\,
            ltout => OPEN,
            carryin => \eeprom.n4092\,
            carryout => \eeprom.n4093\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_8_lut_LC_20_29_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18544\,
            in2 => \_gnd_net_\,
            in3 => \N__18521\,
            lcout => \eeprom.n2980\,
            ltout => OPEN,
            carryin => \eeprom.n4093\,
            carryout => \eeprom.n4094\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_9_lut_LC_20_29_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28433\,
            in2 => \N__19325\,
            in3 => \N__18506\,
            lcout => \eeprom.n2979\,
            ltout => OPEN,
            carryin => \eeprom.n4094\,
            carryout => \eeprom.n4095\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_10_lut_LC_20_30_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19447\,
            in2 => \N__28919\,
            in3 => \N__18497\,
            lcout => \eeprom.n2978\,
            ltout => OPEN,
            carryin => \bfn_20_30_0_\,
            carryout => \eeprom.n4096\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_11_lut_LC_20_30_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18493\,
            in2 => \N__28923\,
            in3 => \N__18464\,
            lcout => \eeprom.n2977\,
            ltout => OPEN,
            carryin => \eeprom.n4096\,
            carryout => \eeprom.n4097\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_12_lut_LC_20_30_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18460\,
            in2 => \N__28920\,
            in3 => \N__18431\,
            lcout => \eeprom.n2976\,
            ltout => OPEN,
            carryin => \eeprom.n4097\,
            carryout => \eeprom.n4098\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_13_lut_LC_20_30_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18428\,
            in2 => \N__28924\,
            in3 => \N__18875\,
            lcout => \eeprom.n2975\,
            ltout => OPEN,
            carryin => \eeprom.n4098\,
            carryout => \eeprom.n4099\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_14_lut_LC_20_30_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19578\,
            in2 => \N__28921\,
            in3 => \N__18863\,
            lcout => \eeprom.n2974\,
            ltout => OPEN,
            carryin => \eeprom.n4099\,
            carryout => \eeprom.n4100\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_15_lut_LC_20_30_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18856\,
            in2 => \N__28925\,
            in3 => \N__18827\,
            lcout => \eeprom.n2973\,
            ltout => OPEN,
            carryin => \eeprom.n4100\,
            carryout => \eeprom.n4101\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_16_lut_LC_20_30_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19741\,
            in2 => \N__28922\,
            in3 => \N__18812\,
            lcout => \eeprom.n2972\,
            ltout => OPEN,
            carryin => \eeprom.n4101\,
            carryout => \eeprom.n4102\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_17_lut_LC_20_30_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19771\,
            in2 => \N__28926\,
            in3 => \N__18803\,
            lcout => \eeprom.n2971\,
            ltout => OPEN,
            carryin => \eeprom.n4102\,
            carryout => \eeprom.n4103\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_18_lut_LC_20_31_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19714\,
            in2 => \N__28927\,
            in3 => \N__18788\,
            lcout => \eeprom.n2970\,
            ltout => OPEN,
            carryin => \bfn_20_31_0_\,
            carryout => \eeprom.n4104\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1955_19_lut_LC_20_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28440\,
            in1 => \N__19802\,
            in2 => \N__18785\,
            in3 => \N__18677\,
            lcout => \eeprom.n3001\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_41_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__18653\,
            in1 => \N__18647\,
            in2 => \_gnd_net_\,
            in3 => \N__18641\,
            lcout => OPEN,
            ltout => \eeprom.n4847_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_45_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18635\,
            in1 => \N__18626\,
            in2 => \N__18983\,
            in3 => \N__18980\,
            lcout => OPEN,
            ltout => \eeprom.n4853_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_46_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18974\,
            in1 => \N__18968\,
            in2 => \N__18962\,
            in3 => \N__18959\,
            lcout => OPEN,
            ltout => \eeprom.n4859_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_47_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__18953\,
            in1 => \N__18947\,
            in2 => \N__18941\,
            in3 => \N__18938\,
            lcout => \eeprom.n4865\,
            ltout => \eeprom.n4865_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4699_4_lut_LC_21_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18925\,
            in1 => \N__18904\,
            in2 => \N__18932\,
            in3 => \N__18916\,
            lcout => OPEN,
            ltout => \eeprom.enable_N_59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rw_16_LC_21_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__27895\,
            in1 => \_gnd_net_\,
            in2 => \N__18929\,
            in3 => \_gnd_net_\,
            lcout => rw,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.enable_14_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18926\,
            in1 => \N__18917\,
            in2 => \N__18908\,
            in3 => \N__18893\,
            lcout => \eeprom.enable\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29860\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1423_3_lut_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22730\,
            in2 => \N__22700\,
            in3 => \N__23139\,
            lcout => \eeprom.n2211\,
            ltout => \eeprom.n2211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1490_3_lut_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19820\,
            in2 => \N__18887\,
            in3 => \N__21734\,
            lcout => \eeprom.n2310\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4676_3_lut_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22819\,
            in2 => \N__22844\,
            in3 => \N__23137\,
            lcout => \eeprom.n2215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1430_3_lut_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22373\,
            in1 => \N__24638\,
            in2 => \_gnd_net_\,
            in3 => \N__23138\,
            lcout => \eeprom.n2218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1493_3_lut_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19855\,
            in2 => \N__19841\,
            in3 => \N__21722\,
            lcout => \eeprom.n2313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1495_3_lut_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19889\,
            in2 => \N__19991\,
            in3 => \N__21723\,
            lcout => \eeprom.n2315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1426_3_lut_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22793\,
            in2 => \N__23315\,
            in3 => \N__23147\,
            lcout => \eeprom.n2214\,
            ltout => \eeprom.n2214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_52_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20226\,
            in1 => \N__19873\,
            in2 => \N__19004\,
            in3 => \N__19983\,
            lcout => \eeprom.n5045\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1497_3_lut_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19907\,
            in2 => \N__21738\,
            in3 => \N__19955\,
            lcout => \eeprom.n2317\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i6_3_lut_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__25802\,
            in1 => \N__29206\,
            in2 => \_gnd_net_\,
            in3 => \N__25360\,
            lcout => \eeprom.n3720\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_2_lut_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__24602\,
            in1 => \N__24601\,
            in2 => \N__20319\,
            in3 => \N__18992\,
            lcout => \eeprom.n2418\,
            ltout => OPEN,
            carryin => \bfn_21_20_0_\,
            carryout => \eeprom.n4007\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_3_lut_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20108\,
            in1 => \N__20107\,
            in2 => \N__20367\,
            in3 => \N__18989\,
            lcout => \eeprom.n2417\,
            ltout => OPEN,
            carryin => \eeprom.n4007\,
            carryout => \eeprom.n4008\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_4_lut_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20147\,
            in1 => \N__20146\,
            in2 => \N__20320\,
            in3 => \N__18986\,
            lcout => \eeprom.n2416\,
            ltout => OPEN,
            carryin => \eeprom.n4008\,
            carryout => \eeprom.n4009\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_5_lut_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20164\,
            in1 => \N__20165\,
            in2 => \N__20323\,
            in3 => \N__19031\,
            lcout => \eeprom.n2415\,
            ltout => OPEN,
            carryin => \eeprom.n4009\,
            carryout => \eeprom.n4010\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_6_lut_LC_21_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20062\,
            in1 => \N__20061\,
            in2 => \N__20321\,
            in3 => \N__19028\,
            lcout => \eeprom.n2414\,
            ltout => OPEN,
            carryin => \eeprom.n4010\,
            carryout => \eeprom.n4011\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_7_lut_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__20127\,
            in2 => \N__20324\,
            in3 => \N__19025\,
            lcout => \eeprom.n2413\,
            ltout => OPEN,
            carryin => \eeprom.n4011\,
            carryout => \eeprom.n4012\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_8_lut_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20042\,
            in1 => \N__20041\,
            in2 => \N__20322\,
            in3 => \N__19022\,
            lcout => \eeprom.n2412\,
            ltout => OPEN,
            carryin => \eeprom.n4012\,
            carryout => \eeprom.n4013\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_9_lut_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20405\,
            in1 => \N__20404\,
            in2 => \N__20368\,
            in3 => \N__19019\,
            lcout => \eeprom.n2411\,
            ltout => OPEN,
            carryin => \eeprom.n4013\,
            carryout => \eeprom.n4014\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_10_lut_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20273\,
            in1 => \N__20272\,
            in2 => \N__20369\,
            in3 => \N__19016\,
            lcout => \eeprom.n2410\,
            ltout => OPEN,
            carryin => \bfn_21_21_0_\,
            carryout => \eeprom.n4015\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_11_lut_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20087\,
            in1 => \N__20086\,
            in2 => \N__20371\,
            in3 => \N__19013\,
            lcout => \eeprom.n2409\,
            ltout => OPEN,
            carryin => \eeprom.n4015\,
            carryout => \eeprom.n4016\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_12_lut_LC_21_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20009\,
            in1 => \N__20008\,
            in2 => \N__20370\,
            in3 => \N__19010\,
            lcout => \eeprom.n2408\,
            ltout => OPEN,
            carryin => \eeprom.n4016\,
            carryout => \eeprom.n4017\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1553_13_lut_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20428\,
            in1 => \N__20429\,
            in2 => \N__20372\,
            in3 => \N__19007\,
            lcout => \eeprom.n2407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i2298_3_lut_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19258\,
            in2 => \N__19238\,
            in3 => \N__19207\,
            lcout => \eeprom.n3502\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1627_3_lut_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20582\,
            in2 => \N__20558\,
            in3 => \N__23486\,
            lcout => \eeprom.n2511\,
            ltout => \eeprom.n2511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1694_3_lut_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23969\,
            in2 => \N__19055\,
            in3 => \N__24434\,
            lcout => \eeprom.n2610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1702_3_lut_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23723\,
            in1 => \N__24320\,
            in2 => \_gnd_net_\,
            in3 => \N__24433\,
            lcout => \eeprom.n2618\,
            ltout => \eeprom.n2618_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1769_3_lut_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19046\,
            in2 => \N__19052\,
            in3 => \N__22563\,
            lcout => \eeprom.n2717\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_2_lut_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24286\,
            in2 => \_gnd_net_\,
            in3 => \N__19049\,
            lcout => \eeprom.n2686\,
            ltout => OPEN,
            carryin => \bfn_21_23_0_\,
            carryout => \eeprom.n4043\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_3_lut_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28134\,
            in2 => \N__22273\,
            in3 => \N__19040\,
            lcout => \eeprom.n2685\,
            ltout => OPEN,
            carryin => \eeprom.n4043\,
            carryout => \eeprom.n4044\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_4_lut_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23816\,
            in3 => \N__19037\,
            lcout => \eeprom.n2684\,
            ltout => OPEN,
            carryin => \eeprom.n4044\,
            carryout => \eeprom.n4045\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_5_lut_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23759\,
            in3 => \N__19034\,
            lcout => \eeprom.n2683\,
            ltout => OPEN,
            carryin => \eeprom.n4045\,
            carryout => \eeprom.n4046\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_6_lut_LC_21_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23876\,
            in3 => \N__19289\,
            lcout => \eeprom.n2682\,
            ltout => OPEN,
            carryin => \eeprom.n4046\,
            carryout => \eeprom.n4047\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_7_lut_LC_21_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23789\,
            in3 => \N__19286\,
            lcout => \eeprom.n2681\,
            ltout => OPEN,
            carryin => \eeprom.n4047\,
            carryout => \eeprom.n4048\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_8_lut_LC_21_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23846\,
            in3 => \N__19283\,
            lcout => \eeprom.n2680\,
            ltout => OPEN,
            carryin => \eeprom.n4048\,
            carryout => \eeprom.n4049\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_9_lut_LC_21_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22358\,
            in2 => \N__28287\,
            in3 => \N__19280\,
            lcout => \eeprom.n2679\,
            ltout => OPEN,
            carryin => \eeprom.n4049\,
            carryout => \eeprom.n4050\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_10_lut_LC_21_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22342\,
            in2 => \N__28288\,
            in3 => \N__19277\,
            lcout => \eeprom.n2678\,
            ltout => OPEN,
            carryin => \bfn_21_24_0_\,
            carryout => \eeprom.n4051\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_11_lut_LC_21_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28141\,
            in2 => \N__22309\,
            in3 => \N__19274\,
            lcout => \eeprom.n2677\,
            ltout => OPEN,
            carryin => \eeprom.n4051\,
            carryout => \eeprom.n4052\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_12_lut_LC_21_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22139\,
            in2 => \N__28289\,
            in3 => \N__19271\,
            lcout => \eeprom.n2676\,
            ltout => OPEN,
            carryin => \eeprom.n4052\,
            carryout => \eeprom.n4053\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_13_lut_LC_21_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22643\,
            in2 => \N__28290\,
            in3 => \N__19268\,
            lcout => \eeprom.n2675\,
            ltout => OPEN,
            carryin => \eeprom.n4053\,
            carryout => \eeprom.n4054\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_14_lut_LC_21_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28149\,
            in2 => \N__22622\,
            in3 => \N__19265\,
            lcout => \eeprom.n2674\,
            ltout => OPEN,
            carryin => \eeprom.n4054\,
            carryout => \eeprom.n4055\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_15_lut_LC_21_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22244\,
            in2 => \N__28291\,
            in3 => \N__19355\,
            lcout => \eeprom.n2673\,
            ltout => OPEN,
            carryin => \eeprom.n4055\,
            carryout => \eeprom.n4056\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1754_16_lut_LC_21_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28145\,
            in1 => \N__24335\,
            in2 => \N__22590\,
            in3 => \N__19352\,
            lcout => \eeprom.n2704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1761_3_lut_LC_21_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19349\,
            in2 => \N__22310\,
            in3 => \N__22580\,
            lcout => \eeprom.n2709\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1762_3_lut_LC_21_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19343\,
            in2 => \N__22592\,
            in3 => \N__22343\,
            lcout => \eeprom.n2710\,
            ltout => \eeprom.n2710_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_adj_84_LC_21_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21489\,
            in1 => \N__21177\,
            in2 => \N__19337\,
            in3 => \N__21223\,
            lcout => \eeprom.n17_adj_339\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1770_3_lut_LC_21_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__19334\,
            in1 => \_gnd_net_\,
            in2 => \N__22591\,
            in3 => \N__24282\,
            lcout => \eeprom.n2718\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1900_3_lut_LC_21_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19556\,
            in2 => \N__20786\,
            in3 => \N__19681\,
            lcout => \eeprom.n2912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_61_LC_21_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20889\,
            in1 => \N__20802\,
            in2 => \N__20958\,
            in3 => \N__19484\,
            lcout => OPEN,
            ltout => \eeprom.n5157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_LC_21_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__24256\,
            in1 => \N__20982\,
            in2 => \N__19301\,
            in3 => \N__20709\,
            lcout => \eeprom.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_60_LC_21_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20847\,
            in3 => \N__20778\,
            lcout => \eeprom.n5153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1906_3_lut_LC_21_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__24257\,
            in1 => \_gnd_net_\,
            in2 => \N__19421\,
            in3 => \N__19674\,
            lcout => \eeprom.n2918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1899_3_lut_LC_21_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__20710\,
            in1 => \_gnd_net_\,
            in2 => \N__19682\,
            in3 => \N__19544\,
            lcout => \eeprom.n2911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_2_lut_LC_21_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24255\,
            in2 => \_gnd_net_\,
            in3 => \N__19412\,
            lcout => \eeprom.n2886\,
            ltout => OPEN,
            carryin => \bfn_21_27_0_\,
            carryout => \eeprom.n4072\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_3_lut_LC_21_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20986\,
            in2 => \N__28841\,
            in3 => \N__19403\,
            lcout => \eeprom.n2885\,
            ltout => OPEN,
            carryin => \eeprom.n4072\,
            carryout => \eeprom.n4073\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_4_lut_LC_21_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20959\,
            in3 => \N__19391\,
            lcout => \eeprom.n2884\,
            ltout => OPEN,
            carryin => \eeprom.n4073\,
            carryout => \eeprom.n4074\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_5_lut_LC_21_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20896\,
            in2 => \_gnd_net_\,
            in3 => \N__19382\,
            lcout => \eeprom.n2883\,
            ltout => OPEN,
            carryin => \eeprom.n4074\,
            carryout => \eeprom.n4075\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_6_lut_LC_21_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20854\,
            in3 => \N__19367\,
            lcout => \eeprom.n2882\,
            ltout => OPEN,
            carryin => \eeprom.n4075\,
            carryout => \eeprom.n4076\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_7_lut_LC_21_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20815\,
            in3 => \N__19358\,
            lcout => \eeprom.n2881\,
            ltout => OPEN,
            carryin => \eeprom.n4076\,
            carryout => \eeprom.n4077\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_8_lut_LC_21_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20785\,
            in2 => \_gnd_net_\,
            in3 => \N__19547\,
            lcout => \eeprom.n2880\,
            ltout => OPEN,
            carryin => \eeprom.n4077\,
            carryout => \eeprom.n4078\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_9_lut_LC_21_27_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28721\,
            in2 => \N__20717\,
            in3 => \N__19538\,
            lcout => \eeprom.n2879\,
            ltout => OPEN,
            carryin => \eeprom.n4078\,
            carryout => \eeprom.n4079\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_10_lut_LC_21_28_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21360\,
            in2 => \N__28842\,
            in3 => \N__19529\,
            lcout => \eeprom.n2878\,
            ltout => OPEN,
            carryin => \bfn_21_28_0_\,
            carryout => \eeprom.n4080\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_11_lut_LC_21_28_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21304\,
            in2 => \N__28844\,
            in3 => \N__19517\,
            lcout => \eeprom.n2877\,
            ltout => OPEN,
            carryin => \eeprom.n4080\,
            carryout => \eeprom.n4081\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_12_lut_LC_21_28_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28733\,
            in2 => \N__21274\,
            in3 => \N__19505\,
            lcout => \eeprom.n2876\,
            ltout => OPEN,
            carryin => \eeprom.n4081\,
            carryout => \eeprom.n4082\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_13_lut_LC_21_28_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21211\,
            in2 => \N__28845\,
            in3 => \N__19502\,
            lcout => \eeprom.n2875\,
            ltout => OPEN,
            carryin => \eeprom.n4082\,
            carryout => \eeprom.n4083\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_14_lut_LC_21_28_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28737\,
            in2 => \N__21164\,
            in3 => \N__19490\,
            lcout => \eeprom.n2874\,
            ltout => OPEN,
            carryin => \eeprom.n4083\,
            carryout => \eeprom.n4084\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_15_lut_LC_21_28_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28725\,
            in2 => \N__21110\,
            in3 => \N__19487\,
            lcout => \eeprom.n2873\,
            ltout => OPEN,
            carryin => \eeprom.n4084\,
            carryout => \eeprom.n4085\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_16_lut_LC_21_28_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21072\,
            in2 => \N__28843\,
            in3 => \N__19811\,
            lcout => \eeprom.n2872\,
            ltout => OPEN,
            carryin => \eeprom.n4085\,
            carryout => \eeprom.n4086\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_17_lut_LC_21_28_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28729\,
            in2 => \N__21029\,
            in3 => \N__19808\,
            lcout => \eeprom.n2871\,
            ltout => OPEN,
            carryin => \eeprom.n4086\,
            carryout => \eeprom.n4087\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1888_18_lut_LC_21_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28153\,
            in1 => \N__21400\,
            in2 => \N__19680\,
            in3 => \N__19805\,
            lcout => \eeprom.n2902\,
            ltout => \eeprom.n2902_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_adj_62_LC_21_29_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__19770\,
            in1 => \N__19740\,
            in2 => \N__19793\,
            in3 => \N__19707\,
            lcout => \eeprom.n19_adj_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1892_3_lut_LC_21_29_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21073\,
            in1 => \_gnd_net_\,
            in2 => \N__19678\,
            in3 => \N__19781\,
            lcout => \eeprom.n2904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1893_3_lut_LC_21_29_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21102\,
            in1 => \_gnd_net_\,
            in2 => \N__19679\,
            in3 => \N__19754\,
            lcout => \eeprom.n2905\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1891_3_lut_LC_21_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__19724\,
            in1 => \_gnd_net_\,
            in2 => \N__21028\,
            in3 => \N__19656\,
            lcout => \eeprom.n2903\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1895_3_lut_LC_21_29_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21212\,
            in2 => \N__19691\,
            in3 => \N__19666\,
            lcout => \eeprom.n2907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_2_lut_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21998\,
            in3 => \N__19559\,
            lcout => \eeprom.n2286\,
            ltout => OPEN,
            carryin => \bfn_22_17_0_\,
            carryout => \eeprom.n3997\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_3_lut_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28190\,
            in2 => \N__19954\,
            in3 => \N__19895\,
            lcout => \eeprom.n2285\,
            ltout => OPEN,
            carryin => \eeprom.n3997\,
            carryout => \eeprom.n3998\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_4_lut_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20231\,
            in3 => \N__19892\,
            lcout => \eeprom.n2284\,
            ltout => OPEN,
            carryin => \eeprom.n3998\,
            carryout => \eeprom.n3999\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_5_lut_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19990\,
            in3 => \N__19880\,
            lcout => \eeprom.n2283\,
            ltout => OPEN,
            carryin => \eeprom.n3999\,
            carryout => \eeprom.n4000\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_6_lut_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19877\,
            in3 => \N__19862\,
            lcout => \eeprom.n2282\,
            ltout => OPEN,
            carryin => \eeprom.n4000\,
            carryout => \eeprom.n4001\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_7_lut_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19859\,
            in3 => \N__19829\,
            lcout => \eeprom.n2281\,
            ltout => OPEN,
            carryin => \eeprom.n4001\,
            carryout => \eeprom.n4002\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_8_lut_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20189\,
            in3 => \N__19826\,
            lcout => \eeprom.n2280\,
            ltout => OPEN,
            carryin => \eeprom.n4002\,
            carryout => \eeprom.n4003\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_9_lut_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21640\,
            in2 => \N__28352\,
            in3 => \N__19823\,
            lcout => \eeprom.n2279\,
            ltout => OPEN,
            carryin => \eeprom.n4003\,
            carryout => \eeprom.n4004\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_10_lut_LC_22_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28264\,
            in2 => \N__19925\,
            in3 => \N__19814\,
            lcout => \eeprom.n2278\,
            ltout => OPEN,
            carryin => \bfn_22_18_0_\,
            carryout => \eeprom.n4005\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_11_lut_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21955\,
            in2 => \N__28411\,
            in3 => \N__19997\,
            lcout => \eeprom.n2277\,
            ltout => OPEN,
            carryin => \eeprom.n4005\,
            carryout => \eeprom.n4006\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1486_12_lut_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__21737\,
            in1 => \N__28268\,
            in2 => \N__23090\,
            in3 => \N__19994\,
            lcout => \eeprom.n2308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1425_3_lut_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22777\,
            in2 => \N__23154\,
            in3 => \N__22757\,
            lcout => \eeprom.n2213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1428_3_lut_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22882\,
            in2 => \N__22862\,
            in3 => \N__23140\,
            lcout => \eeprom.n2216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_adj_51_LC_22_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23167\,
            in1 => \N__23026\,
            in2 => \N__22726\,
            in3 => \N__21647\,
            lcout => \eeprom.n2143\,
            ltout => \eeprom.n2143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1429_rep_44_3_lut_LC_22_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22912\,
            in2 => \N__19967\,
            in3 => \N__22898\,
            lcout => \eeprom.n2217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1498_3_lut_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21993\,
            in2 => \N__21739\,
            in3 => \N__19964\,
            lcout => \eeprom.n2318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_54_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__20184\,
            in1 => \N__19950\,
            in2 => \N__21997\,
            in3 => \N__19931\,
            lcout => OPEN,
            ltout => \eeprom.n4797_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4_4_lut_adj_55_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21636\,
            in1 => \N__19921\,
            in2 => \N__19910\,
            in3 => \N__21938\,
            lcout => \eeprom.n2242\,
            ltout => \eeprom.n2242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1427_rep_42_3_lut_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20171\,
            in2 => \N__20246\,
            in3 => \N__20243\,
            lcout => OPEN,
            ltout => \eeprom.n5400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4677_3_lut_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22977\,
            in2 => \N__20234\,
            in3 => \N__21680\,
            lcout => \eeprom.n2314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4679_3_lut_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20230\,
            in2 => \N__20210\,
            in3 => \N__21727\,
            lcout => \eeprom.n2316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1492_3_lut_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__20198\,
            in1 => \N__20185\,
            in2 => \N__21740\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1360_rep_47_3_lut_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22820\,
            in2 => \N__23155\,
            in3 => \N__21542\,
            lcout => \eeprom.n5405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_57_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20163\,
            in1 => \N__20145\,
            in2 => \N__20129\,
            in3 => \N__20024\,
            lcout => OPEN,
            ltout => \eeprom.n5085_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_58_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__24600\,
            in1 => \N__20106\,
            in2 => \N__20090\,
            in3 => \N__20085\,
            lcout => \eeprom.n7_adj_323\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_56_LC_22_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20063\,
            in3 => \N__20040\,
            lcout => \eeprom.n5081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1489_3_lut_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20018\,
            in2 => \N__21959\,
            in3 => \N__21736\,
            lcout => \eeprom.n2309\,
            ltout => \eeprom.n2309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2_2_lut_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20432\,
            in3 => \N__20271\,
            lcout => OPEN,
            ltout => \eeprom.n8_adj_322_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_59_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20421\,
            in1 => \N__20392\,
            in2 => \N__20381\,
            in3 => \N__20378\,
            lcout => \eeprom.n2341\,
            ltout => \eeprom.n2341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4746_1_lut_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20327\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1491_3_lut_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20282\,
            in2 => \N__21641\,
            in3 => \N__21735\,
            lcout => \eeprom.n2311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_26_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20454\,
            in2 => \N__21921\,
            in3 => \N__20607\,
            lcout => OPEN,
            ltout => \eeprom.n5073_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_27_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__21876\,
            in1 => \N__22441\,
            in2 => \N__20255\,
            in3 => \N__20483\,
            lcout => OPEN,
            ltout => \eeprom.n4782_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_28_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23526\,
            in1 => \N__20535\,
            in2 => \N__20252\,
            in3 => \N__21837\,
            lcout => OPEN,
            ltout => \eeprom.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_4_lut_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20577\,
            in1 => \N__21813\,
            in2 => \N__20249\,
            in3 => \N__20500\,
            lcout => \eeprom.n2440\,
            ltout => \eeprom.n2440_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1629_3_lut_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20455\,
            in2 => \N__20486\,
            in3 => \N__20441\,
            lcout => \eeprom.n2513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_25_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21765\,
            in3 => \N__22095\,
            lcout => \eeprom.n5071\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1628_3_lut_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20608\,
            in2 => \N__20594\,
            in3 => \N__23479\,
            lcout => \eeprom.n2512\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1624_3_lut_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__20536\,
            in1 => \N__20522\,
            in2 => \N__23493\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_2_lut_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22440\,
            in3 => \N__20477\,
            lcout => \eeprom.n2486\,
            ltout => OPEN,
            carryin => \bfn_22_22_0_\,
            carryout => \eeprom.n4018\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_3_lut_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21880\,
            in2 => \N__28549\,
            in3 => \N__20474\,
            lcout => \eeprom.n2485\,
            ltout => OPEN,
            carryin => \eeprom.n4018\,
            carryout => \eeprom.n4019\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_4_lut_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21772\,
            in3 => \N__20471\,
            lcout => \eeprom.n2484\,
            ltout => OPEN,
            carryin => \eeprom.n4019\,
            carryout => \eeprom.n4020\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_5_lut_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21925\,
            in3 => \N__20468\,
            lcout => \eeprom.n2483\,
            ltout => OPEN,
            carryin => \eeprom.n4020\,
            carryout => \eeprom.n4021\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_6_lut_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22108\,
            in3 => \N__20465\,
            lcout => \eeprom.n2482\,
            ltout => OPEN,
            carryin => \eeprom.n4021\,
            carryout => \eeprom.n4022\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_7_lut_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20462\,
            in3 => \N__20435\,
            lcout => \eeprom.n2481\,
            ltout => OPEN,
            carryin => \eeprom.n4022\,
            carryout => \eeprom.n4023\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_8_lut_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20612\,
            in2 => \_gnd_net_\,
            in3 => \N__20585\,
            lcout => \eeprom.n2480\,
            ltout => OPEN,
            carryin => \eeprom.n4023\,
            carryout => \eeprom.n4024\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_9_lut_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20581\,
            in2 => \N__28550\,
            in3 => \N__20549\,
            lcout => \eeprom.n2479\,
            ltout => OPEN,
            carryin => \eeprom.n4024\,
            carryout => \eeprom.n4025\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_10_lut_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28400\,
            in2 => \N__23539\,
            in3 => \N__20546\,
            lcout => \eeprom.n2478\,
            ltout => OPEN,
            carryin => \bfn_22_23_0_\,
            carryout => \eeprom.n4026\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_11_lut_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21844\,
            in2 => \N__28551\,
            in3 => \N__20543\,
            lcout => \eeprom.n2477\,
            ltout => OPEN,
            carryin => \eeprom.n4026\,
            carryout => \eeprom.n4027\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_12_lut_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20540\,
            in2 => \N__28553\,
            in3 => \N__20513\,
            lcout => \eeprom.n2476\,
            ltout => OPEN,
            carryin => \eeprom.n4027\,
            carryout => \eeprom.n4028\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_13_lut_LC_22_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21820\,
            in2 => \N__28552\,
            in3 => \N__20510\,
            lcout => \eeprom.n2475\,
            ltout => OPEN,
            carryin => \eeprom.n4028\,
            carryout => \eeprom.n4029\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1620_14_lut_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000101000"
        )
    port map (
            in0 => \N__23495\,
            in1 => \N__28407\,
            in2 => \N__20507\,
            in3 => \N__20489\,
            lcout => \eeprom.n2506\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i8_4_lut_adj_75_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22638\,
            in1 => \N__22615\,
            in2 => \N__22253\,
            in3 => \N__22280\,
            lcout => \eeprom.n2638\,
            ltout => \eeprom.n2638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1768_3_lut_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23809\,
            in2 => \N__20675\,
            in3 => \N__20672\,
            lcout => \eeprom.n2716\,
            ltout => \eeprom.n2716_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_81_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__22155\,
            in1 => \N__20916\,
            in2 => \N__20666\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1764_3_lut_LC_22_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23842\,
            in2 => \N__20663\,
            in3 => \N__22575\,
            lcout => \eeprom.n2712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1763_3_lut_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__20654\,
            in1 => \N__22357\,
            in2 => \N__22588\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1760_3_lut_LC_22_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22138\,
            in1 => \_gnd_net_\,
            in2 => \N__20648\,
            in3 => \N__22568\,
            lcout => \eeprom.n2708\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1759_3_lut_LC_22_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20639\,
            in2 => \N__22589\,
            in3 => \N__22642\,
            lcout => \eeprom.n2707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1757_3_lut_LC_22_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22243\,
            in2 => \N__20633\,
            in3 => \N__22576\,
            lcout => \eeprom.n2705\,
            ltout => \eeprom.n2705_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i6_4_lut_adj_83_LC_22_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21324\,
            in1 => \N__22500\,
            in2 => \N__20624\,
            in3 => \N__22175\,
            lcout => OPEN,
            ltout => \eeprom.n16_adj_338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i9_4_lut_adj_86_LC_22_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21126\,
            in1 => \N__20621\,
            in2 => \N__20615\,
            in3 => \N__20691\,
            lcout => \eeprom.n2737\,
            ltout => \eeprom.n2737_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4745_1_lut_LC_22_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20993\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_2_lut_LC_22_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22485\,
            in1 => \N__22487\,
            in2 => \N__20754\,
            in3 => \N__20963\,
            lcout => \eeprom.n2818\,
            ltout => OPEN,
            carryin => \bfn_22_25_0_\,
            carryout => \eeprom.n4057\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_3_lut_LC_22_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22209\,
            in1 => \N__22213\,
            in2 => \N__21443\,
            in3 => \N__20930\,
            lcout => \eeprom.n2817\,
            ltout => OPEN,
            carryin => \eeprom.n4057\,
            carryout => \eeprom.n4058\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_4_lut_LC_22_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20926\,
            in1 => \N__20927\,
            in2 => \N__20755\,
            in3 => \N__20876\,
            lcout => \eeprom.n2816\,
            ltout => OPEN,
            carryin => \eeprom.n4058\,
            carryout => \eeprom.n4059\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_5_lut_LC_22_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20873\,
            in1 => \N__20872\,
            in2 => \N__20758\,
            in3 => \N__20822\,
            lcout => \eeprom.n2815\,
            ltout => OPEN,
            carryin => \eeprom.n4059\,
            carryout => \eeprom.n4060\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_6_lut_LC_22_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22025\,
            in1 => \N__22024\,
            in2 => \N__20756\,
            in3 => \N__20789\,
            lcout => \eeprom.n2814\,
            ltout => OPEN,
            carryin => \eeprom.n4060\,
            carryout => \eeprom.n4061\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_7_lut_LC_22_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22157\,
            in1 => \N__22156\,
            in2 => \N__20759\,
            in3 => \N__20762\,
            lcout => \eeprom.n2813\,
            ltout => OPEN,
            carryin => \eeprom.n4061\,
            carryout => \eeprom.n4062\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_8_lut_LC_22_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22046\,
            in1 => \N__22042\,
            in2 => \N__20757\,
            in3 => \N__20696\,
            lcout => \eeprom.n2812\,
            ltout => OPEN,
            carryin => \eeprom.n4062\,
            carryout => \eeprom.n4063\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_9_lut_LC_22_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__20693\,
            in1 => \N__20692\,
            in2 => \N__21444\,
            in3 => \N__21335\,
            lcout => \eeprom.n2811\,
            ltout => OPEN,
            carryin => \eeprom.n4063\,
            carryout => \eeprom.n4064\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_10_lut_LC_22_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21332\,
            in1 => \N__21331\,
            in2 => \N__21469\,
            in3 => \N__21290\,
            lcout => \eeprom.n2810\,
            ltout => OPEN,
            carryin => \bfn_22_26_0_\,
            carryout => \eeprom.n4065\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_11_lut_LC_22_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21287\,
            in1 => \N__21286\,
            in2 => \N__21473\,
            in3 => \N__21239\,
            lcout => \eeprom.n2809\,
            ltout => OPEN,
            carryin => \eeprom.n4065\,
            carryout => \eeprom.n4066\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_12_lut_LC_22_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21236\,
            in1 => \N__21235\,
            in2 => \N__21470\,
            in3 => \N__21188\,
            lcout => \eeprom.n2808\,
            ltout => OPEN,
            carryin => \eeprom.n4066\,
            carryout => \eeprom.n4067\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_13_lut_LC_22_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21185\,
            in1 => \N__21184\,
            in2 => \N__21474\,
            in3 => \N__21137\,
            lcout => \eeprom.n2807\,
            ltout => OPEN,
            carryin => \eeprom.n4067\,
            carryout => \eeprom.n4068\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_14_lut_LC_22_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21134\,
            in1 => \N__21133\,
            in2 => \N__21471\,
            in3 => \N__21077\,
            lcout => \eeprom.n2806\,
            ltout => OPEN,
            carryin => \eeprom.n4068\,
            carryout => \eeprom.n4069\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_15_lut_LC_22_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__22510\,
            in1 => \N__22511\,
            in2 => \N__21475\,
            in3 => \N__21047\,
            lcout => \eeprom.n2805\,
            ltout => OPEN,
            carryin => \eeprom.n4069\,
            carryout => \eeprom.n4070\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_16_lut_LC_22_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21044\,
            in1 => \N__21043\,
            in2 => \N__21472\,
            in3 => \N__20996\,
            lcout => \eeprom.n2804\,
            ltout => OPEN,
            carryin => \eeprom.n4070\,
            carryout => \eeprom.n4071\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1821_17_lut_LC_22_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__21496\,
            in1 => \N__21497\,
            in2 => \N__21476\,
            in3 => \N__21404\,
            lcout => \eeprom.n2803\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_105_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23049\,
            in2 => \N__22978\,
            in3 => \N__23392\,
            lcout => OPEN,
            ltout => \eeprom.n5005_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_106_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__22941\,
            in1 => \N__21617\,
            in2 => \N__21380\,
            in3 => \N__22998\,
            lcout => OPEN,
            ltout => \eeprom.n5009_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_107_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__23231\,
            in1 => \N__23257\,
            in2 => \N__21377\,
            in3 => \N__23561\,
            lcout => \eeprom.n2044\,
            ltout => \eeprom.n2044_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1358_3_lut_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23050\,
            in1 => \_gnd_net_\,
            in2 => \N__21374\,
            in3 => \N__21524\,
            lcout => \eeprom.n2114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1360_3_lut_LC_23_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21541\,
            in2 => \N__22979\,
            in3 => \N__23341\,
            lcout => \eeprom.n2116\,
            ltout => \eeprom.n2116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_3_lut_adj_49_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22773\,
            in2 => \N__21371\,
            in3 => \N__22878\,
            lcout => \eeprom.n5061\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1361_3_lut_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21551\,
            in2 => \N__23003\,
            in3 => \N__23340\,
            lcout => \eeprom.n2117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1356_3_lut_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__21512\,
            in1 => \_gnd_net_\,
            in2 => \N__23358\,
            in3 => \N__23258\,
            lcout => \eeprom.n2112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_2_lut_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21616\,
            in2 => \_gnd_net_\,
            in3 => \N__21368\,
            lcout => \eeprom.n2086\,
            ltout => OPEN,
            carryin => \bfn_23_18_0_\,
            carryout => \eeprom.n3980\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_3_lut_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28242\,
            in2 => \N__23002\,
            in3 => \N__21545\,
            lcout => \eeprom.n2085\,
            ltout => OPEN,
            carryin => \eeprom.n3980\,
            carryout => \eeprom.n3981\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_4_lut_LC_23_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22976\,
            in3 => \N__21530\,
            lcout => \eeprom.n2084\,
            ltout => OPEN,
            carryin => \eeprom.n3981\,
            carryout => \eeprom.n3982\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_5_lut_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23393\,
            in3 => \N__21527\,
            lcout => \eeprom.n2083\,
            ltout => OPEN,
            carryin => \eeprom.n3982\,
            carryout => \eeprom.n3983\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_6_lut_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23054\,
            in3 => \N__21518\,
            lcout => \eeprom.n2082\,
            ltout => OPEN,
            carryin => \eeprom.n3983\,
            carryout => \eeprom.n3984\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_7_lut_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22942\,
            in3 => \N__21515\,
            lcout => \eeprom.n2081\,
            ltout => OPEN,
            carryin => \eeprom.n3984\,
            carryout => \eeprom.n3985\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_8_lut_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23256\,
            in3 => \N__21506\,
            lcout => \eeprom.n2080\,
            ltout => OPEN,
            carryin => \eeprom.n3985\,
            carryout => \eeprom.n3986\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_9_lut_LC_23_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23229\,
            in2 => \N__28393\,
            in3 => \N__21503\,
            lcout => \eeprom.n2079\,
            ltout => OPEN,
            carryin => \eeprom.n3986\,
            carryout => \eeprom.n3987\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1352_10_lut_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__28243\,
            in1 => \N__23363\,
            in2 => \N__23560\,
            in3 => \N__21500\,
            lcout => \eeprom.n2110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4671_3_lut_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__23364\,
            in1 => \N__23146\,
            in2 => \_gnd_net_\,
            in3 => \N__21721\,
            lcout => \eeprom.n5501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1422_3_lut_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__23144\,
            in1 => \N__23025\,
            in2 => \N__22682\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1357_3_lut_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21674\,
            in2 => \N__22943\,
            in3 => \N__23359\,
            lcout => \eeprom.n2113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1362_3_lut_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21615\,
            in1 => \_gnd_net_\,
            in2 => \N__23366\,
            in3 => \N__21668\,
            lcout => \eeprom.n2118\,
            ltout => \eeprom.n2118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_50_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__24634\,
            in1 => \N__21659\,
            in2 => \N__21650\,
            in3 => \N__23264\,
            lcout => \eeprom.n4788\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1424_3_lut_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22742\,
            in1 => \N__23284\,
            in2 => \_gnd_net_\,
            in3 => \N__23145\,
            lcout => \eeprom.n2212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i24_3_lut_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26429\,
            in1 => \N__29208\,
            in2 => \_gnd_net_\,
            in3 => \N__24983\,
            lcout => \eeprom.n2019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i5_3_lut_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__29212\,
            in1 => \_gnd_net_\,
            in2 => \N__25835\,
            in3 => \N__24763\,
            lcout => \eeprom.n3721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i8_3_lut_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26096\,
            in1 => \N__29210\,
            in2 => \_gnd_net_\,
            in3 => \N__25544\,
            lcout => \eeprom.n3619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i22_3_lut_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29209\,
            in1 => \N__26150\,
            in2 => \_gnd_net_\,
            in3 => \N__25025\,
            lcout => \eeprom.n2219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i3_3_lut_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__25883\,
            in1 => \N__29211\,
            in2 => \_gnd_net_\,
            in3 => \N__24808\,
            lcout => \eeprom.n3723\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_53_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23089\,
            in3 => \N__21954\,
            lcout => \eeprom.n6_adj_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1631_3_lut_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21932\,
            in2 => \N__23490\,
            in3 => \N__21926\,
            lcout => \eeprom.n2515\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1633_3_lut_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21893\,
            in2 => \N__21887\,
            in3 => \N__23467\,
            lcout => \eeprom.n2517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1625_3_lut_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21857\,
            in2 => \N__21848\,
            in3 => \N__23475\,
            lcout => \eeprom.n2509\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1623_3_lut_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21821\,
            in2 => \N__23492\,
            in3 => \N__21797\,
            lcout => \eeprom.n2507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1634_3_lut_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22442\,
            in1 => \N__21788\,
            in2 => \_gnd_net_\,
            in3 => \N__23466\,
            lcout => \eeprom.n2518\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1632_3_lut_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21779\,
            in2 => \N__23491\,
            in3 => \N__21773\,
            lcout => \eeprom.n2516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1630_3_lut_LC_23_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22118\,
            in2 => \N__22112\,
            in3 => \N__23474\,
            lcout => \eeprom.n2514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1695_3_lut_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__24019\,
            in1 => \_gnd_net_\,
            in2 => \N__24432\,
            in3 => \N__24002\,
            lcout => \eeprom.n2611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1701_3_lut_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23681\,
            in2 => \N__23707\,
            in3 => \N__24408\,
            lcout => \eeprom.n2617\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i5_4_lut_adj_66_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24493\,
            in1 => \N__23907\,
            in2 => \N__24355\,
            in3 => \N__24462\,
            lcout => OPEN,
            ltout => \eeprom.n13_adj_329_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_adj_69_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23989\,
            in1 => \N__24018\,
            in2 => \N__22079\,
            in3 => \N__23882\,
            lcout => \eeprom.n2539\,
            ltout => \eeprom.n2539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1697_3_lut_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24094\,
            in2 => \N__22076\,
            in3 => \N__24074\,
            lcout => \eeprom.n2613\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1767_3_lut_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23752\,
            in2 => \N__22073\,
            in3 => \N__22564\,
            lcout => \eeprom.n2715\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1765_3_lut_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23782\,
            in2 => \N__22587\,
            in3 => \N__22058\,
            lcout => \eeprom.n2713\,
            ltout => \eeprom.n2713_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_80_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22028\,
            in3 => \N__22011\,
            lcout => \eeprom.n5213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1696_3_lut_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__24061\,
            in1 => \N__24035\,
            in2 => \N__24436\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2612\,
            ltout => \eeprom.n2612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i7_4_lut_adj_74_LC_23_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22329\,
            in1 => \N__22220\,
            in2 => \N__22313\,
            in3 => \N__22308\,
            lcout => \eeprom.n16_adj_334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i21_1_lut_LC_23_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24920\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_adj_73_LC_23_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__24287\,
            in1 => \N__22134\,
            in2 => \N__23732\,
            in3 => \N__22274\,
            lcout => \eeprom.n12_adj_333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1690_3_lut_LC_23_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24470\,
            in2 => \N__24449\,
            in3 => \N__24422\,
            lcout => \eeprom.n2606\,
            ltout => \eeprom.n2606_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_72_LC_23_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22223\,
            in3 => \N__24331\,
            lcout => \eeprom.n10_adj_332\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_82_LC_23_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__22486\,
            in1 => \N__22214\,
            in2 => \N__22190\,
            in3 => \N__22181\,
            lcout => \eeprom.n4830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1766_3_lut_LC_23_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22169\,
            in2 => \N__23875\,
            in3 => \N__22561\,
            lcout => \eeprom.n2714\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1693_3_lut_LC_23_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23927\,
            in2 => \N__23954\,
            in3 => \N__24427\,
            lcout => \eeprom.n2609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i11_3_lut_LC_23_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26051\,
            in1 => \N__29204\,
            in2 => \_gnd_net_\,
            in3 => \N__25625\,
            lcout => \eeprom.n3319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1692_3_lut_LC_23_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__23917\,
            in1 => \_gnd_net_\,
            in2 => \N__24437\,
            in3 => \N__23894\,
            lcout => \eeprom.n2608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1691_3_lut_LC_23_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24508\,
            in2 => \N__24482\,
            in3 => \N__24431\,
            lcout => \eeprom.n2607\,
            ltout => \eeprom.n2607_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1758_3_lut_LC_23_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__22604\,
            in1 => \_gnd_net_\,
            in2 => \N__22595\,
            in3 => \N__22562\,
            lcout => \eeprom.n2706\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i17_3_lut_LC_23_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29176\,
            in1 => \N__26258\,
            in2 => \_gnd_net_\,
            in3 => \N__24956\,
            lcout => \eeprom.n2719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i15_3_lut_LC_23_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25967\,
            in1 => \N__29177\,
            in2 => \_gnd_net_\,
            in3 => \N__27581\,
            lcout => \eeprom.n2919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i20_3_lut_LC_23_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26201\,
            in1 => \N__29175\,
            in2 => \_gnd_net_\,
            in3 => \N__29348\,
            lcout => \eeprom.n2419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i13_3_lut_LC_23_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26012\,
            in1 => \N__29207\,
            in2 => \_gnd_net_\,
            in3 => \N__25691\,
            lcout => \eeprom.n3119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_2_lut_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24633\,
            in2 => \_gnd_net_\,
            in3 => \N__22361\,
            lcout => \eeprom.n2186\,
            ltout => OPEN,
            carryin => \bfn_24_17_0_\,
            carryout => \eeprom.n3988\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_3_lut_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28031\,
            in2 => \N__22916\,
            in3 => \N__22886\,
            lcout => \eeprom.n2185\,
            ltout => OPEN,
            carryin => \eeprom.n3988\,
            carryout => \eeprom.n3989\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_4_lut_LC_24_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22883\,
            in3 => \N__22847\,
            lcout => \eeprom.n2184\,
            ltout => OPEN,
            carryin => \eeprom.n3989\,
            carryout => \eeprom.n3990\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_5_lut_LC_24_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22837\,
            in3 => \N__22796\,
            lcout => \eeprom.n2183\,
            ltout => OPEN,
            carryin => \eeprom.n3990\,
            carryout => \eeprom.n3991\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_6_lut_LC_24_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23314\,
            in3 => \N__22781\,
            lcout => \eeprom.n2182\,
            ltout => OPEN,
            carryin => \eeprom.n3991\,
            carryout => \eeprom.n3992\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_7_lut_LC_24_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22778\,
            in3 => \N__22745\,
            lcout => \eeprom.n2181\,
            ltout => OPEN,
            carryin => \eeprom.n3992\,
            carryout => \eeprom.n3993\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_8_lut_LC_24_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23288\,
            in3 => \N__22733\,
            lcout => \eeprom.n2180\,
            ltout => OPEN,
            carryin => \eeprom.n3993\,
            carryout => \eeprom.n3994\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_9_lut_LC_24_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28032\,
            in2 => \N__22725\,
            in3 => \N__22685\,
            lcout => \eeprom.n2179\,
            ltout => OPEN,
            carryin => \eeprom.n3994\,
            carryout => \eeprom.n3995\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_10_lut_LC_24_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28318\,
            in2 => \N__23027\,
            in3 => \N__22673\,
            lcout => \eeprom.n2178\,
            ltout => OPEN,
            carryin => \bfn_24_18_0_\,
            carryout => \eeprom.n3996\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1419_11_lut_LC_24_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28319\,
            in1 => \N__23168\,
            in2 => \N__23156\,
            in3 => \N__23093\,
            lcout => \eeprom.n2209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i2_3_lut_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__25916\,
            in1 => \N__29213\,
            in2 => \_gnd_net_\,
            in3 => \N__25663\,
            lcout => \eeprom.n3724\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1291_3_lut_LC_24_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23180\,
            in2 => \N__25739\,
            in3 => \N__23596\,
            lcout => \eeprom.n2015\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1355_3_lut_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__23357\,
            in1 => \N__23230\,
            in2 => \N__23036\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1294_3_lut_LC_24_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__25145\,
            in1 => \_gnd_net_\,
            in2 => \N__23605\,
            in3 => \N__23210\,
            lcout => \eeprom.n2018\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3487_4_lut_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__25144\,
            in1 => \N__25459\,
            in2 => \N__25520\,
            in3 => \N__25703\,
            lcout => \eeprom.n1945\,
            ltout => \eeprom.n1945_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1293_3_lut_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23198\,
            in1 => \_gnd_net_\,
            in2 => \N__22982\,
            in3 => \N__25519\,
            lcout => \eeprom.n2017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1290_3_lut_LC_24_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__27808\,
            in1 => \_gnd_net_\,
            in2 => \N__23603\,
            in3 => \N__23636\,
            lcout => \eeprom.n2014\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1292_3_lut_LC_24_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23189\,
            in2 => \N__27701\,
            in3 => \N__23588\,
            lcout => \eeprom.n2016\,
            ltout => \eeprom.n2016_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1359_3_lut_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23375\,
            in2 => \N__23369\,
            in3 => \N__23365\,
            lcout => \eeprom.n2115\,
            ltout => \eeprom.n2115_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_48_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23291\,
            in3 => \N__23280\,
            lcout => \eeprom.n5059\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4674_3_lut_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__23627\,
            in1 => \_gnd_net_\,
            in2 => \N__23604\,
            in3 => \N__27613\,
            lcout => \eeprom.n2013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1288_3_lut_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25568\,
            in2 => \N__23618\,
            in3 => \N__23592\,
            lcout => \eeprom.n2012\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_2_lut_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25143\,
            in2 => \_gnd_net_\,
            in3 => \N__23201\,
            lcout => \eeprom.n1986\,
            ltout => OPEN,
            carryin => \bfn_24_20_0_\,
            carryout => \eeprom.n3973\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_3_lut_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25515\,
            in2 => \N__28594\,
            in3 => \N__23192\,
            lcout => \eeprom.n1985\,
            ltout => OPEN,
            carryin => \eeprom.n3973\,
            carryout => \eeprom.n3974\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_4_lut_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27700\,
            in3 => \N__23183\,
            lcout => \eeprom.n1984\,
            ltout => OPEN,
            carryin => \eeprom.n3974\,
            carryout => \eeprom.n3975\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_5_lut_LC_24_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25735\,
            in2 => \_gnd_net_\,
            in3 => \N__23171\,
            lcout => \eeprom.n1983\,
            ltout => OPEN,
            carryin => \eeprom.n3975\,
            carryout => \eeprom.n3976\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_6_lut_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27809\,
            in3 => \N__23630\,
            lcout => \eeprom.n1982\,
            ltout => OPEN,
            carryin => \eeprom.n3976\,
            carryout => \eeprom.n3977\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_7_lut_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27614\,
            in3 => \N__23621\,
            lcout => \eeprom.n1981\,
            ltout => OPEN,
            carryin => \eeprom.n3977\,
            carryout => \eeprom.n3978\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_8_lut_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25564\,
            in2 => \_gnd_net_\,
            in3 => \N__23609\,
            lcout => \eeprom.n1980\,
            ltout => OPEN,
            carryin => \eeprom.n3978\,
            carryout => \eeprom.n3979\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1285_9_lut_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__28477\,
            in1 => \N__25460\,
            in2 => \N__23606\,
            in3 => \N__23564\,
            lcout => \eeprom.n2011\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1626_3_lut_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23540\,
            in2 => \N__23510\,
            in3 => \N__23494\,
            lcout => \eeprom.n2510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i10_3_lut_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__29738\,
            in1 => \N__26078\,
            in2 => \_gnd_net_\,
            in3 => \N__29199\,
            lcout => \eeprom.n3419\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_63_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24130\,
            in3 => \N__24057\,
            lcout => OPEN,
            ltout => \eeprom.n5169_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_64_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24093\,
            in1 => \N__23664\,
            in2 => \N__23396\,
            in3 => \N__24162\,
            lcout => OPEN,
            ltout => \eeprom.n5173_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i3_4_lut_adj_65_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__24319\,
            in1 => \N__23940\,
            in2 => \N__23885\,
            in3 => \N__23700\,
            lcout => \eeprom.n11_adj_328\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1700_3_lut_LC_24_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__24418\,
            in1 => \N__23645\,
            in2 => \N__23671\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n2616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1698_3_lut_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24107\,
            in1 => \N__24129\,
            in2 => \_gnd_net_\,
            in3 => \N__24417\,
            lcout => \eeprom.n2614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1699_3_lut_LC_24_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24163\,
            in2 => \N__24435\,
            in3 => \N__24143\,
            lcout => \eeprom.n2615\,
            ltout => \eeprom.n2615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_70_LC_24_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23849\,
            in3 => \N__23832\,
            lcout => OPEN,
            ltout => \eeprom.n5101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_71_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23805\,
            in1 => \N__23778\,
            in2 => \N__23762\,
            in3 => \N__23748\,
            lcout => \eeprom.n5105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_2_lut_LC_24_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24312\,
            in3 => \N__23711\,
            lcout => \eeprom.n2586\,
            ltout => OPEN,
            carryin => \bfn_24_23_0_\,
            carryout => \eeprom.n4030\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_3_lut_LC_24_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28478\,
            in2 => \N__23708\,
            in3 => \N__23675\,
            lcout => \eeprom.n2585\,
            ltout => OPEN,
            carryin => \eeprom.n4030\,
            carryout => \eeprom.n4031\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_4_lut_LC_24_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23672\,
            in3 => \N__23639\,
            lcout => \eeprom.n2584\,
            ltout => OPEN,
            carryin => \eeprom.n4031\,
            carryout => \eeprom.n4032\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_5_lut_LC_24_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24167\,
            in3 => \N__24137\,
            lcout => \eeprom.n2583\,
            ltout => OPEN,
            carryin => \eeprom.n4032\,
            carryout => \eeprom.n4033\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_6_lut_LC_24_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24134\,
            in3 => \N__24101\,
            lcout => \eeprom.n2582\,
            ltout => OPEN,
            carryin => \eeprom.n4033\,
            carryout => \eeprom.n4034\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_7_lut_LC_24_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24098\,
            in3 => \N__24068\,
            lcout => \eeprom.n2581\,
            ltout => OPEN,
            carryin => \eeprom.n4034\,
            carryout => \eeprom.n4035\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_8_lut_LC_24_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24065\,
            in3 => \N__24029\,
            lcout => \eeprom.n2580\,
            ltout => OPEN,
            carryin => \eeprom.n4035\,
            carryout => \eeprom.n4036\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_9_lut_LC_24_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28479\,
            in2 => \N__24026\,
            in3 => \N__23996\,
            lcout => \eeprom.n2579\,
            ltout => OPEN,
            carryin => \eeprom.n4036\,
            carryout => \eeprom.n4037\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_10_lut_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28595\,
            in2 => \N__23993\,
            in3 => \N__23957\,
            lcout => \eeprom.n2578\,
            ltout => OPEN,
            carryin => \bfn_24_24_0_\,
            carryout => \eeprom.n4038\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_11_lut_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23947\,
            in2 => \N__28717\,
            in3 => \N__23921\,
            lcout => \eeprom.n2577\,
            ltout => OPEN,
            carryin => \eeprom.n4038\,
            carryout => \eeprom.n4039\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_12_lut_LC_24_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28599\,
            in2 => \N__23918\,
            in3 => \N__23888\,
            lcout => \eeprom.n2576\,
            ltout => OPEN,
            carryin => \eeprom.n4039\,
            carryout => \eeprom.n4040\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_13_lut_LC_24_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28500\,
            in2 => \N__24509\,
            in3 => \N__24473\,
            lcout => \eeprom.n2575\,
            ltout => OPEN,
            carryin => \eeprom.n4040\,
            carryout => \eeprom.n4041\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_14_lut_LC_24_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24469\,
            in2 => \N__28632\,
            in3 => \N__24440\,
            lcout => \eeprom.n2574\,
            ltout => OPEN,
            carryin => \eeprom.n4041\,
            carryout => \eeprom.n4042\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_add_1687_15_lut_LC_24_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001001000"
        )
    port map (
            in0 => \N__28600\,
            in1 => \N__24426\,
            in2 => \N__24362\,
            in3 => \N__24338\,
            lcout => \eeprom.n2605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i19_3_lut_LC_24_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26216\,
            in1 => \N__29198\,
            in2 => \_gnd_net_\,
            in3 => \N__25103\,
            lcout => \eeprom.n2519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i18_3_lut_LC_24_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26237\,
            in1 => \N__29178\,
            in2 => \_gnd_net_\,
            in3 => \N__25076\,
            lcout => \eeprom.n2619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i16_3_lut_LC_24_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29179\,
            in1 => \N__26282\,
            in2 => \_gnd_net_\,
            in3 => \N__29984\,
            lcout => \eeprom.n2819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i12_3_lut_LC_24_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26039\,
            in1 => \N__29180\,
            in2 => \_gnd_net_\,
            in3 => \N__29549\,
            lcout => \eeprom.n3219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i14_3_lut_LC_24_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25982\,
            in1 => \N__29203\,
            in2 => \_gnd_net_\,
            in3 => \N__24860\,
            lcout => \eeprom.n3019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_adj_9_LC_26_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__27423\,
            in1 => \N__27143\,
            in2 => \_gnd_net_\,
            in3 => \N__26886\,
            lcout => \eeprom.i2c.n534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3200_2_lut_LC_26_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26986\,
            in2 => \_gnd_net_\,
            in3 => \N__27028\,
            lcout => n3585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_adj_10_LC_26_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__25245\,
            in1 => \N__25168\,
            in2 => \_gnd_net_\,
            in3 => \N__26948\,
            lcout => n1805,
            ltout => \n1805_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i1_LC_26_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__24542\,
            in1 => \N__26560\,
            in2 => \N__24545\,
            in3 => \N__26521\,
            lcout => n170,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_adj_11_LC_26_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__25246\,
            in1 => \N__25169\,
            in2 => \_gnd_net_\,
            in3 => \N__26949\,
            lcout => n1800,
            ltout => \n1800_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i4_LC_26_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__24533\,
            in1 => \N__24527\,
            in2 => \N__24536\,
            in3 => \N__26522\,
            lcout => n164,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_36_i4_2_lut_LC_26_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__26987\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27032\,
            lcout => n4_adj_361,
            ltout => \n4_adj_361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i5_LC_26_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__24705\,
            in1 => \N__24518\,
            in2 => \N__24521\,
            in3 => \N__26523\,
            lcout => n162,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4589_3_lut_4_lut_4_lut_LC_26_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111111111"
        )
    port map (
            in0 => \N__27152\,
            in1 => \N__27516\,
            in2 => \N__26897\,
            in3 => \N__27419\,
            lcout => OPEN,
            ltout => \n5361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_26_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__26498\,
            in1 => \N__25183\,
            in2 => \N__24512\,
            in3 => \N__27884\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i0_LC_26_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__26499\,
            in1 => \N__24670\,
            in2 => \N__26564\,
            in3 => \N__24581\,
            lcout => n172,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29688\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_4_lut_LC_26_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100110011"
        )
    port map (
            in0 => \N__29785\,
            in1 => \N__27515\,
            in2 => \N__26519\,
            in3 => \N__27418\,
            lcout => OPEN,
            ltout => \n22_adj_367_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_26_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__26497\,
            in1 => \N__25182\,
            in2 => \N__24575\,
            in3 => \N__25166\,
            lcout => OPEN,
            ltout => \n4_adj_369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2_3_lut_4_lut_LC_26_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__27153\,
            in1 => \N__26891\,
            in2 => \N__24572\,
            in3 => \N__25247\,
            lcout => n4733,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_140_i11_2_lut_3_lut_4_lut_LC_26_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__27514\,
            in1 => \N__27151\,
            in2 => \N__27424\,
            in3 => \N__26887\,
            lcout => n11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_38_i4_2_lut_LC_26_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__27037\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26993\,
            lcout => n4,
            ltout => \n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i3_LC_26_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__24566\,
            in1 => \N__24712\,
            in2 => \N__24569\,
            in3 => \N__26514\,
            lcout => n166,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_143_i10_2_lut_LC_26_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27144\,
            in2 => \_gnd_net_\,
            in3 => \N__26893\,
            lcout => n10_adj_360,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i2_LC_26_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__24551\,
            in1 => \N__24676\,
            in2 => \N__24560\,
            in3 => \N__26513\,
            lcout => n168,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i7_LC_26_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__24692\,
            in1 => \N__24658\,
            in2 => \N__26524\,
            in3 => \N__24713\,
            lcout => n158,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4649_3_lut_4_lut_LC_26_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111011"
        )
    port map (
            in0 => \N__26894\,
            in1 => \N__27425\,
            in2 => \N__27160\,
            in3 => \N__27520\,
            lcout => OPEN,
            ltout => \n5461_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i1_LC_26_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111111"
        )
    port map (
            in0 => \N__27521\,
            in1 => \N__24686\,
            in2 => \N__24680\,
            in3 => \N__27176\,
            lcout => state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.data_out_i0_i6_LC_26_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__24644\,
            in1 => \N__24677\,
            in2 => \N__24659\,
            in3 => \N__26515\,
            lcout => n160,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29695\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i23_3_lut_LC_26_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26123\,
            in1 => \N__29173\,
            in2 => \_gnd_net_\,
            in3 => \N__25049\,
            lcout => \eeprom.n2119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i5_1_lut_LC_26_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24749\,
            lcout => \eeprom.n29_adj_278\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i14_1_lut_LC_26_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24856\,
            lcout => \eeprom.n20_adj_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i21_3_lut_LC_26_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__29174\,
            in1 => \N__26174\,
            in2 => \_gnd_net_\,
            in3 => \N__24919\,
            lcout => \eeprom.n2319\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i3_1_lut_LC_26_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24794\,
            lcout => \eeprom.n31_adj_286\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i0_LC_26_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25485\,
            in2 => \_gnd_net_\,
            in3 => \N__24818\,
            lcout => \eeprom.eeprom_counter_0\,
            ltout => OPEN,
            carryin => \bfn_26_21_0_\,
            carryout => \eeprom.n3931\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i1_LC_26_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25653\,
            in2 => \_gnd_net_\,
            in3 => \N__24815\,
            lcout => \eeprom.eeprom_counter_1\,
            ltout => OPEN,
            carryin => \eeprom.n3931\,
            carryout => \eeprom.n3932\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i2_LC_26_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24798\,
            in2 => \_gnd_net_\,
            in3 => \N__24773\,
            lcout => \eeprom.eeprom_counter_2\,
            ltout => OPEN,
            carryin => \eeprom.n3932\,
            carryout => \eeprom.n3933\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i3_LC_26_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25762\,
            in2 => \_gnd_net_\,
            in3 => \N__24770\,
            lcout => \eeprom.eeprom_counter_3\,
            ltout => OPEN,
            carryin => \eeprom.n3933\,
            carryout => \eeprom.n3934\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i4_LC_26_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24753\,
            in2 => \_gnd_net_\,
            in3 => \N__24728\,
            lcout => \eeprom.eeprom_counter_4\,
            ltout => OPEN,
            carryin => \eeprom.n3934\,
            carryout => \eeprom.n3935\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i5_LC_26_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25344\,
            in2 => \_gnd_net_\,
            in3 => \N__24725\,
            lcout => \eeprom.eeprom_counter_5\,
            ltout => OPEN,
            carryin => \eeprom.n3935\,
            carryout => \eeprom.n3936\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i6_LC_26_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29394\,
            in2 => \_gnd_net_\,
            in3 => \N__24722\,
            lcout => \eeprom.eeprom_counter_6\,
            ltout => OPEN,
            carryin => \eeprom.n3936\,
            carryout => \eeprom.n3937\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i7_LC_26_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25540\,
            in2 => \_gnd_net_\,
            in3 => \N__24719\,
            lcout => \eeprom.eeprom_counter_7\,
            ltout => OPEN,
            carryin => \eeprom.n3937\,
            carryout => \eeprom.n3938\,
            clk => \N__29861\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i8_LC_26_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29244\,
            in2 => \_gnd_net_\,
            in3 => \N__24716\,
            lcout => \eeprom.eeprom_counter_8\,
            ltout => OPEN,
            carryin => \bfn_26_22_0_\,
            carryout => \eeprom.n3939\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i9_LC_26_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29730\,
            in2 => \_gnd_net_\,
            in3 => \N__24872\,
            lcout => \eeprom.eeprom_counter_9\,
            ltout => OPEN,
            carryin => \eeprom.n3939\,
            carryout => \eeprom.n3940\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i10_LC_26_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25621\,
            in2 => \_gnd_net_\,
            in3 => \N__24869\,
            lcout => \eeprom.eeprom_counter_10\,
            ltout => OPEN,
            carryin => \eeprom.n3940\,
            carryout => \eeprom.n3941\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i11_LC_26_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29544\,
            in2 => \_gnd_net_\,
            in3 => \N__24866\,
            lcout => \eeprom.eeprom_counter_11\,
            ltout => OPEN,
            carryin => \eeprom.n3941\,
            carryout => \eeprom.n3942\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i12_LC_26_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25687\,
            in2 => \_gnd_net_\,
            in3 => \N__24863\,
            lcout => \eeprom.eeprom_counter_12\,
            ltout => OPEN,
            carryin => \eeprom.n3942\,
            carryout => \eeprom.n3943\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i13_LC_26_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24855\,
            in2 => \_gnd_net_\,
            in3 => \N__24833\,
            lcout => \eeprom.eeprom_counter_13\,
            ltout => OPEN,
            carryin => \eeprom.n3943\,
            carryout => \eeprom.n3944\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i14_LC_26_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27573\,
            in2 => \_gnd_net_\,
            in3 => \N__24830\,
            lcout => \eeprom.eeprom_counter_14\,
            ltout => OPEN,
            carryin => \eeprom.n3944\,
            carryout => \eeprom.n3945\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i15_LC_26_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29976\,
            in2 => \_gnd_net_\,
            in3 => \N__24827\,
            lcout => \eeprom.eeprom_counter_15\,
            ltout => OPEN,
            carryin => \eeprom.n3945\,
            carryout => \eeprom.n3946\,
            clk => \N__29863\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i16_LC_26_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24948\,
            in2 => \_gnd_net_\,
            in3 => \N__24824\,
            lcout => \eeprom.eeprom_counter_16\,
            ltout => OPEN,
            carryin => \bfn_26_23_0_\,
            carryout => \eeprom.n3947\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i17_LC_26_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25071\,
            in2 => \_gnd_net_\,
            in3 => \N__24821\,
            lcout => \eeprom.eeprom_counter_17\,
            ltout => OPEN,
            carryin => \eeprom.n3947\,
            carryout => \eeprom.n3948\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i18_LC_26_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25102\,
            in2 => \_gnd_net_\,
            in3 => \N__24926\,
            lcout => \eeprom.eeprom_counter_18\,
            ltout => OPEN,
            carryin => \eeprom.n3948\,
            carryout => \eeprom.n3949\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i19_LC_26_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29340\,
            in2 => \_gnd_net_\,
            in3 => \N__24923\,
            lcout => \eeprom.eeprom_counter_19\,
            ltout => OPEN,
            carryin => \eeprom.n3949\,
            carryout => \eeprom.n3950\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i20_LC_26_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24915\,
            in2 => \_gnd_net_\,
            in3 => \N__24893\,
            lcout => \eeprom.eeprom_counter_20\,
            ltout => OPEN,
            carryin => \eeprom.n3950\,
            carryout => \eeprom.n3951\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i21_LC_26_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25020\,
            in2 => \_gnd_net_\,
            in3 => \N__24890\,
            lcout => \eeprom.eeprom_counter_21\,
            ltout => OPEN,
            carryin => \eeprom.n3951\,
            carryout => \eeprom.n3952\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i22_LC_26_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25044\,
            in2 => \_gnd_net_\,
            in3 => \N__24887\,
            lcout => \eeprom.eeprom_counter_22\,
            ltout => OPEN,
            carryin => \eeprom.n3952\,
            carryout => \eeprom.n3953\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i23_LC_26_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24978\,
            in2 => \_gnd_net_\,
            in3 => \N__24884\,
            lcout => \eeprom.eeprom_counter_23\,
            ltout => OPEN,
            carryin => \eeprom.n3953\,
            carryout => \eeprom.n3954\,
            clk => \N__29865\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i24_LC_26_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25120\,
            in2 => \_gnd_net_\,
            in3 => \N__24881\,
            lcout => \eeprom.eeprom_counter_24\,
            ltout => OPEN,
            carryin => \bfn_26_24_0_\,
            carryout => \eeprom.n3955\,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i25_LC_26_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29496\,
            in2 => \_gnd_net_\,
            in3 => \N__24878\,
            lcout => \eeprom.eeprom_counter_25\,
            ltout => OPEN,
            carryin => \eeprom.n3955\,
            carryout => \eeprom.n3956\,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i26_LC_26_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29312\,
            in2 => \_gnd_net_\,
            in3 => \N__24875\,
            lcout => \eeprom.eeprom_counter_26\,
            ltout => OPEN,
            carryin => \eeprom.n3956\,
            carryout => \eeprom.n3957\,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i27_LC_26_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25438\,
            in2 => \_gnd_net_\,
            in3 => \N__24998\,
            lcout => \eeprom.eeprom_counter_27\,
            ltout => OPEN,
            carryin => \eeprom.n3957\,
            carryout => \eeprom.n3958\,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i28_LC_26_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25593\,
            in2 => \_gnd_net_\,
            in3 => \N__24995\,
            lcout => \eeprom.eeprom_counter_28\,
            ltout => OPEN,
            carryin => \eeprom.n3958\,
            carryout => \eeprom.n3959\,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i29_LC_26_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27778\,
            in2 => \_gnd_net_\,
            in3 => \N__24992\,
            lcout => \eeprom.eeprom_counter_29\,
            ltout => OPEN,
            carryin => \eeprom.n3959\,
            carryout => \eeprom.n3960\,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i30_LC_26_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25300\,
            in2 => \_gnd_net_\,
            in3 => \N__24989\,
            lcout => \eeprom.eeprom_counter_30\,
            ltout => OPEN,
            carryin => \eeprom.n3960\,
            carryout => \eeprom.n3961\,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.eeprom_counter_228__i31_LC_26_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29094\,
            in2 => \_gnd_net_\,
            in3 => \N__24986\,
            lcout => \eeprom.eeprom_counter_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29866\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i30_1_lut_LC_26_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27774\,
            lcout => \eeprom.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i27_1_lut_LC_26_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29304\,
            lcout => \eeprom.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i24_1_lut_LC_26_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24979\,
            lcout => \eeprom.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i17_1_lut_LC_26_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24955\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i28_1_lut_LC_26_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25434\,
            lcout => \eeprom.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i31_1_lut_LC_26_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25296\,
            lcout => \eeprom.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i25_3_lut_LC_26_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29090\,
            in2 => \N__26405\,
            in3 => \N__25119\,
            lcout => \eeprom.n1919\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i25_1_lut_LC_26_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25121\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i19_1_lut_LC_26_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25098\,
            lcout => \eeprom.n15_adj_295\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i18_1_lut_LC_26_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25072\,
            lcout => \eeprom.n16_adj_294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i23_1_lut_LC_26_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25045\,
            lcout => \eeprom.n11_adj_299\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i29_1_lut_LC_26_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25600\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i32_1_lut_LC_26_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29095\,
            lcout => \eeprom.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i22_1_lut_LC_26_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25021\,
            lcout => \eeprom.n12_adj_298\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter_i0_LC_27_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26947\,
            in2 => \_gnd_net_\,
            in3 => \N__25208\,
            lcout => \eeprom.i2c.counter_0\,
            ltout => OPEN,
            carryin => \bfn_27_17_0_\,
            carryout => \eeprom.i2c.n3899\,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.counter_i1_LC_27_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28003\,
            in2 => \N__27038\,
            in3 => \N__25205\,
            lcout => \eeprom.i2c.counter_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3899\,
            carryout => \eeprom.i2c.n3900\,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.counter_i2_LC_27_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26988\,
            in2 => \N__28103\,
            in3 => \N__25202\,
            lcout => \eeprom.i2c.counter_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3900\,
            carryout => \eeprom.i2c.n3901\,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.counter_i3_LC_27_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28007\,
            in2 => \N__26645\,
            in3 => \N__25199\,
            lcout => \eeprom.i2c.counter_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3901\,
            carryout => \eeprom.i2c.n3902\,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.counter_i4_LC_27_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26615\,
            in2 => \N__28104\,
            in3 => \N__25196\,
            lcout => \eeprom.i2c.counter_4\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3902\,
            carryout => \eeprom.i2c.n3903\,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.counter_i5_LC_27_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28011\,
            in2 => \N__26630\,
            in3 => \N__25193\,
            lcout => \eeprom.i2c.counter_5\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3903\,
            carryout => \eeprom.i2c.n3904\,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.counter_i6_LC_27_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26591\,
            in2 => \N__28105\,
            in3 => \N__25190\,
            lcout => \eeprom.i2c.counter_6\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3904\,
            carryout => \eeprom.i2c.n3905\,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.counter_i7_LC_27_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__26603\,
            in1 => \N__28015\,
            in2 => \_gnd_net_\,
            in3 => \N__25187\,
            lcout => \eeprom.i2c.counter_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29693\,
            ce => \N__25256\,
            sr => \N__25274\
        );

    \eeprom.i2c.i4657_3_lut_4_lut_LC_27_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001000"
        )
    port map (
            in0 => \N__25184\,
            in1 => \N__25167\,
            in2 => \N__26520\,
            in3 => \N__25244\,
            lcout => n5458,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i56_3_lut_LC_27_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__27367\,
            in1 => \N__27129\,
            in2 => \_gnd_net_\,
            in3 => \N__26815\,
            lcout => \eeprom.i2c.n33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i3_LC_27_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110101000"
        )
    port map (
            in0 => \N__27132\,
            in1 => \N__26753\,
            in2 => \N__25223\,
            in3 => \N__25280\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3794_2_lut_4_lut_LC_27_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__27369\,
            in1 => \N__27130\,
            in2 => \N__26895\,
            in3 => \N__26446\,
            lcout => \eeprom.i2c.n1913\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i20_4_lut_LC_27_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010001000100"
        )
    port map (
            in0 => \N__26447\,
            in1 => \N__25262\,
            in2 => \N__26576\,
            in3 => \N__25415\,
            lcout => \eeprom.i2c.n1829\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_144_i9_2_lut_LC_27_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__27368\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27513\,
            lcout => \eeprom.i2c.n9\,
            ltout => \eeprom.i2c.n9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_4_lut_LC_27_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101010"
        )
    port map (
            in0 => \N__26572\,
            in1 => \N__27065\,
            in2 => \N__25226\,
            in3 => \N__27055\,
            lcout => n1814,
            ltout => \n1814_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_LC_27_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__26752\,
            in1 => \_gnd_net_\,
            in2 => \N__25211\,
            in3 => \N__27131\,
            lcout => n471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_adj_8_LC_27_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__25400\,
            in1 => \N__25414\,
            in2 => \_gnd_net_\,
            in3 => \N__27526\,
            lcout => \eeprom.i2c.n1901\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i321_2_lut_LC_27_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27301\,
            in2 => \_gnd_net_\,
            in3 => \N__26912\,
            lcout => \state_7_N_162_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_4_lut_LC_27_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110010"
        )
    port map (
            in0 => \N__27385\,
            in1 => \N__27138\,
            in2 => \N__27522\,
            in3 => \N__26816\,
            lcout => \eeprom.i2c.n37\,
            ltout => \eeprom.i2c.n37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_adj_7_LC_27_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27493\,
            in2 => \N__25403\,
            in3 => \N__25399\,
            lcout => \eeprom.i2c.n39\,
            ltout => \eeprom.i2c.n39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4684_4_lut_LC_27_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__26819\,
            in1 => \N__27527\,
            in2 => \N__25391\,
            in3 => \N__25550\,
            lcout => \eeprom.i2c.n4513\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3_4_lut_4_lut_LC_27_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000010100"
        )
    port map (
            in0 => \N__26817\,
            in1 => \N__27386\,
            in2 => \N__27159\,
            in3 => \N__27494\,
            lcout => \eeprom.i2c.n407\,
            ltout => \eeprom.i2c.n407_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4692_4_lut_LC_27_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__27495\,
            in1 => \N__25388\,
            in2 => \N__25382\,
            in3 => \N__26818\,
            lcout => \eeprom.i2c.n524\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i1_3_lut_LC_27_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__25937\,
            in1 => \N__29171\,
            in2 => \_gnd_net_\,
            in3 => \N__25484\,
            lcout => \eeprom.n917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i6_1_lut_LC_27_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25340\,
            lcout => \eeprom.n28_adj_279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i4_3_lut_LC_27_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__25761\,
            in1 => \N__29172\,
            in2 => \_gnd_net_\,
            in3 => \N__25859\,
            lcout => \eeprom.n3722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i31_3_lut_LC_27_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29170\,
            in1 => \N__25304\,
            in2 => \_gnd_net_\,
            in3 => \N__26297\,
            lcout => \eeprom.n1256\,
            ltout => \eeprom.n1256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4559_2_lut_LC_27_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25571\,
            in3 => \N__27208\,
            lcout => \eeprom.n1913\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_3_lut_3_lut_LC_27_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__27406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27157\,
            lcout => \eeprom.i2c.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i8_1_lut_LC_27_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25536\,
            lcout => \eeprom.n26_adj_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2c_scl_enable_124_LC_27_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__27407\,
            in1 => \N__26892\,
            in2 => \N__27538\,
            in3 => \N__27158\,
            lcout => scl_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.i2c_scl_enable_124C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1226_3_lut_LC_27_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27268\,
            in2 => \N__27254\,
            in3 => \N__27636\,
            lcout => \eeprom.n1918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i1_1_lut_LC_27_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25489\,
            in3 => \_gnd_net_\,
            lcout => \eeprom.n33_adj_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1220_3_lut_4_lut_LC_27_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__29169\,
            in1 => \N__27854\,
            in2 => \N__28985\,
            in3 => \N__27637\,
            lcout => \eeprom.n1912\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i28_3_lut_LC_27_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29168\,
            in1 => \N__25442\,
            in2 => \_gnd_net_\,
            in3 => \N__26357\,
            lcout => \eeprom.n1139\,
            ltout => \eeprom.n1139_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1224_3_lut_LC_27_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__27230\,
            in1 => \_gnd_net_\,
            in2 => \N__25418\,
            in3 => \N__27635\,
            lcout => \eeprom.n1916\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i4_1_lut_LC_27_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25760\,
            lcout => \eeprom.n30_adj_277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_3_lut_LC_27_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27843\,
            in2 => \N__27209\,
            in3 => \N__27793\,
            lcout => OPEN,
            ltout => \eeprom.n5035_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_87_LC_27_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27681\,
            in1 => \N__25722\,
            in2 => \N__25706\,
            in3 => \N__27597\,
            lcout => \eeprom.n5039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i13_1_lut_LC_27_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25683\,
            lcout => \eeprom.n21_adj_264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i7_1_lut_LC_27_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29390\,
            lcout => \eeprom.n27_adj_280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i2_1_lut_LC_27_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25649\,
            lcout => \eeprom.n32_adj_288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i26_3_lut_LC_27_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__29096\,
            in1 => \_gnd_net_\,
            in2 => \N__29507\,
            in3 => \N__26393\,
            lcout => \eeprom.n892\,
            ltout => \eeprom.n892_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_42_LC_27_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__29291\,
            in1 => \N__29098\,
            in2 => \N__25628\,
            in3 => \N__26356\,
            lcout => \eeprom.n4977\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i11_1_lut_LC_27_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25617\,
            lcout => \eeprom.n23_adj_268\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i29_3_lut_LC_27_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29097\,
            in2 => \N__25601\,
            in3 => \N__26330\,
            lcout => \eeprom.n1138\,
            ltout => \eeprom.n1138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4557_1_lut_4_lut_LC_27_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__27654\,
            in1 => \N__28981\,
            in2 => \N__25952\,
            in3 => \N__27725\,
            lcout => \eeprom.n5327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_2_lut_LC_27_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25949\,
            in3 => \N__25928\,
            lcout => \eeprom.n33\,
            ltout => OPEN,
            carryin => \bfn_27_23_0_\,
            carryout => \eeprom.n4242\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_3_lut_LC_27_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25925\,
            in3 => \N__25901\,
            lcout => \eeprom.n32_adj_287\,
            ltout => OPEN,
            carryin => \eeprom.n4242\,
            carryout => \eeprom.n4243\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_4_lut_LC_27_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25898\,
            in3 => \N__25871\,
            lcout => \eeprom.n31_adj_285\,
            ltout => OPEN,
            carryin => \eeprom.n4243\,
            carryout => \eeprom.n4244\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_5_lut_LC_27_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25868\,
            in2 => \_gnd_net_\,
            in3 => \N__25850\,
            lcout => \eeprom.n30_adj_284\,
            ltout => OPEN,
            carryin => \eeprom.n4244\,
            carryout => \eeprom.n4245\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_6_lut_LC_27_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25847\,
            in3 => \N__25820\,
            lcout => \eeprom.n29_adj_283\,
            ltout => OPEN,
            carryin => \eeprom.n4245\,
            carryout => \eeprom.n4246\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_7_lut_LC_27_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25817\,
            in3 => \N__25787\,
            lcout => \eeprom.n28_adj_282\,
            ltout => OPEN,
            carryin => \eeprom.n4246\,
            carryout => \eeprom.n4247\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_8_lut_LC_27_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25784\,
            in3 => \N__25775\,
            lcout => \eeprom.n27_adj_281\,
            ltout => OPEN,
            carryin => \eeprom.n4247\,
            carryout => \eeprom.n4248\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_9_lut_LC_27_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26108\,
            in3 => \N__26084\,
            lcout => \eeprom.n26_adj_275\,
            ltout => OPEN,
            carryin => \eeprom.n4248\,
            carryout => \eeprom.n4249\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_10_lut_LC_27_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29222\,
            in3 => \N__26081\,
            lcout => \eeprom.n25_adj_271\,
            ltout => OPEN,
            carryin => \bfn_27_24_0_\,
            carryout => \eeprom.n4250\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_11_lut_LC_27_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29711\,
            in3 => \N__26066\,
            lcout => \eeprom.n24_adj_269\,
            ltout => OPEN,
            carryin => \eeprom.n4250\,
            carryout => \eeprom.n4251\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_12_lut_LC_27_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26063\,
            in3 => \N__26042\,
            lcout => \eeprom.n23\,
            ltout => OPEN,
            carryin => \eeprom.n4251\,
            carryout => \eeprom.n4252\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_13_lut_LC_27_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29522\,
            in3 => \N__26027\,
            lcout => \eeprom.n22_adj_265\,
            ltout => OPEN,
            carryin => \eeprom.n4252\,
            carryout => \eeprom.n4253\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_14_lut_LC_27_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26024\,
            in3 => \N__26000\,
            lcout => \eeprom.n21\,
            ltout => OPEN,
            carryin => \eeprom.n4253\,
            carryout => \eeprom.n4254\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_15_lut_LC_27_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25997\,
            in3 => \N__25970\,
            lcout => \eeprom.n20\,
            ltout => OPEN,
            carryin => \eeprom.n4254\,
            carryout => \eeprom.n4255\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_16_lut_LC_27_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27551\,
            in3 => \N__25955\,
            lcout => \eeprom.n19_adj_320\,
            ltout => OPEN,
            carryin => \eeprom.n4255\,
            carryout => \eeprom.n4256\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_17_lut_LC_27_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29957\,
            in3 => \N__26270\,
            lcout => \eeprom.n18_adj_326\,
            ltout => OPEN,
            carryin => \eeprom.n4256\,
            carryout => \eeprom.n4257\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_18_lut_LC_27_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26267\,
            in3 => \N__26249\,
            lcout => \eeprom.n17_adj_324\,
            ltout => OPEN,
            carryin => \bfn_27_25_0_\,
            carryout => \eeprom.n4258\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_19_lut_LC_27_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26246\,
            in3 => \N__26228\,
            lcout => \eeprom.n16_adj_325\,
            ltout => OPEN,
            carryin => \eeprom.n4258\,
            carryout => \eeprom.n4259\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_20_lut_LC_27_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26225\,
            in3 => \N__26204\,
            lcout => \eeprom.n15\,
            ltout => OPEN,
            carryin => \eeprom.n4259\,
            carryout => \eeprom.n4260\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_21_lut_LC_27_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29318\,
            in2 => \_gnd_net_\,
            in3 => \N__26192\,
            lcout => \eeprom.n14\,
            ltout => OPEN,
            carryin => \eeprom.n4260\,
            carryout => \eeprom.n4261\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_22_lut_LC_27_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26189\,
            in3 => \N__26162\,
            lcout => \eeprom.n13_adj_318\,
            ltout => OPEN,
            carryin => \eeprom.n4261\,
            carryout => \eeprom.n4262\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_23_lut_LC_27_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26159\,
            in3 => \N__26135\,
            lcout => \eeprom.n12_adj_319\,
            ltout => OPEN,
            carryin => \eeprom.n4262\,
            carryout => \eeprom.n4263\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_24_lut_LC_27_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26132\,
            in3 => \N__26111\,
            lcout => \eeprom.n11\,
            ltout => OPEN,
            carryin => \eeprom.n4263\,
            carryout => \eeprom.n4264\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_25_lut_LC_27_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26438\,
            in3 => \N__26417\,
            lcout => \eeprom.n10_adj_343\,
            ltout => OPEN,
            carryin => \eeprom.n4264\,
            carryout => \eeprom.n4265\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_26_lut_LC_27_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26414\,
            in3 => \N__26396\,
            lcout => \eeprom.n9_adj_308\,
            ltout => OPEN,
            carryin => \bfn_27_26_0_\,
            carryout => \eeprom.n4266\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_27_lut_LC_27_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29480\,
            in3 => \N__26381\,
            lcout => \eeprom.n8_adj_311\,
            ltout => OPEN,
            carryin => \eeprom.n4266\,
            carryout => \eeprom.n4267\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_28_lut_LC_27_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26378\,
            in3 => \N__26369\,
            lcout => \eeprom.n7_adj_309\,
            ltout => OPEN,
            carryin => \eeprom.n4267\,
            carryout => \eeprom.n4268\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_29_lut_LC_27_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26366\,
            in3 => \N__26342\,
            lcout => \eeprom.n6_adj_306\,
            ltout => OPEN,
            carryin => \eeprom.n4268\,
            carryout => \eeprom.n4269\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_30_lut_LC_27_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26339\,
            in3 => \N__26321\,
            lcout => \eeprom.n5_adj_317\,
            ltout => OPEN,
            carryin => \eeprom.n4269\,
            carryout => \eeprom.n4270\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_31_lut_LC_27_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26318\,
            in3 => \N__26309\,
            lcout => \eeprom.n4_adj_310\,
            ltout => OPEN,
            carryin => \eeprom.n4270\,
            carryout => \eeprom.n4271\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_32_lut_LC_27_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__26306\,
            in3 => \N__26285\,
            lcout => \eeprom.n3_adj_312\,
            ltout => OPEN,
            carryin => \eeprom.n4271\,
            carryout => \eeprom.n4272\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_add_3_33_lut_LC_27_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26659\,
            in2 => \_gnd_net_\,
            in3 => \N__26648\,
            lcout => \eeprom.n2_adj_307\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4695_2_lut_3_lut_4_lut_LC_28_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27405\,
            in1 => \N__26853\,
            in2 => \N__27161\,
            in3 => \N__27542\,
            lcout => n174,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i5_4_lut_LC_28_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26641\,
            in1 => \N__26626\,
            in2 => \N__26951\,
            in3 => \N__26614\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i6_4_lut_LC_28_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__26602\,
            in1 => \N__26590\,
            in2 => \N__26579\,
            in3 => \N__26550\,
            lcout => \eeprom.i2c.n464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.equal_41_i4_2_lut_LC_28_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26982\,
            lcout => n4_adj_358,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_142_i11_2_lut_3_lut_4_lut_LC_28_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__27541\,
            in1 => \N__27402\,
            in2 => \N__26877\,
            in3 => \N__27149\,
            lcout => n11_adj_359,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_7__I_0_137_i10_2_lut_LC_28_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27142\,
            in2 => \_gnd_net_\,
            in3 => \N__26839\,
            lcout => n10,
            ltout => \n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3809_3_lut_4_lut_LC_28_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__27539\,
            in1 => \N__27400\,
            in2 => \N__26534\,
            in3 => \N__26493\,
            lcout => \eeprom.i2c.n4579\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i2_LC_28_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110111"
        )
    port map (
            in0 => \N__27191\,
            in1 => \N__27185\,
            in2 => \N__26896\,
            in3 => \N__27175\,
            lcout => state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i2_2_lut_3_lut_4_lut_LC_28_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111101"
        )
    port map (
            in0 => \N__27540\,
            in1 => \N__27403\,
            in2 => \N__26878\,
            in3 => \N__27150\,
            lcout => OPEN,
            ltout => \n6_adj_365_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.state_i0_i0_LC_28_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111111"
        )
    port map (
            in0 => \N__27404\,
            in1 => \N__27044\,
            in2 => \N__27179\,
            in3 => \N__27174\,
            lcout => state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29687\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3258_2_lut_3_lut_LC_28_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__26840\,
            in1 => \N__27401\,
            in2 => \_gnd_net_\,
            in3 => \N__27148\,
            lcout => n3587,
            ltout => \n3587_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4641_4_lut_LC_28_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__29798\,
            in1 => \N__27443\,
            in2 => \N__27059\,
            in3 => \N__27056\,
            lcout => n5454,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4645_2_lut_LC_28_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27880\,
            in2 => \_gnd_net_\,
            in3 => \N__27036\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n5464_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4644_4_lut_LC_28_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000000000"
        )
    port map (
            in0 => \N__26989\,
            in1 => \N__26950\,
            in2 => \N__26918\,
            in3 => \N__27523\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n5451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.sda_out_133_LC_28_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000010111010"
        )
    port map (
            in0 => \N__27437\,
            in1 => \N__26854\,
            in2 => \N__26915\,
            in3 => \N__27408\,
            lcout => \eeprom.i2c.sda_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.sda_out_133C_net\,
            ce => \N__26906\,
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3210_2_lut_3_lut_LC_28_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111000"
        )
    port map (
            in0 => \N__27410\,
            in1 => \N__27525\,
            in2 => \N__26885\,
            in3 => \_gnd_net_\,
            lcout => n3595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3196_2_lut_LC_28_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__27524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27409\,
            lcout => n3581,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.write_enable_132_LC_28_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27436\,
            in2 => \_gnd_net_\,
            in3 => \N__27411\,
            lcout => sda_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeeprom.i2c.write_enable_132C_net\,
            ce => \N__27290\,
            sr => \N__27278\
        );

    \eeprom.add_822_2_lut_LC_28_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27269\,
            in3 => \N__27245\,
            lcout => \eeprom.n1198\,
            ltout => OPEN,
            carryin => \bfn_28_21_0_\,
            carryout => \eeprom.n4273\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_822_3_lut_LC_28_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28169\,
            in2 => \N__29273\,
            in3 => \N__27242\,
            lcout => \eeprom.n1197\,
            ltout => OPEN,
            carryin => \eeprom.n4273\,
            carryout => \eeprom.n4274\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_822_4_lut_LC_28_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27239\,
            in3 => \N__27224\,
            lcout => \eeprom.n1196\,
            ltout => OPEN,
            carryin => \eeprom.n4274\,
            carryout => \eeprom.n4275\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_822_5_lut_LC_28_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27746\,
            in3 => \N__27221\,
            lcout => \eeprom.n1195\,
            ltout => OPEN,
            carryin => \eeprom.n4275\,
            carryout => \eeprom.n4276\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_822_6_lut_LC_28_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27655\,
            in2 => \_gnd_net_\,
            in3 => \N__27218\,
            lcout => \eeprom.n1194\,
            ltout => OPEN,
            carryin => \eeprom.n4276\,
            carryout => \eeprom.n4277\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_822_7_lut_LC_28_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__27215\,
            in1 => \_gnd_net_\,
            in2 => \N__27844\,
            in3 => \N__27194\,
            lcout => \eeprom.n5328\,
            ltout => OPEN,
            carryin => \eeprom.n4277\,
            carryout => \eeprom.n4278\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.add_822_8_lut_LC_28_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28946\,
            in2 => \_gnd_net_\,
            in3 => \N__27857\,
            lcout => \eeprom.n1192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_2_lut_adj_44_LC_28_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27845\,
            in3 => \N__27713\,
            lcout => \eeprom.n1843\,
            ltout => \eeprom.n1843_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1223_3_lut_LC_28_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27742\,
            in2 => \N__27818\,
            in3 => \N__27815\,
            lcout => \eeprom.n1915\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i30_3_lut_LC_28_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__29185\,
            in1 => \N__27782\,
            in2 => \_gnd_net_\,
            in3 => \N__27758\,
            lcout => \eeprom.n1137\,
            ltout => \eeprom.n1137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i1_4_lut_adj_43_LC_28_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28980\,
            in1 => \N__27741\,
            in2 => \N__27728\,
            in3 => \N__27724\,
            lcout => \eeprom.n4983\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_i1225_3_lut_LC_28_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27707\,
            in2 => \N__27638\,
            in3 => \N__29272\,
            lcout => \eeprom.n1917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i4673_3_lut_LC_28_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27665\,
            in2 => \N__27659\,
            in3 => \N__27631\,
            lcout => \eeprom.n1914\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i15_1_lut_LC_28_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27580\,
            lcout => \eeprom.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i9_3_lut_LC_28_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29465\,
            in1 => \N__29205\,
            in2 => \_gnd_net_\,
            in3 => \N__29252\,
            lcout => \eeprom.n3519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i7_3_lut_LC_28_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__29414\,
            in1 => \N__29137\,
            in2 => \_gnd_net_\,
            in3 => \N__29404\,
            lcout => \eeprom.n3719\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i20_1_lut_LC_28_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29347\,
            lcout => \eeprom.n14_adj_297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_mux_3_i27_3_lut_LC_28_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29311\,
            in2 => \N__29184\,
            in3 => \N__29287\,
            lcout => \eeprom.n1140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i9_1_lut_LC_28_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29251\,
            lcout => \eeprom.n25_adj_272\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i401_2_lut_LC_28_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28967\,
            lcout => \eeprom.n1135\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_29_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.saved_addr__i1_LC_29_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__29797\,
            in1 => \N__27908\,
            in2 => \N__27902\,
            in3 => \N__27879\,
            lcout => saved_addr_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29658\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.enable_slow_121_LC_29_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__29632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29824\,
            lcout => \state_7_N_146_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29862\,
            ce => \N__29753\,
            sr => \N__29786\
        );

    \eeprom.i2c.i2c_clk_122_LC_29_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__29817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29625\,
            lcout => \eeprom.i2c.i2c_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29864\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_3_lut_LC_29_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__29624\,
            in1 => \N__29781\,
            in2 => \_gnd_net_\,
            in3 => \N__29816\,
            lcout => \eeprom.i2c.n1832\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i1_2_lut_LC_29_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29896\,
            in2 => \_gnd_net_\,
            in3 => \N__29941\,
            lcout => OPEN,
            ltout => \eeprom.i2c.n6_adj_255_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i4_4_lut_LC_29_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__29911\,
            in1 => \N__29878\,
            in2 => \N__29741\,
            in3 => \N__29926\,
            lcout => \eeprom.i2c.counter2_7__N_133\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i10_1_lut_LC_29_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29737\,
            lcout => \eeprom.n24_adj_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.i3188_2_lut_LC_29_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__29657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29578\,
            lcout => scl_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i12_1_lut_LC_29_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29545\,
            lcout => \eeprom.n22_adj_266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i26_1_lut_LC_29_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29503\,
            lcout => \eeprom.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.rem_4_unary_minus_2_inv_0_i16_1_lut_LC_29_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29983\,
            lcout => \eeprom.n18_adj_293\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eeprom.i2c.counter2_229_230__i1_LC_30_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29942\,
            in2 => \_gnd_net_\,
            in3 => \N__29930\,
            lcout => \eeprom.i2c.counter2_0\,
            ltout => OPEN,
            carryin => \bfn_30_20_0_\,
            carryout => \eeprom.i2c.n3962\,
            clk => \N__29867\,
            ce => 'H',
            sr => \N__29825\
        );

    \eeprom.i2c.counter2_229_230__i2_LC_30_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29927\,
            in2 => \_gnd_net_\,
            in3 => \N__29915\,
            lcout => \eeprom.i2c.counter2_1\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3962\,
            carryout => \eeprom.i2c.n3963\,
            clk => \N__29867\,
            ce => 'H',
            sr => \N__29825\
        );

    \eeprom.i2c.counter2_229_230__i3_LC_30_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29912\,
            in2 => \_gnd_net_\,
            in3 => \N__29900\,
            lcout => \eeprom.i2c.counter2_2\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3963\,
            carryout => \eeprom.i2c.n3964\,
            clk => \N__29867\,
            ce => 'H',
            sr => \N__29825\
        );

    \eeprom.i2c.counter2_229_230__i4_LC_30_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29897\,
            in2 => \_gnd_net_\,
            in3 => \N__29885\,
            lcout => \eeprom.i2c.counter2_3\,
            ltout => OPEN,
            carryin => \eeprom.i2c.n3964\,
            carryout => \eeprom.i2c.n3965\,
            clk => \N__29867\,
            ce => 'H',
            sr => \N__29825\
        );

    \eeprom.i2c.counter2_229_230__i5_LC_30_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29879\,
            in2 => \_gnd_net_\,
            in3 => \N__29882\,
            lcout => \eeprom.i2c.counter2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__29867\,
            ce => 'H',
            sr => \N__29825\
        );
end \INTERFACE\;
