// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Wed Oct  2 00:23:42 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    input PIN_3 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    input PIN_4 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    input PIN_5 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    output PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    output PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    output PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    output PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    output PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    input PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    inout PIN_20 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    inout PIN_21 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    inout PIN_22 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    input PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    input PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire GND_net, VCC_net, CLK_c, LED_c, PIN_6_c_0, PIN_7_c_1, PIN_8_c_2, 
        PIN_9_c_3, PIN_10_c_4, PIN_11_c_5, PIN_13_c, PIN_18_c_1, PIN_19_c_0, 
        PIN_23_c_1, PIN_24_c_0, tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(66[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(67[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(68[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(69[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(70[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(71[22:24])
    wire [23:0]Kd;   // verilog/TinyFPGA_B.v(72[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(73[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(74[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(75[22:35])
    wire [23:0]deadband;   // verilog/TinyFPGA_B.v(76[22:30])
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(77[22:34])
    
    wire hall1, hall2, hall3;
    wire [23:0]pwm;   // verilog/TinyFPGA_B.v(85[10:13])
    wire [31:0]motor_state;   // verilog/TinyFPGA_B.v(134[22:33])
    
    wire n47968;
    wire [31:0]motor_state_23__N_25;
    wire [24:0]displacement_23__N_91;
    wire [23:0]displacement_23__N_1;
    
    wire rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(88[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(92[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(92[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(92[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(92[12:19])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(93[12:25])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(94[12:26])
    
    wire n47840, n20136;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(94[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(99[12:33])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(109[11:16])
    
    wire n249, n248, n47838, n6, n38028, n38027, n38026, n38025, 
        n122, n38024, n48719, n38023, n4, n38022, n38021, n2, 
        n38020, n38019, n38018, n37168, n48713, n49157, n49266, 
        n38017, n38016, n38015, n47795, n37167, n2298, n2297, 
        n37166, n37165, n37164, n38014, n37163, n37162, n38013, 
        n37161, n38012, n37160, n37159, n37158, n38011, n37157, 
        n37156, n38010, n37155, n37154, n38009, n37153, n47783, 
        n47781, n38008, n38007, n37152, n37151, n47775, n38006, 
        n38005, n38004, n47773, n38003, n47755, n37150, n37149, 
        n24351, n24350, n24349, n6932, n48920, n47747, n22552, 
        n22549, n47743, n22546, n38002, n37148, n43238, n47722, 
        n47718, n22543, n22540, n37147, n22537, n38001, n22534, 
        n22531, n38000, n49264, n37999, n22528, n37998, n47690, 
        n29726, n22525, n37997, n22522, n2242, n47, n2296, n2295, 
        n2294, n2293, n2292, n2265, n2264, n2241, n37996, n37995, 
        n22519, n22516, n48753, n37146, n22513, n22510, n24332, 
        n22507, n37994, n44019, n37993, n47639, n44009, n47631, 
        Kp_23__N_515, n37992, n47628, n37991, n47623, n48548, n28794, 
        n37990, n28760, Kp_23__N_865, n47615, n103, n49262, n37989, 
        n4_adj_3960, n37988, n24253, n37987, n37986, n37985, n37984, 
        n37983, n24252, n24251, n24250, n47589, n24249, n24248, 
        n48779, n47581, n47571, n24068, n24067, n24066, n24065, 
        n24064, n24063, n24062, n24061, n24052, n24051, n24050, 
        n24049, n24048, n24047, n24046, n24045, n24036, n24035, 
        n24034, n24033, n24032, n24031, n24030, n24029, n24004, 
        n24003, n24002, n24001, n24000, n23999, n23998, n23997, 
        n23988, n23987, n23986, n23985, n23984, n23983, n23982, 
        n23981, n23972, n23971, n23970, n23969, n23968, n23967, 
        n23966, n23965, n224, n6837, n99, n98, n97, n96, n95, 
        n94, n93, n92, n91, n90, n89, n88, n87, n86, n85, 
        n84, n83, n82, n81, n80, n79, n78, n77, n75, n74, 
        n73, n72, n71, n70, n69, n68, n67, n66, n65, n64, 
        n63, n62, n61, n60, n59, n58, n57, n56, n55, n54, 
        n53, n25, n24, n23, n22, n21, n20, n19, n18, n17, 
        n16, n15, n14, n13, n12, n11, n10, n9, n8, n7, n6_adj_3961, 
        n5, n4_adj_3962, n3, n23940, n23939, n23938, n47557, n48782, 
        n24334, n42561, n24344, n47543, n7026, n7001, n6977, n6954, 
        n23937, n3822, n3821, n3820, n3818, n3817, n3816, n3815, 
        n3814, n3813, n3812, n3811, n3810, n3809, n3808, n3807, 
        n3806, n3805, n3804, n3803, n3802, n3801, n3800, n3799, 
        n47541, n2_adj_3963, n44238, n47539, n43909, n43907, n15_adj_3964, 
        n15_adj_3965, n2263, n2262, n2261, n4015, n2260, n2259, 
        n2258;
    wire [31:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(23[23:26])
    wire [31:0]\PID_CONTROLLER.err_prev ;   // verilog/motorControl.v(24[23:31])
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(25[23:29])
    wire [8:0]pwm_count;   // verilog/motorControl.v(55[13:22])
    
    wire n47529, n25_adj_3966, n24_adj_3967, n23_adj_3968, n22_adj_3969, 
        n21_adj_3970, n20_adj_3971, n19_adj_3972, n18_adj_3973, n17_adj_3974, 
        n16_adj_3975, n15_adj_3976, n14_adj_3977, n13_adj_3978, n12_adj_3979, 
        n11_adj_3980, n10_adj_3981, n9_adj_3982, n8_adj_3983, n7_adj_3984, 
        n6_adj_3985, n22470;
    wire [31:0]pwm_23__N_2951;
    
    wire pwm_23__N_2948, n387, n413, n414, n415, n421, n3839, 
        n48720, n455, n456, n457, n458, n459, n460, n461, n462, 
        n463, n467, n468, n469, n470, n471, n4_adj_3986, n4_adj_3987, 
        n2257, n2256, n2255, n2254, n2253, n2252, n2251, n2250, 
        n2_adj_3988, n2243, n2244, n24335, n24336, n24337, n24338, 
        n24339, n24321, n868, n869, n870, n871, n872, n873, 
        n874, n875, n24348, n24347, n23716, quadA_debounced, quadB_debounced, 
        count_enable, n49260, n47498, n47494, quadA_debounced_adj_3989, 
        quadB_debounced_adj_3990, count_enable_adj_3991, n4037, n2315, 
        n2314, n2313, n2312, n2311, n15_adj_3992, n48788, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n4_adj_3993, n47484, n2249, n24245, n24244, n24243, n23936, 
        n23935, n23934, n23933, n2248, n2247, n47478;
    wire [2:0]r_Bit_Index_adj_4419;   // verilog/uart_tx.v(33[16:27])
    
    wire n24242, n24241, n24240, n2246, n2245, n23924, n23923, 
        n23922, n23921, n23920, n23919, n2310, n2309, n2308, n2307, 
        n2306, n2305, n2304, n2303, n2302, n2301, n48875, n47471, 
        n2300, n48918;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n43905;
    wire [1:0]reg_B_adj_4426;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n2299, n6911, n47460, n24333, n47450, n48611, n47446, 
        n3_adj_3999, n47442, n43255, n369, n370, n371, n372, n373, 
        n374, n375, n376, n377, n378, n379, n380, n381, n382, 
        n383, n384, n385, n386, n387_adj_4000, n388, n389, n390, 
        n391, n392, n393, n48694, n510, n533, n534, n558, n48693, 
        n648, n649, n47434, n43253, n671, n672, n30, n6854, 
        n783, n784, n785, n806, n807, n29, n914, n915, n916, 
        n917, n918, n938, n939, n40155, n47427, n24_adj_4001, 
        n47425, n1043, n1044, n1045, n1046, n1047, n1048, n1067, 
        n1068, n47423, n23714, n23_adj_4002, n22_adj_4003, n21_adj_4004, 
        n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1193, 
        n1194, n20_adj_4005, n47419, n19_adj_4006, n1292, n1293, 
        n1294, n1295, n1296, n1297, n1298, n1299, n18_adj_4007, 
        n1316, n1317, n48887, n17_adj_4008, n6872, n1412, n1413, 
        n1414, n1415, n1416, n1417, n1418, n1419, n1420, n47411, 
        n1436, n1437, n47407, n43251, n1529, n1530, n1531, n1532, 
        n1533, n1534, n1535, n1536, n1537, n1538, n1553, n1554, 
        n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, 
        n6750, n6751, n6752, n1643, n1644, n1645, n1646, n1647, 
        n1648, n1649, n1650, n1651, n1652, n1653, n1667, n1668, 
        n1, n1754, n1755, n1756, n1757, n1758, n1759, n1760, 
        n1761, n1762, n1763, n1764, n1765, n1778, n1779, n48629, 
        n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
        n1870, n1871, n1872, n1873, n1874, n37885, n1886, n1887, 
        n37884, n37883, n37882, n6840, n6841, n6842, n6843, n6844, 
        n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, 
        n6853, n37881, n37880, n1967, n1968, n1969, n1970, n1971, 
        n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
        n1980, n1991, n1992, n37879, n6857, n6858, n6859, n6860, 
        n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, 
        n6869, n6870, n6871, n37878, n2069, n2070, n2071, n2072, 
        n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, 
        n2081, n2082, n2083, n2093, n2094, n48926, n37877, n6875, 
        n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, 
        n6884, n6885, n6886, n6887, n6888, n6889, n6890, n47396, 
        n37876, n2168, n2169, n2170, n2171, n2172, n2173, n2174, 
        n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
        n2183, n5825, n2192, n2193, n47394, n47392, n6894, n6895, 
        n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, 
        n6904, n6905, n6906, n6907, n6908, n6909, n6910, n37875, 
        n37874, n2264_adj_4009, n2265_adj_4010, n2266, n2267, n2268, 
        n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, 
        n2277, n2278, n2279, n2280, n2288, n2289, n37873, n6914, 
        n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, 
        n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, 
        n6931, n6217, n2357, n2358, n2359, n2360, n2361, n2362, 
        n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
        n2371, n2372, n2373, n2374, n2381, n2382, n20342, n6935, 
        n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, 
        n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
        n6952, n6953, n37872, n37871, n22462, n2447, n2448, n2449, 
        n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, 
        n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, 
        n2471, n2472, n37870, n6957, n6958, n6959, n6960, n6961, 
        n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, 
        n6970, n6971, n6972, n6973, n6974, n6975, n6976, n37869, 
        n6578, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
        n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, 
        n2549, n2550, n2551, n2552, n2553, n2558, n2559, n6980, 
        n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, 
        n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, 
        n6997, n6998, n6999, n7000, n5826, n2618, n2619, n2620, 
        n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, 
        n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, 
        n2637, n2638, n2642, n2643, n37868, n47386, n7004, n7005, 
        n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, 
        n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
        n7022, n7023, n7024, n7025, n37867, n2699, n2700, n2701, 
        n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, 
        n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, 
        n2718, n2719, n2720, n2723, n2724, n37866, n37865, n2777, 
        n2798, n2799, n2801, n2802, n37864, n37863, n22458, n23918, 
        n23917, n37862, n37861, n37860, n37859, n37858, n23900, 
        n37857, n23899, n23898, n23897, n23896, n23895, n23894, 
        n28052, n23893, n23892, n37856, n23891, n37855, n23890, 
        n37854, n6218, n23889, n48895, n37853, n37852, n37851, 
        n37850, n37849, n37848, n37847, n37846, n37845, n6579, 
        n37844, n37843, n37842, n37841, n37840, n37839, n47361, 
        n6649, n5827, n47357, n47355, n37838, n37837, n37836, 
        n37835, n37834, n37833, n37832, n37831, n37830, n47351, 
        n37829, n6219, n37828, n37827, n47349, n5_adj_4011, n7_adj_4012, 
        n37826, n37825, n37824, n37823, n37385, n37822, n37384, 
        n37383, n37821, n37382, n37381, n37820, n37380, n6580, 
        n37819, n37818, n37817, n6689, n22504, n6650, n43231, 
        n5828, n37816, n49155, n37815, n37814, n37813, n37812, 
        n6220, n37811, n10_adj_4013, n37810, n37809, n37808, n37807, 
        n37806, n37805, n37804, n37803, n37802, n6581, n6729, 
        n37801, n6690, n6651, n5829, n37800, n37799, n37798, n37797, 
        n37796, n37795, n37794, n37793, n37792, n37791, n37790, 
        n37789, n37788, n37787, n11_adj_4014, n13_adj_4015, n15_adj_4016, 
        n48649, n11_adj_4017, n13_adj_4018, n48725, n15_adj_4019, 
        n37786, n37785, n37784, n37783, n11_adj_4020, n13_adj_4021, 
        n15_adj_4022, n11_adj_4023, n13_adj_4024, n15_adj_4025, n1_adj_4026, 
        n47335, n22_adj_4027, n37782, n48259, n37781, n6836, n22459, 
        n37780, n37779, n4_adj_4028, n6_adj_4029, n8_adj_4030, n9_adj_4031, 
        n11_adj_4032, n13_adj_4033, n15_adj_4034, n23888, n23887, 
        n23886, n37778, n23885, n37777, n23884, n23883, n23882, 
        n37776, n23881, n37775, n23880, n23879, n23878, n23877, 
        n23875, n23874, n23873, n23872, n23871, n23870, n23869, 
        n23868, n23867, n23866, n23865, n23864, n23863, n23862, 
        n23861, n23860, n37774, n23859, n37773, n23858, n23857, 
        n23856, n23855, n48653, n23854, n37772, n23853, n23850, 
        n37771, n23849, n37770, n23846, n23845, n23844, n23840, 
        n37769, n23838, n23837, n37768, n23835, n23834, n23832, 
        n23825, n23823, n23822, n23820, n23819, n37767, n23818, 
        n23817, n23816, n23815, n37766, n23814, n23813, n23812, 
        n37765, n23809, n23806, n23803, n23799, n23797, n23796, 
        n23794, n23793, n23791, n23790, n23788, n23787, n23785, 
        n23784, n23782, n23781, n23779, n23778, n6891, n37764, 
        n37763, n37762, n47320, n10_adj_4035, n6221, n37761, n49153, 
        n37760, n37759, n37758, n6582, n6783, n37757, n6730, n6691, 
        n37756, n47318, n6652, n5830, n37755, n37754, n37753, 
        n37752, n37751, n37750, n37749, n37748, n6222, n37747, 
        n37746, n22456, n37745, n47316, n37744, n6583, n6824, 
        n37743, n6784, n6731, n37742, n8_adj_4036, n6692, n6_adj_4037, 
        n6653, n37741, n43229, n37740, n37739, n37738, n37737, 
        n47312, n37736, n47310, n37735, n6223, n4_adj_4038, n6_adj_4039, 
        n8_adj_4040, n9_adj_4041, n11_adj_4042, n13_adj_4043, n15_adj_4044, 
        n37734, n5022, n47308, n37733, n37732, n37731, n6795, 
        n6835, n23776, n47304, n37730, n37729, n6584, n37728, 
        n6825, n6785, n6732, n6693, n48905, n6654, n49149, n37727, 
        n37726, n37725, n37724, n37723, n4_adj_4045, n37722, n2_adj_4046, 
        n3_adj_4047, n4_adj_4048, n5_adj_4049, n6_adj_4050, n7_adj_4051, 
        n8_adj_4052, n9_adj_4053, n10_adj_4054, n11_adj_4055, n12_adj_4056, 
        n13_adj_4057, n14_adj_4058, n15_adj_4059, n16_adj_4060, n17_adj_4061, 
        n18_adj_4062, n19_adj_4063, n20_adj_4064, n21_adj_4065, n22_adj_4066, 
        n23_adj_4067, n24_adj_4068, n25_adj_4069, n2_adj_4070, n3_adj_4071, 
        n4_adj_4072, n5_adj_4073, n6_adj_4074, n7_adj_4075, n8_adj_4076, 
        n9_adj_4077, n10_adj_4078, n11_adj_4079, n12_adj_4080, n13_adj_4081, 
        n14_adj_4082, n15_adj_4083, n16_adj_4084, n17_adj_4085, n18_adj_4086, 
        n19_adj_4087, n20_adj_4088, n21_adj_4089, n22_adj_4090, n23_adj_4091, 
        n24_adj_4092, n25_adj_4093, n37721, n37720, n6585, n37719, 
        n6826, n6786, n6733, n6694, n37718, n6655, n37717, n37716, 
        n2_adj_4094, n37715, n37714, n37713, n37712, n37711, n37710, 
        n37709, n37708, n37707, n37706, n37705, n37704, n6827, 
        n6787, n6734, n6695, n6656, n47290, n37703, n46, n47288, 
        n37702, n37701, n37700, n37699, n37698, n37697, n37696, 
        n37695, n37694, n6828, n6788, n37693, n6735, n44, n48787, 
        n6696, n6657, n37692, n37691, n37690, n37689, n37688, 
        n37687, n37686, n47284, n37685, n37684, n42, n47282, n37683, 
        n6829, n6789, n6736, n6697, n37682, n40, n42_adj_4095, 
        n44_adj_4096, n45, n49115, n24412, n24411, n24410, n24408, 
        n24407, n37681, n38, n40_adj_4097, n42_adj_4098, n43, n48578, 
        n48967, n24406, n24405, n24404, n24403, n24402, n24401, 
        n24400, n24399, n24398, n24397, n24396, n24395, n24394, 
        n24393, n24392, n24391, n37680, n6830, n6790, n6737, n6698, 
        n24390, n37679, n36, n38_adj_4099, n40_adj_4100, n41, n49019, 
        n24388, n24385, n24384, n24383, n24382, n24381, n24380, 
        n24377, n24376, n24375, n24374, n24373, n24372, n34, n36_adj_4101, 
        n38_adj_4102, n39, n41_adj_4103, n43_adj_4104, n44_adj_4105, 
        n45_adj_4106, n48580, n24371, n24370, n24369, n24365, n24364, 
        n24363, n24362, n24359, n24358, n24357, n6831, n6791, 
        n6738, n37678, n24353, n32, n34_adj_4107, n37, n39_adj_4108, 
        n41_adj_4109, n48961, n43_adj_4110, n48582, n48959, n24352, 
        n24236, n24234, n23756, n24233, n37677, n30_adj_4111, n31, 
        n32_adj_4112, n33, n34_adj_4113, n35, n37_adj_4114, n39_adj_4115, 
        n48957, n41_adj_4116, n42_adj_4117, n43_adj_4118, n45_adj_4119, 
        n49150, n48977, n23752, n23751, n23750, n24228, n24227, 
        n24226, n6832, n6792, n28, n29_adj_4120, n30_adj_4121, n31_adj_4122, 
        n32_adj_4123, n33_adj_4124, n35_adj_4125, n37_adj_4126, n48955, 
        n39_adj_4127, n40_adj_4128, n41_adj_4129, n43_adj_4130, n48953, 
        n49135, n24225, n6739, n23746, n23602, n24223, n24222, 
        n37676, n47276, n23596, n26, n27, n28_adj_4131, n29_adj_4132, 
        n30_adj_4133, n31_adj_4134, n33_adj_4135, n35_adj_4136, n48951, 
        n37_adj_4137, n38_adj_4138, n39_adj_4139, n41_adj_4140, n49152, 
        n24221, n24220, n37675, n23745, n24_adj_4141, n25_adj_4142, 
        n26_adj_4143, n27_adj_4144, n28_adj_4145, n29_adj_4146, n30_adj_4147, 
        n31_adj_4148, n32_adj_4149, n33_adj_4150, n35_adj_4151, n36_adj_4152, 
        n37_adj_4153, n39_adj_4154, n41_adj_4155, n48813, n43_adj_4156, 
        n44_adj_4157, n45_adj_4158, n48815, n47274, n23743, n22_adj_4159, 
        n23_adj_4160, n24_adj_4161, n25_adj_4162, n26_adj_4163, n27_adj_4164, 
        n28_adj_4165, n29_adj_4166, n30_adj_4167, n31_adj_4168, n33_adj_4169, 
        n34_adj_4170, n35_adj_4171, n37_adj_4172, n39_adj_4173, n41_adj_4174, 
        n42_adj_4175, n43_adj_4176, n49119, n48943, n6833, n6793, 
        n24217, n23563, n37674, n37673, n20_adj_4177, n21_adj_4178, 
        n22_adj_4179, n23_adj_4180, n24_adj_4181, n25_adj_4182, n26_adj_4183, 
        n27_adj_4184, n28_adj_4185, n29_adj_4186, n31_adj_4187, n32_adj_4188, 
        n33_adj_4189, n35_adj_4190, n37_adj_4191, n39_adj_4192, n41_adj_4193, 
        n49231, n49160, n37672, n18_adj_4194, n19_adj_4195, n20_adj_4196, 
        n21_adj_4197, n22_adj_4198, n23_adj_4199, n24_adj_4200, n25_adj_4201, 
        n26_adj_4202, n27_adj_4203, n29_adj_4204, n30_adj_4205, n31_adj_4206, 
        n33_adj_4207, n35_adj_4208, n37_adj_4209, n49162, n39_adj_4210, 
        n41_adj_4211, n42_adj_4212, n43_adj_4213, n45_adj_4214, n48588, 
        n16_adj_4215, n17_adj_4216, n18_adj_4217, n19_adj_4218, n20_adj_4219, 
        n21_adj_4220, n22_adj_4221, n23_adj_4222, n25_adj_4223, n27_adj_4224, 
        n28_adj_4225, n29_adj_4226, n31_adj_4227, n33_adj_4228, n35_adj_4229, 
        n37_adj_4230, n39_adj_4231, n41_adj_4232, n43_adj_4233, n14_adj_4234, 
        n16_adj_4235, n17_adj_4236, n18_adj_4237, n19_adj_4238, n20_adj_4239, 
        n21_adj_4240, n22_adj_4241, n23_adj_4242, n25_adj_4243, n26_adj_4244, 
        n27_adj_4245, n29_adj_4246, n31_adj_4247, n49109, n33_adj_4248, 
        n35_adj_4249, n37_adj_4250, n39_adj_4251, n40_adj_4252, n41_adj_4253, 
        n43_adj_4254, n45_adj_4255, n49137, n23533, n12_adj_4256, 
        n14_adj_4257, n15_adj_4258, n16_adj_4259, n17_adj_4260, n18_adj_4261, 
        n19_adj_4262, n20_adj_4263, n21_adj_4264, n23_adj_4265, n24_adj_4266, 
        n25_adj_4267, n27_adj_4268, n29_adj_4269, n49111, n31_adj_4270, 
        n33_adj_4271, n35_adj_4272, n37_adj_4273, n38_adj_4274, n39_adj_4275, 
        n41_adj_4276, n48935, n43_adj_4277, n49087, n49268, n6834, 
        n6794, n10_adj_4278, n12_adj_4279, n13_adj_4280, n14_adj_4281, 
        n15_adj_4282, n16_adj_4283, n17_adj_4284, n18_adj_4285, n19_adj_4286, 
        n21_adj_4287, n22_adj_4288, n23_adj_4289, n25_adj_4290, n27_adj_4291, 
        n48974, n29_adj_4292, n48700, n31_adj_4293, n33_adj_4294, 
        n35_adj_4295, n36_adj_4296, n37_adj_4297, n39_adj_4298, n41_adj_4299, 
        n49263, n6753, n8_adj_4300, n10_adj_4301, n11_adj_4302, n12_adj_4303, 
        n13_adj_4304, n14_adj_4305, n15_adj_4306, n16_adj_4307, n17_adj_4308, 
        n19_adj_4309, n20_adj_4310, n21_adj_4311, n23_adj_4312, n25_adj_4313, 
        n48933, n27_adj_4314, n29_adj_4315, n31_adj_4316, n48931, 
        n33_adj_4317, n34_adj_4318, n35_adj_4319, n37_adj_4320, n39_adj_4321, 
        n48845, n49164, n48847, n37671, n6_adj_4322, n8_adj_4323, 
        n9_adj_4324, n10_adj_4325, n11_adj_4326, n12_adj_4327, n13_adj_4328, 
        n14_adj_4329, n15_adj_4330, n17_adj_4331, n19_adj_4332, n21_adj_4333, 
        n23_adj_4334, n48851, n25_adj_4335, n48927, n27_adj_4336, 
        n29_adj_4337, n48925, n31_adj_4338, n32_adj_4339, n33_adj_4340, 
        n35_adj_4341, n37_adj_4342, n49166, n49117, n48921, n4_adj_4343, 
        n6_adj_4344, n7_adj_4345, n8_adj_4346, n9_adj_4347, n10_adj_4348, 
        n11_adj_4349, n12_adj_4350, n13_adj_4351, n15_adj_4352, n16_adj_4353, 
        n17_adj_4354, n19_adj_4355, n21_adj_4356, n48919, n23_adj_4357, 
        n24_adj_4358, n25_adj_4359, n27_adj_4360, n48917, n29_adj_4361, 
        n30_adj_4362, n31_adj_4363, n33_adj_4364, n35_adj_4365, n48867, 
        n37_adj_4366, n49043, n39_adj_4367, n40_adj_4368, n41_adj_4369, 
        n43_adj_4370, n45_adj_4371, n49045, n37670, n48714, n37669, 
        n37668, n47266, n37667, n37666, n37665, n37664, n47258, 
        n37663, n37662, n37661, n37660, n47252, n37659, n37658, 
        n37657, n37656, n37655, n49121, n37654, n37653, n47236, 
        n37652, n45225, n37651, n48778, n37650, n37649, n37648, 
        n48747, n37647, n47225, n37646, n37645, n37644, n37643, 
        n37642, n37641, n37640, n37639, n37638, n37637, n22833, 
        n48749, n28350, n22561, n22558, n22555, n44576, n22429, 
        n37221, n37220, n37219, n37218, n37217, n47207, n47206, 
        n44626, n22467, n37606, n37605, n37604, n37603, n37602, 
        n1_adj_4372, n24346, n37601, n24345, n37600, n47647, n48928, 
        n7_adj_4373, n50101, n24343, n24342, n24341, n43236, n24340, 
        n47188, n47186, n47184, n48544, n47182, n47180, n49256, 
        n49254, n49248, n48777, n49247, n49267, n49232, n49220, 
        n49249, n47157, n47156, n49212, n49255, n49253, n49251, 
        n49217, n49191, n49190, n49229, n49173, n49172, n48785, 
        n49169, n49120, n49118, n49116, n49112, n49110, n49108, 
        n49102, n49098, n49096, n49094, n49158, n49090, n44902, 
        n5_adj_4374, n42011, n49265, n48781, n49034, n49028, n49156, 
        n49154, n44586, n48993, n49107, n48980, n48976, n48972, 
        n49113, n48968, n48964, n48962, n48960, n48958, n48956, 
        n48952, n48936, n48934, n48932, n48864, n48862, n48854, 
        n48850, n48842, n48840, n48835, n48833, n48789, n48808, 
        n42279, n49148, n48415, n48574, n48411, n48401, n48586, 
        n5_adj_4375, n48589, n48365, n43709, n49961, n41_adj_4376, 
        n40_adj_4377, n44311, n43459, n43441, n48710, n48317, n48273, 
        n48709, n48265, n48242, n48240, n48236, n48234, n48228, 
        n48226, n48218, n48216, n48200, n48197, n48715, n48186, 
        n48176, n48704, n48171, n48116, n48703, n48096, n48613, 
        n48040, n48032, n47972, n48804, n48633, n48699, n48802, 
        n49258, n48798, n48963, n48508, n49161;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n2291({n2292, n2293, n2294, 
            n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
            n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
            n2311, n2312, n2313, n2314, n2315}), .encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .data_o({quadA_debounced, quadB_debounced}), 
            .clk32MHz(clk32MHz), .n23875(n23875), .n23874(n23874), .n23873(n23873), 
            .n23872(n23872), .n23871(n23871), .n23870(n23870), .n23869(n23869), 
            .n23868(n23868), .n23867(n23867), .n23866(n23866), .n23865(n23865), 
            .n23864(n23864), .n23863(n23863), .n23862(n23862), .n23861(n23861), 
            .n23860(n23860), .n23859(n23859), .n23858(n23858), .n23857(n23857), 
            .n23856(n23856), .n23855(n23855), .n23854(n23854), .n23850(n23850), 
            .n23745(n23745), .count_enable(count_enable), .n24359(n24359), 
            .reg_B({reg_B}), .PIN_23_c_1(PIN_23_c_1), .PIN_24_c_0(PIN_24_c_0), 
            .n23750(n23750), .n44902(n44902)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(166[15] 171[4])
    SB_IO hall1_input (.PACKAGE_PIN(PIN_20), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall2_input (.PACKAGE_PIN(PIN_21), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_22), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_3024_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n37701), 
            .O(n6852)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31812_4_lut (.I0(n33_adj_4189), .I1(n31_adj_4187), .I2(n29_adj_4186), 
            .I3(n47320), .O(n47312));
    defparam i31812_4_lut.LUT_INIT = 16'haaab;
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3024_4 (.CI(n37701), .I0(n1979), .I1(n98), .CO(n37702));
    SB_LUT4 add_3024_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n37700), 
            .O(n6853)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_3 (.CI(n37700), .I0(n1980), .I1(n99), .CO(n37701));
    motorControl control (.GND_net(GND_net), .\PWMLimit[4] (PWMLimit[4]), 
            .\PWMLimit[0] (PWMLimit[0]), .\PWMLimit[1] (PWMLimit[1]), .\PID_CONTROLLER.result[5] (\PID_CONTROLLER.result [5]), 
            .n11(n11_adj_4020), .\PID_CONTROLLER.result[6] (\PID_CONTROLLER.result [6]), 
            .n13(n13_adj_4021), .\PID_CONTROLLER.result[7] (\PID_CONTROLLER.result [7]), 
            .n15(n15_adj_4022), .\PWMLimit[8] (PWMLimit[8]), .\PWMLimit[9] (PWMLimit[9]), 
            .\PID_CONTROLLER.err[31] (\PID_CONTROLLER.err [31]), .n387(n387), 
            .n11_adj_10(n11_adj_4017), .n24384(n24384), .pwm({pwm}), .clk32MHz(clk32MHz), 
            .n24383(n24383), .n24382(n24382), .n24381(n24381), .n24380(n24380), 
            .n42011(n42011), .n24377(n24377), .n24376(n24376), .n24375(n24375), 
            .n24374(n24374), .n24373(n24373), .n24372(n24372), .n24371(n24371), 
            .n24370(n24370), .n24369(n24369), .n24365(n24365), .n24364(n24364), 
            .n24363(n24363), .n24362(n24362), .n24358(n24358), .\deadband[9] (deadband[9]), 
            .\pwm_23__N_2951[5] (pwm_23__N_2951[5]), .\pwm_23__N_2951[6] (pwm_23__N_2951[6]), 
            .n13_adj_11(n13_adj_4018), .n15_adj_12(n15_adj_4019), .\pwm_23__N_2951[7] (pwm_23__N_2951[7]), 
            .pwm_23__N_2948(pwm_23__N_2948), .\Ki[7] (Ki[7]), .\Ki[3] (Ki[3]), 
            .\Kp[1] (Kp[1]), .\PID_CONTROLLER.err[7] (\PID_CONTROLLER.err [7]), 
            .\Kp[0] (Kp[0]), .\PID_CONTROLLER.err[8] (\PID_CONTROLLER.err [8]), 
            .\Kp[2] (Kp[2]), .n11_adj_13(n11_adj_4023), .\Kp[3] (Kp[3]), 
            .\PID_CONTROLLER.err[3] (\PID_CONTROLLER.err [3]), .\PID_CONTROLLER.err[13] (\PID_CONTROLLER.err [13]), 
            .n415(n415), .n414(n414), .n13_adj_14(n13_adj_4024), .\PID_CONTROLLER.err[14] (\PID_CONTROLLER.err [14]), 
            .\deadband[0] (deadband[0]), .n15_adj_15(n15_adj_4025), .\PID_CONTROLLER.err[0] (\PID_CONTROLLER.err [0]), 
            .PIN_7_c_1(PIN_7_c_1), .n413(n413), .\Kp[4] (Kp[4]), .n421(n421), 
            .\Ki[4] (Ki[4]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), .\Ki[5] (Ki[5]), 
            .\Kp[7] (Kp[7]), .\Kd[1] (Kd[1]), .\Kd[0] (Kd[0]), .VCC_net(VCC_net), 
            .\Ki[6] (Ki[6]), .\Kd[2] (Kd[2]), .\Kd[3] (Kd[3]), .\Kd[4] (Kd[4]), 
            .\deadband[1] (deadband[1]), .\Kd[5] (Kd[5]), .\Kd[6] (Kd[6]), 
            .\Kd[7] (Kd[7]), .\Ki[0] (Ki[0]), .\deadband[2] (deadband[2]), 
            .\deadband[3] (deadband[3]), .\deadband[4] (deadband[4]), .\Ki[1] (Ki[1]), 
            .\PID_CONTROLLER.err[9] (\PID_CONTROLLER.err [9]), .\PID_CONTROLLER.err[6] (\PID_CONTROLLER.err [6]), 
            .\PID_CONTROLLER.err[5] (\PID_CONTROLLER.err [5]), .\PID_CONTROLLER.err[4] (\PID_CONTROLLER.err [4]), 
            .\PID_CONTROLLER.err[2] (\PID_CONTROLLER.err [2]), .\PID_CONTROLLER.err[1] (\PID_CONTROLLER.err [1]), 
            .pwm_count({pwm_count}), .\Ki[2] (Ki[2]), .\deadband[5] (deadband[5]), 
            .\deadband[6] (deadband[6]), .\deadband[7] (deadband[7]), .\deadband[8] (deadband[8]), 
            .\PID_CONTROLLER.err[19] (\PID_CONTROLLER.err [19]), .\PID_CONTROLLER.err[20] (\PID_CONTROLLER.err [20]), 
            .\PID_CONTROLLER.err[18] (\PID_CONTROLLER.err [18]), .\PID_CONTROLLER.err[17] (\PID_CONTROLLER.err [17]), 
            .IntegralLimit({IntegralLimit}), .\motor_state[23] (motor_state[23]), 
            .\motor_state[22] (motor_state[22]), .\motor_state[21] (motor_state[21]), 
            .\motor_state[20] (motor_state[20]), .\motor_state[19] (motor_state[19]), 
            .\motor_state[18] (motor_state[18]), .\motor_state[17] (motor_state[17]), 
            .\motor_state[16] (motor_state[16]), .\motor_state[15] (motor_state[15]), 
            .\motor_state[14] (motor_state[14]), .\PID_CONTROLLER.err[22] (\PID_CONTROLLER.err [22]), 
            .\PID_CONTROLLER.err[23] (\PID_CONTROLLER.err [23]), .\motor_state[13] (motor_state[13]), 
            .\motor_state[12] (motor_state[12]), .\motor_state[11] (motor_state[11]), 
            .\motor_state[10] (motor_state[10]), .\motor_state[9] (motor_state[9]), 
            .\motor_state[8] (motor_state[8]), .\motor_state[7] (motor_state[7]), 
            .\motor_state[6] (motor_state[6]), .\motor_state[5] (motor_state[5]), 
            .\motor_state[4] (motor_state[4]), .\motor_state[3] (motor_state[3]), 
            .\motor_state[2] (motor_state[2]), .\motor_state[1] (motor_state[1]), 
            .\PID_CONTROLLER.err[12] (\PID_CONTROLLER.err [12]), .\motor_state[0] (motor_state[0]), 
            .\PID_CONTROLLER.err_prev[31] (\PID_CONTROLLER.err_prev [31]), 
            .\PID_CONTROLLER.err_prev[23] (\PID_CONTROLLER.err_prev [23]), 
            .\PID_CONTROLLER.err_prev[22] (\PID_CONTROLLER.err_prev [22]), 
            .\PID_CONTROLLER.err_prev[21] (\PID_CONTROLLER.err_prev [21]), 
            .\PID_CONTROLLER.err_prev[20] (\PID_CONTROLLER.err_prev [20]), 
            .\PID_CONTROLLER.err_prev[19] (\PID_CONTROLLER.err_prev [19]), 
            .\PID_CONTROLLER.err_prev[18] (\PID_CONTROLLER.err_prev [18]), 
            .\PID_CONTROLLER.err_prev[17] (\PID_CONTROLLER.err_prev [17]), 
            .\PID_CONTROLLER.err_prev[16] (\PID_CONTROLLER.err_prev [16]), 
            .\PID_CONTROLLER.err_prev[15] (\PID_CONTROLLER.err_prev [15]), 
            .\PID_CONTROLLER.err_prev[14] (\PID_CONTROLLER.err_prev [14]), 
            .\PID_CONTROLLER.err_prev[13] (\PID_CONTROLLER.err_prev [13]), 
            .\PID_CONTROLLER.err_prev[12] (\PID_CONTROLLER.err_prev [12]), 
            .\PID_CONTROLLER.err_prev[11] (\PID_CONTROLLER.err_prev [11]), 
            .\PID_CONTROLLER.err_prev[10] (\PID_CONTROLLER.err_prev [10]), 
            .\PID_CONTROLLER.err_prev[9] (\PID_CONTROLLER.err_prev [9]), .\PID_CONTROLLER.err_prev[8] (\PID_CONTROLLER.err_prev [8]), 
            .\PID_CONTROLLER.err_prev[7] (\PID_CONTROLLER.err_prev [7]), .\PID_CONTROLLER.err_prev[6] (\PID_CONTROLLER.err_prev [6]), 
            .\PID_CONTROLLER.err_prev[5] (\PID_CONTROLLER.err_prev [5]), .\PID_CONTROLLER.err_prev[4] (\PID_CONTROLLER.err_prev [4]), 
            .\PID_CONTROLLER.err_prev[3] (\PID_CONTROLLER.err_prev [3]), .\PID_CONTROLLER.err_prev[2] (\PID_CONTROLLER.err_prev [2]), 
            .\PID_CONTROLLER.err_prev[1] (\PID_CONTROLLER.err_prev [1]), .\PID_CONTROLLER.err_prev[0] (\PID_CONTROLLER.err_prev [0]), 
            .n22(n22_adj_4003), .n21(n21_adj_4004), .n23900(n23900), .n23899(n23899), 
            .n23898(n23898), .n23897(n23897), .n23896(n23896), .n23895(n23895), 
            .n23894(n23894), .n23893(n23893), .n23892(n23892), .n23891(n23891), 
            .n23890(n23890), .n23889(n23889), .n24(n24_adj_4001), .n23888(n23888), 
            .n23887(n23887), .n23886(n23886), .n23885(n23885), .n23884(n23884), 
            .n23883(n23883), .n23882(n23882), .n23881(n23881), .n23880(n23880), 
            .n23879(n23879), .n23878(n23878), .n20(n20_adj_4005), .n23877(n23877), 
            .n23(n23_adj_4002), .n19(n19_adj_4006), .n17(n17_adj_4008), 
            .n48782(n48782), .n18(n18_adj_4007), .PIN_8_c_2(PIN_8_c_2), 
            .PIN_9_c_3(PIN_9_c_3), .PIN_10_c_4(PIN_10_c_4), .PIN_11_c_5(PIN_11_c_5), 
            .n868(n868), .\PID_CONTROLLER.err[10] (\PID_CONTROLLER.err [10]), 
            .\PID_CONTROLLER.err[11] (\PID_CONTROLLER.err [11]), .\PID_CONTROLLER.err[15] (\PID_CONTROLLER.err [15]), 
            .\PID_CONTROLLER.err[16] (\PID_CONTROLLER.err [16]), .\PID_CONTROLLER.err[21] (\PID_CONTROLLER.err [21]), 
            .n869(n869), .n870(n870), .n871(n871), .PIN_6_c_0(PIN_6_c_0), 
            .n872(n872), .n873(n873), .n874(n874), .n875(n875), .n47156(n47156), 
            .n23743(n23743), .\PWMLimit[2] (PWMLimit[2]), .\PWMLimit[3] (PWMLimit[3]), 
            .hall3(hall3), .\PWMLimit[5] (PWMLimit[5]), .hall1(hall1), 
            .\PWMLimit[6] (PWMLimit[6]), .hall2(hall2), .\PWMLimit[7] (PWMLimit[7]), 
            .n29(n29), .n30(n30), .n48778(n48778), .n471(n471), .n470(n470), 
            .n469(n469), .n468(n468), .n467(n467), .n1(n1_adj_4026), 
            .n28052(n28052), .n1_adj_16(n1), .n463(n463), .n44626(n44626), 
            .n462(n462), .n461(n461), .n460(n460), .n459(n459), .n458(n458), 
            .n457(n457), .n456(n456), .n455(n455), .n15_adj_17(n15_adj_4016), 
            .n13_adj_18(n13_adj_4015), .n11_adj_19(n11_adj_4014), .setpoint({setpoint}), 
            .n47225(n47225), .n47180(n47180), .n47182(n47182), .n47188(n47188), 
            .n47186(n47186), .n47184(n47184)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(143[16] 159[4])
    SB_LUT4 add_3024_2_lut (.I0(GND_net), .I1(n382), .I2(n558), .I3(VCC_net), 
            .O(n6854)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_2_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_10_pad (.PACKAGE_PIN(PIN_10), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_10_c_4)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_10_pad.PIN_TYPE = 6'b011001;
    defparam PIN_10_pad.PULLUP = 1'b0;
    defparam PIN_10_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_10_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3024_2 (.CI(VCC_net), .I0(n382), .I1(n558), .CO(n37700));
    SB_LUT4 add_3023_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n37699), 
            .O(n6824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3023_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n37698), 
            .O(n6825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1350_i20_4_lut (.I0(n383), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4177));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_1350_i28_3_lut (.I0(n26_adj_4183), .I1(n93), 
            .I2(n31_adj_4187), .I3(GND_net), .O(n28_adj_4185));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1463_3_lut_3_lut (.I0(n2192), .I1(n6879), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1462_3_lut_3_lut (.I0(n2192), .I1(n6878), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3023_14 (.CI(n37698), .I0(n1863), .I1(n88), .CO(n37699));
    SB_LUT4 div_12_i1461_3_lut_3_lut (.I0(n2192), .I1(n6877), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1350_i32_3_lut (.I0(n24_adj_4181), .I1(n91), 
            .I2(n35_adj_4190), .I3(GND_net), .O(n32_adj_4188));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3023_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n37697), 
            .O(n6826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33654_4_lut (.I0(n32_adj_4188), .I1(n22_adj_4179), .I2(n35_adj_4190), 
            .I3(n47310), .O(n49156));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33654_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3023_13 (.CI(n37697), .I0(n1864), .I1(n89), .CO(n37698));
    SB_LUT4 div_12_i1464_3_lut_3_lut (.I0(n2192), .I1(n6880), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33655_3_lut (.I0(n49156), .I1(n90), .I2(n37_adj_4191), .I3(GND_net), 
            .O(n49157));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33655_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33592_3_lut (.I0(n49157), .I1(n89), .I2(n39_adj_4192), .I3(GND_net), 
            .O(n49094));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33592_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3023_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n37696), 
            .O(n6827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33223_4_lut (.I0(n39_adj_4192), .I1(n37_adj_4191), .I2(n35_adj_4190), 
            .I3(n47312), .O(n48725));
    defparam i33223_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33656_4_lut (.I0(n28_adj_4185), .I1(n20_adj_4177), .I2(n31_adj_4187), 
            .I3(n47316), .O(n49158));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33656_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3023_12 (.CI(n37696), .I0(n1865), .I1(n90), .CO(n37697));
    SB_LUT4 i33526_3_lut (.I0(n49094), .I1(n88), .I2(n41_adj_4193), .I3(GND_net), 
            .O(n49028));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33526_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1472_3_lut_3_lut (.I0(n2192), .I1(n6888), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3023_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n37695), 
            .O(n6828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1473_3_lut_3_lut (.I0(n2192), .I1(n6889), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3023_11 (.CI(n37695), .I0(n1866), .I1(n91), .CO(n37696));
    SB_LUT4 div_12_i1471_3_lut_3_lut (.I0(n2192), .I1(n6887), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33729_4_lut (.I0(n49028), .I1(n49158), .I2(n41_adj_4193), 
            .I3(n48725), .O(n49231));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33729_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33730_3_lut (.I0(n49231), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n49232));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33730_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33667_3_lut (.I0(n49232), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n49169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33667_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_3023_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n37694), 
            .O(n6829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_10 (.CI(n37694), .I0(n1867), .I1(n92), .CO(n37695));
    SB_LUT4 i1_4_lut (.I0(n49169), .I1(n22543), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1470_3_lut_3_lut (.I0(n2192), .I1(n6886), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1469_3_lut_3_lut (.I0(n2192), .I1(n6885), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1468_3_lut_3_lut (.I0(n2192), .I1(n6884), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1527_3_lut_3_lut (.I0(n2288), .I1(n6899), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i6_2_lut (.I0(pwm_23__N_2951[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4018));   // verilog/motorControl.v(25[23:29])
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_2_lut (.I0(pwm_23__N_2951[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4017));   // verilog/motorControl.v(25[23:29])
    defparam i14_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3023_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n37693), 
            .O(n6830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_9 (.CI(n37693), .I0(n1868), .I1(n93), .CO(n37694));
    SB_LUT4 add_3023_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n37692), 
            .O(n6831)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_8 (.CI(n37692), .I0(n1869), .I1(n94), .CO(n37693));
    SB_LUT4 add_3023_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n37691), 
            .O(n6832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_7 (.CI(n37691), .I0(n1870), .I1(n95), .CO(n37692));
    SB_LUT4 div_12_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4176));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3023_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n37690), 
            .O(n6833)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_6 (.CI(n37690), .I0(n1871), .I1(n96), .CO(n37691));
    SB_LUT4 i21_2_lut (.I0(PWMLimit[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4022));   // verilog/motorControl.v(25[23:29])
    defparam i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3023_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n37689), 
            .O(n6834)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_5 (.CI(n37689), .I0(n1872), .I1(n97), .CO(n37690));
    SB_LUT4 add_3023_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n37688), 
            .O(n6835)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_4 (.CI(n37688), .I0(n1873), .I1(n98), .CO(n37689));
    SB_LUT4 add_3023_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n37687), 
            .O(n6836)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_3 (.CI(n37687), .I0(n1874), .I1(n99), .CO(n37688));
    SB_LUT4 add_3023_2_lut (.I0(GND_net), .I1(n381), .I2(n558), .I3(VCC_net), 
            .O(n6837)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3023_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3023_2 (.CI(VCC_net), .I0(n381), .I1(n558), .CO(n37687));
    SB_LUT4 div_12_i1522_3_lut_3_lut (.I0(n2288), .I1(n6894), .I2(n2264_adj_4009), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3021_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n37686), 
            .O(n6783)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3021_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n37685), 
            .O(n6784)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_13 (.CI(n37685), .I0(n1755), .I1(n89), .CO(n37686));
    SB_LUT4 add_3021_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n37684), 
            .O(n6785)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_12 (.CI(n37684), .I0(n1756), .I1(n90), .CO(n37685));
    SB_LUT4 add_3021_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n37683), 
            .O(n6786)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_11 (.CI(n37683), .I0(n1757), .I1(n91), .CO(n37684));
    SB_LUT4 add_3021_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n37682), 
            .O(n6787)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_2_lut (.I0(PWMLimit[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4021));   // verilog/motorControl.v(25[23:29])
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1525_3_lut_3_lut (.I0(n2288), .I1(n6897), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3021_10 (.CI(n37682), .I0(n1758), .I1(n92), .CO(n37683));
    SB_LUT4 add_3021_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n37681), 
            .O(n6788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_2_lut (.I0(PWMLimit[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4020));   // verilog/motorControl.v(25[23:29])
    defparam i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3021_9 (.CI(n37681), .I0(n1759), .I1(n93), .CO(n37682));
    SB_LUT4 add_3021_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n37680), 
            .O(n6789)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_8 (.CI(n37680), .I0(n1760), .I1(n94), .CO(n37681));
    SB_LUT4 add_3021_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n37679), 
            .O(n6790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_7 (.CI(n37679), .I0(n1761), .I1(n95), .CO(n37680));
    SB_LUT4 add_3021_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n37678), 
            .O(n6791)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_6 (.CI(n37678), .I0(n1762), .I1(n96), .CO(n37679));
    SB_LUT4 add_3021_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n37677), 
            .O(n6792)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2986_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n37221), 
            .O(n5825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3021_5 (.CI(n37677), .I0(n1763), .I1(n97), .CO(n37678));
    SB_LUT4 add_3021_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n37676), 
            .O(n6793)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_4 (.CI(n37676), .I0(n1764), .I1(n98), .CO(n37677));
    SB_LUT4 div_12_i1523_3_lut_3_lut (.I0(n2288), .I1(n6895), .I2(n2265_adj_4010), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3021_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n37675), 
            .O(n6794)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_3 (.CI(n37675), .I0(n1765), .I1(n99), .CO(n37676));
    SB_LUT4 add_3021_2_lut (.I0(GND_net), .I1(n380), .I2(n558), .I3(VCC_net), 
            .O(n6795)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3021_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3021_2 (.CI(VCC_net), .I0(n380), .I1(n558), .CO(n37675));
    SB_LUT4 add_3019_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n37674), 
            .O(n6742)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3019_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n37673), 
            .O(n6743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_12 (.CI(n37673), .I0(n1644), .I1(n90), .CO(n37674));
    SB_LUT4 div_12_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3019_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n37672), 
            .O(n6744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_11 (.CI(n37672), .I0(n1645), .I1(n91), .CO(n37673));
    SB_LUT4 add_3019_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n37671), 
            .O(n6745)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_10 (.CI(n37671), .I0(n1646), .I1(n92), .CO(n37672));
    SB_LUT4 add_3019_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n37670), 
            .O(n6746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_9 (.CI(n37670), .I0(n1647), .I1(n93), .CO(n37671));
    SB_LUT4 add_3019_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n37669), 
            .O(n6747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_8 (.CI(n37669), .I0(n1648), .I1(n94), .CO(n37670));
    SB_LUT4 add_3019_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n37668), 
            .O(n6748)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_7 (.CI(n37668), .I0(n1649), .I1(n95), .CO(n37669));
    SB_LUT4 add_3019_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n37667), 
            .O(n6749)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_6 (.CI(n37667), .I0(n1650), .I1(n96), .CO(n37668));
    SB_LUT4 add_3019_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n37666), 
            .O(n6750)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_5 (.CI(n37666), .I0(n1651), .I1(n97), .CO(n37667));
    SB_LUT4 add_3019_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n37665), 
            .O(n6751)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_4 (.CI(n37665), .I0(n1652), .I1(n98), .CO(n37666));
    SB_LUT4 add_3019_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n37664), 
            .O(n6752)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3019_3 (.CI(n37664), .I0(n1653), .I1(n99), .CO(n37665));
    SB_LUT4 add_3019_2_lut (.I0(GND_net), .I1(n379), .I2(n558), .I3(VCC_net), 
            .O(n6753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3019_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1526_3_lut_3_lut (.I0(n2288), .I1(n6898), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3019_2 (.CI(VCC_net), .I0(n379), .I1(n558), .CO(n37664));
    SB_LUT4 add_3018_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n37663), 
            .O(n6729)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3018_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n37662), 
            .O(n6730)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_11 (.CI(n37662), .I0(n1530), .I1(n91), .CO(n37663));
    SB_LUT4 add_3018_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n37661), 
            .O(n6731)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_10 (.CI(n37661), .I0(n1531), .I1(n92), .CO(n37662));
    SB_LUT4 add_3018_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n37660), 
            .O(n6732)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_9 (.CI(n37660), .I0(n1532), .I1(n93), .CO(n37661));
    SB_LUT4 add_3018_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n37659), 
            .O(n6733)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_8 (.CI(n37659), .I0(n1533), .I1(n94), .CO(n37660));
    SB_LUT4 add_3018_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n37658), 
            .O(n6734)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_7 (.CI(n37658), .I0(n1534), .I1(n95), .CO(n37659));
    SB_LUT4 add_3018_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n37657), 
            .O(n6735)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_6 (.CI(n37657), .I0(n1535), .I1(n96), .CO(n37658));
    SB_LUT4 add_3018_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n37656), 
            .O(n6736)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1338_3_lut_3_lut (.I0(n1991), .I1(n6851), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3018_5 (.CI(n37656), .I0(n1536), .I1(n97), .CO(n37657));
    SB_LUT4 add_3018_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n37655), 
            .O(n6737)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_4 (.CI(n37655), .I0(n1537), .I1(n98), .CO(n37656));
    SB_LUT4 add_3018_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n37654), 
            .O(n6738)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_3 (.CI(n37654), .I0(n1538), .I1(n99), .CO(n37655));
    SB_LUT4 add_3018_2_lut (.I0(GND_net), .I1(n378), .I2(n558), .I3(VCC_net), 
            .O(n6739)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3018_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3018_2 (.CI(VCC_net), .I0(n378), .I1(n558), .CO(n37654));
    SB_LUT4 add_3016_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n37653), 
            .O(n6689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3016_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n37652), 
            .O(n6690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_10 (.CI(n37652), .I0(n1413), .I1(n92), .CO(n37653));
    SB_LUT4 add_3016_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n37651), 
            .O(n6691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_9 (.CI(n37651), .I0(n1414), .I1(n93), .CO(n37652));
    SB_LUT4 add_3016_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n37650), 
            .O(n6692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_8 (.CI(n37650), .I0(n1415), .I1(n94), .CO(n37651));
    SB_LUT4 add_3016_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n37649), 
            .O(n6693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_7 (.CI(n37649), .I0(n1416), .I1(n95), .CO(n37650));
    SB_LUT4 add_3016_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n37648), 
            .O(n6694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_6 (.CI(n37648), .I0(n1417), .I1(n96), .CO(n37649));
    SB_LUT4 add_3016_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n37647), 
            .O(n6695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_5 (.CI(n37647), .I0(n1418), .I1(n97), .CO(n37648));
    SB_LUT4 add_3016_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n37646), 
            .O(n6696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_4 (.CI(n37646), .I0(n1419), .I1(n98), .CO(n37647));
    SB_LUT4 add_3016_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n37645), 
            .O(n6697)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_3 (.CI(n37645), .I0(n1420), .I1(n99), .CO(n37646));
    SB_LUT4 add_3016_2_lut (.I0(GND_net), .I1(n377), .I2(n558), .I3(VCC_net), 
            .O(n6698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3016_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3016_2 (.CI(VCC_net), .I0(n377), .I1(n558), .CO(n37645));
    SB_LUT4 div_12_i1535_3_lut_3_lut (.I0(n2288), .I1(n6907), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_906_i32_4_lut (.I0(n377), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_i1532_3_lut_3_lut (.I0(n2288), .I1(n6904), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3014_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n37644), 
            .O(n6649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3014_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n37643), 
            .O(n6650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_9 (.CI(n37643), .I0(n1293), .I1(n93), .CO(n37644));
    SB_LUT4 add_3014_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n37642), 
            .O(n6651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1531_3_lut_3_lut (.I0(n2288), .I1(n6903), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1530_3_lut_3_lut (.I0(n2288), .I1(n6902), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3014_8 (.CI(n37642), .I0(n1294), .I1(n94), .CO(n37643));
    SB_LUT4 add_3014_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n37641), 
            .O(n6652)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1529_3_lut_3_lut (.I0(n2288), .I1(n6901), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1528_3_lut_3_lut (.I0(n2288), .I1(n6900), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3014_7 (.CI(n37641), .I0(n1295), .I1(n95), .CO(n37642));
    SB_LUT4 add_3014_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n37640), 
            .O(n6653)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4162));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4164));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1524_3_lut_3_lut (.I0(n2288), .I1(n6896), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3014_6 (.CI(n37640), .I0(n1296), .I1(n96), .CO(n37641));
    SB_LUT4 add_3014_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n37639), 
            .O(n6654)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_5 (.CI(n37639), .I0(n1297), .I1(n97), .CO(n37640));
    SB_LUT4 add_3014_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n37638), 
            .O(n6655)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_4 (.CI(n37638), .I0(n1298), .I1(n98), .CO(n37639));
    SB_LUT4 add_3014_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n37637), 
            .O(n6656)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_3 (.CI(n37637), .I0(n1299), .I1(n99), .CO(n37638));
    SB_LUT4 add_3014_2_lut (.I0(GND_net), .I1(n376), .I2(n558), .I3(VCC_net), 
            .O(n6657)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3014_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3014_2 (.CI(VCC_net), .I0(n376), .I1(n558), .CO(n37637));
    SB_LUT4 div_12_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4166));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3011_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n37606), 
            .O(n6578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3011_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n37605), 
            .O(n6579)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_8 (.CI(n37605), .I0(n1170), .I1(n94), .CO(n37606));
    SB_LUT4 add_3011_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n37604), 
            .O(n6580)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1539_3_lut_3_lut (.I0(n2288), .I1(n6911), .I2(n385), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3011_7 (.CI(n37604), .I0(n1171), .I1(n95), .CO(n37605));
    SB_LUT4 add_3011_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n37603), 
            .O(n6581)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_6 (.CI(n37603), .I0(n1172), .I1(n96), .CO(n37604));
    SB_LUT4 add_3011_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n37602), 
            .O(n6582)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_5 (.CI(n37602), .I0(n1173), .I1(n97), .CO(n37603));
    SB_LUT4 add_3011_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n37601), 
            .O(n6583)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4168));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3011_4 (.CI(n37601), .I0(n1174), .I1(n98), .CO(n37602));
    SB_LUT4 add_3011_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n37600), 
            .O(n6584)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_3 (.CI(n37600), .I0(n1175), .I1(n99), .CO(n37601));
    SB_LUT4 add_3011_2_lut (.I0(GND_net), .I1(n375), .I2(n558), .I3(VCC_net), 
            .O(n6585)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3011_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3011_2 (.CI(VCC_net), .I0(n375), .I1(n558), .CO(n37600));
    SB_LUT4 div_12_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1534_3_lut_3_lut (.I0(n2288), .I1(n6906), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1335_3_lut_3_lut (.I0(n1991), .I1(n6848), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4160));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31861_4_lut (.I0(n29_adj_4166), .I1(n27_adj_4164), .I2(n25_adj_4162), 
            .I3(n23_adj_4160), .O(n47361));
    defparam i31861_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_i1533_3_lut_3_lut (.I0(n2288), .I1(n6905), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1538_3_lut_3_lut (.I0(n2288), .I1(n6910), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1536_3_lut_3_lut (.I0(n2288), .I1(n6908), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31851_4_lut (.I0(n35_adj_4171), .I1(n33_adj_4169), .I2(n31_adj_4168), 
            .I3(n47361), .O(n47351));
    defparam i31851_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2986_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n37220), 
            .O(n5826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1537_3_lut_3_lut (.I0(n2288), .I1(n6909), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1281_i22_4_lut (.I0(n382), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4159));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_1281_i30_3_lut (.I0(n28_adj_4165), .I1(n93), 
            .I2(n33_adj_4169), .I3(GND_net), .O(n30_adj_4167));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1281_i34_3_lut (.I0(n26_adj_4163), .I1(n91), 
            .I2(n37_adj_4172), .I3(GND_net), .O(n34_adj_4170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1595_3_lut_3_lut (.I0(n2381), .I1(n6926), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2986_6 (.CI(n37220), .I0(n915), .I1(n96), .CO(n37221));
    SB_LUT4 i33652_4_lut (.I0(n34_adj_4170), .I1(n24_adj_4161), .I2(n37_adj_4172), 
            .I3(n47349), .O(n49154));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33652_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33653_3_lut (.I0(n49154), .I1(n90), .I2(n39_adj_4173), .I3(GND_net), 
            .O(n49155));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33653_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33594_3_lut (.I0(n49155), .I1(n89), .I2(n41_adj_4174), .I3(GND_net), 
            .O(n49096));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33594_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33245_4_lut (.I0(n41_adj_4174), .I1(n39_adj_4173), .I2(n37_adj_4172), 
            .I3(n47351), .O(n48747));
    defparam i33245_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33441_4_lut (.I0(n30_adj_4167), .I1(n22_adj_4159), .I2(n33_adj_4169), 
            .I3(n47355), .O(n48943));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33441_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33524_3_lut (.I0(n49096), .I1(n88), .I2(n43_adj_4176), .I3(GND_net), 
            .O(n42_adj_4175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33524_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i16_2_lut (.I0(n413), .I1(\PID_CONTROLLER.result [7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4025));   // verilog/motorControl.v(25[23:29])
    defparam i16_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_i1583_3_lut_3_lut (.I0(n2381), .I1(n6914), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33615_4_lut (.I0(n42_adj_4175), .I1(n48943), .I2(n43_adj_4176), 
            .I3(n48747), .O(n49117));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33615_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33616_3_lut (.I0(n49117), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n49118));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33616_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1449 (.I0(n49118), .I1(n22540), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1449.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_3999));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10919_3_lut (.I0(encoder1_position[4]), .I1(n2261), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24334));   // quad.v(35[10] 41[6])
    defparam i10919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1584_3_lut_3_lut (.I0(n2381), .I1(n6915), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_2_lut (.I0(n414), .I1(\PID_CONTROLLER.result [6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4024));   // verilog/motorControl.v(25[23:29])
    defparam i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i16_2_lut_adj_1450 (.I0(n415), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4023));   // verilog/motorControl.v(25[23:29])
    defparam i16_2_lut_adj_1450.LUT_INIT = 16'h6666;
    SB_LUT4 i10827_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24242));   // verilog/coms.v(125[12] 284[6])
    defparam i10827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(n84), .I1(n22546), .I2(GND_net), .I3(GND_net), 
            .O(n22543));
    defparam i1_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_IO PIN_18_pad (.PACKAGE_PIN(PIN_18), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_18_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_18_pad.PIN_TYPE = 6'b000001;
    defparam PIN_18_pad.PULLUP = 1'b0;
    defparam PIN_18_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_18_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_12_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2986_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n37219), 
            .O(n5827)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1587_3_lut_3_lut (.I0(n2381), .I1(n6918), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2986_5 (.CI(n37219), .I0(n916), .I1(n97), .CO(n37220));
    SB_LUT4 add_2986_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n37218), 
            .O(n5828)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1336_3_lut_3_lut (.I0(n1991), .I1(n6849), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1588_3_lut_3_lut (.I0(n2381), .I1(n6919), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1585_3_lut_3_lut (.I0(n2381), .I1(n6916), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1586_3_lut_3_lut (.I0(n2381), .I1(n6917), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10969_4_lut (.I0(pwm_23__N_2948), .I1(n47188), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24384));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10969_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 div_12_i1601_3_lut_3_lut (.I0(n2381), .I1(n6932), .I2(n386), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1597_3_lut_3_lut (.I0(n2381), .I1(n6928), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_2986_4 (.CI(n37218), .I0(n917), .I1(n98), .CO(n37219));
    SB_LUT4 add_2986_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n37217), 
            .O(n5829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_3 (.CI(n37217), .I0(n918), .I1(n99), .CO(n37218));
    SB_LUT4 add_2986_2_lut (.I0(GND_net), .I1(n373), .I2(n558), .I3(VCC_net), 
            .O(n5830)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2986_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2986_2 (.CI(VCC_net), .I0(n373), .I1(n558), .CO(n37217));
    SB_LUT4 div_12_i1599_3_lut_3_lut (.I0(n2381), .I1(n6930), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10970_3_lut (.I0(quadA_debounced_adj_3989), .I1(reg_B_adj_4426[1]), 
            .I2(n44576), .I3(GND_net), .O(n24385));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1593_3_lut_3_lut (.I0(n2381), .I1(n6924), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1594_3_lut_3_lut (.I0(n2381), .I1(n6925), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1592_3_lut_3_lut (.I0(n2381), .I1(n6923), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1591_3_lut_3_lut (.I0(n2381), .I1(n6922), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1590_3_lut_3_lut (.I0(n2381), .I1(n6921), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10973_4_lut (.I0(n29726), .I1(byte_transmit_counter[0]), .I2(n2241), 
            .I3(n3839), .O(n24388));   // verilog/coms.v(125[12] 284[6])
    defparam i10973_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_12_i1589_3_lut_3_lut (.I0(n2381), .I1(n6920), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1596_3_lut_3_lut (.I0(n2381), .I1(n6927), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_1[0]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_LUT4 i10975_3_lut (.I0(setpoint[1]), .I1(n3800), .I2(n23533), .I3(GND_net), 
            .O(n24390));   // verilog/coms.v(125[12] 284[6])
    defparam i10975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1600_3_lut_3_lut (.I0(n2381), .I1(n6931), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i10976_3_lut (.I0(setpoint[2]), .I1(n3801), .I2(n23533), .I3(GND_net), 
            .O(n24391));   // verilog/coms.v(125[12] 284[6])
    defparam i10976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1598_3_lut_3_lut (.I0(n2381), .I1(n6929), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10977_3_lut (.I0(setpoint[3]), .I1(n3802), .I2(n23533), .I3(GND_net), 
            .O(n24392));   // verilog/coms.v(125[12] 284[6])
    defparam i10977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1655_3_lut_3_lut (.I0(n2471), .I1(n6948), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4070), .I3(n38028), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_12_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4071), .I3(n38027), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_24 (.CI(n38027), .I0(GND_net), .I1(n3_adj_4071), 
            .CO(n38028));
    SB_LUT4 div_12_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4072), .I3(n38026), .O(n4_adj_3962)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_23 (.CI(n38026), .I0(GND_net), .I1(n4_adj_4072), 
            .CO(n38027));
    SB_LUT4 div_12_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4073), .I3(n38025), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_22 (.CI(n38025), .I0(GND_net), .I1(n5_adj_4073), 
            .CO(n38026));
    SB_LUT4 div_12_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4074), .I3(n38024), .O(n6_adj_3961)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_21 (.CI(n38024), .I0(GND_net), .I1(n6_adj_4074), 
            .CO(n38025));
    SB_LUT4 div_12_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4075), .I3(n38023), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_20 (.CI(n38023), .I0(GND_net), .I1(n7_adj_4075), 
            .CO(n38024));
    SB_LUT4 div_12_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4076), .I3(n38022), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_19 (.CI(n38022), .I0(GND_net), .I1(n8_adj_4076), 
            .CO(n38023));
    SB_LUT4 div_12_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4077), .I3(n38021), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_18 (.CI(n38021), .I0(GND_net), .I1(n9_adj_4077), 
            .CO(n38022));
    SB_LUT4 div_12_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4078), .I3(n38020), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_17 (.CI(n38020), .I0(GND_net), .I1(n10_adj_4078), 
            .CO(n38021));
    SB_LUT4 div_12_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4079), .I3(n38019), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_16 (.CI(n38019), .I0(GND_net), .I1(n11_adj_4079), 
            .CO(n38020));
    SB_LUT4 i10978_3_lut (.I0(setpoint[4]), .I1(n3803), .I2(n23533), .I3(GND_net), 
            .O(n24393));   // verilog/coms.v(125[12] 284[6])
    defparam i10978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4080), .I3(n38018), .O(n12)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_15 (.CI(n38018), .I0(GND_net), .I1(n12_adj_4080), 
            .CO(n38019));
    SB_LUT4 div_12_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4081), .I3(n38017), .O(n13)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_14 (.CI(n38017), .I0(GND_net), .I1(n13_adj_4081), 
            .CO(n38018));
    SB_LUT4 div_12_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4082), .I3(n38016), .O(n14)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_13 (.CI(n38016), .I0(GND_net), .I1(n14_adj_4082), 
            .CO(n38017));
    SB_LUT4 i10979_3_lut (.I0(setpoint[5]), .I1(n3804), .I2(n23533), .I3(GND_net), 
            .O(n24394));   // verilog/coms.v(125[12] 284[6])
    defparam i10979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4083), .I3(n38015), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_11_pad (.PACKAGE_PIN(PIN_11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_11_c_5)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_11_pad.PIN_TYPE = 6'b011001;
    defparam PIN_11_pad.PULLUP = 1'b0;
    defparam PIN_11_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_23_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b000001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i10980_3_lut (.I0(setpoint[6]), .I1(n3805), .I2(n23533), .I3(GND_net), 
            .O(n24395));   // verilog/coms.v(125[12] 284[6])
    defparam i10980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10981_3_lut (.I0(setpoint[7]), .I1(n3806), .I2(n23533), .I3(GND_net), 
            .O(n24396));   // verilog/coms.v(125[12] 284[6])
    defparam i10981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10982_3_lut (.I0(setpoint[8]), .I1(n3807), .I2(n23533), .I3(GND_net), 
            .O(n24397));   // verilog/coms.v(125[12] 284[6])
    defparam i10982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10983_3_lut (.I0(setpoint[9]), .I1(n3808), .I2(n23533), .I3(GND_net), 
            .O(n24398));   // verilog/coms.v(125[12] 284[6])
    defparam i10983_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1643_3_lut_3_lut (.I0(n2471), .I1(n6936), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1642_3_lut_3_lut (.I0(n2471), .I1(n6935), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10984_3_lut (.I0(setpoint[10]), .I1(n3809), .I2(n23533), 
            .I3(GND_net), .O(n24399));   // verilog/coms.v(125[12] 284[6])
    defparam i10984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33459_3_lut (.I0(n32), .I1(n95), .I2(n39_adj_4108), .I3(GND_net), 
            .O(n48961));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33459_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1644_3_lut_3_lut (.I0(n2471), .I1(n6937), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10985_3_lut (.I0(setpoint[11]), .I1(n3810), .I2(n23533), 
            .I3(GND_net), .O(n24400));   // verilog/coms.v(125[12] 284[6])
    defparam i10985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1647_3_lut_3_lut (.I0(n2471), .I1(n6940), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1645_3_lut_3_lut (.I0(n2471), .I1(n6938), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10986_3_lut (.I0(setpoint[12]), .I1(n3811), .I2(n23533), 
            .I3(GND_net), .O(n24401));   // verilog/coms.v(125[12] 284[6])
    defparam i10986_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_12_unary_minus_2_add_3_12 (.CI(n38015), .I0(GND_net), .I1(n15_adj_4083), 
            .CO(n38016));
    SB_LUT4 i2_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22467), .O(n248));
    defparam i2_4_lut.LUT_INIT = 16'hff37;
    SB_LUT4 div_12_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4084), .I3(n38014), .O(n16)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_11 (.CI(n38014), .I0(GND_net), .I1(n16_adj_4084), 
            .CO(n38015));
    SB_LUT4 div_12_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4085), .I3(n38013), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_10 (.CI(n38013), .I0(GND_net), .I1(n17_adj_4085), 
            .CO(n38014));
    SB_LUT4 div_12_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4086), .I3(n38012), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1648_3_lut_3_lut (.I0(n2471), .I1(n6941), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_12_unary_minus_2_add_3_9 (.CI(n38012), .I0(GND_net), .I1(n18_adj_4086), 
            .CO(n38013));
    SB_LUT4 i34461_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n49961));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i34461_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i10987_3_lut (.I0(setpoint[13]), .I1(n3812), .I2(n23533), 
            .I3(GND_net), .O(n24402));   // verilog/coms.v(125[12] 284[6])
    defparam i10987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4087), .I3(n38011), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_8 (.CI(n38011), .I0(GND_net), .I1(n19_adj_4087), 
            .CO(n38012));
    SB_LUT4 i10988_3_lut (.I0(setpoint[14]), .I1(n3813), .I2(n23533), 
            .I3(GND_net), .O(n24403));   // verilog/coms.v(125[12] 284[6])
    defparam i10988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4088), .I3(n38010), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_7 (.CI(n38010), .I0(GND_net), .I1(n20_adj_4088), 
            .CO(n38011));
    SB_LUT4 div_12_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4089), .I3(n38009), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10989_3_lut (.I0(setpoint[15]), .I1(n3814), .I2(n23533), 
            .I3(GND_net), .O(n24404));   // verilog/coms.v(125[12] 284[6])
    defparam i10989_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_12_unary_minus_2_add_3_6 (.CI(n38009), .I0(GND_net), .I1(n21_adj_4089), 
            .CO(n38010));
    SB_LUT4 div_12_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4090), .I3(n38008), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_5 (.CI(n38008), .I0(GND_net), .I1(n22_adj_4090), 
            .CO(n38009));
    SB_LUT4 div_12_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4091), .I3(n38007), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10990_3_lut (.I0(setpoint[16]), .I1(n3815), .I2(n23533), 
            .I3(GND_net), .O(n24405));   // verilog/coms.v(125[12] 284[6])
    defparam i10990_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_12_unary_minus_2_add_3_4 (.CI(n38007), .I0(GND_net), .I1(n23_adj_4091), 
            .CO(n38008));
    SB_LUT4 div_12_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4092), .I3(n38006), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_2_add_3_3 (.CI(n38006), .I0(GND_net), .I1(n24_adj_4092), 
            .CO(n38007));
    SB_LUT4 div_12_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4093), .I3(VCC_net), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10991_3_lut (.I0(setpoint[17]), .I1(n3816), .I2(n23533), 
            .I3(GND_net), .O(n24406));   // verilog/coms.v(125[12] 284[6])
    defparam i10991_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_12_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4093), 
            .CO(n38006));
    SB_LUT4 div_12_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4046), .I3(n38005), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_12_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4047), .I3(n38004), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10992_3_lut (.I0(setpoint[18]), .I1(n3817), .I2(n23533), 
            .I3(GND_net), .O(n24407));   // verilog/coms.v(125[12] 284[6])
    defparam i10992_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_12_unary_minus_4_add_3_24 (.CI(n38004), .I0(GND_net), .I1(n3_adj_4047), 
            .CO(n38005));
    SB_LUT4 div_12_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4048), .I3(n38003), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_9_pad (.PACKAGE_PIN(PIN_9), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_9_c_3)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_9_pad.PIN_TYPE = 6'b011001;
    defparam PIN_9_pad.PULLUP = 1'b0;
    defparam PIN_9_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_9_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c_2)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i10993_3_lut (.I0(setpoint[19]), .I1(n3818), .I2(n23533), 
            .I3(GND_net), .O(n24408));   // verilog/coms.v(125[12] 284[6])
    defparam i10993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32163_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[14] [4]), 
            .I2(n47), .I3(\FRAME_MATCHER.state [1]), .O(n47236));   // verilog/coms.v(125[12] 284[6])
    defparam i32163_4_lut.LUT_INIT = 16'hcacc;
    SB_LUT4 div_12_i1661_3_lut_3_lut (.I0(n2471), .I1(n6954), .I2(n387_adj_4000), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i24_3_lut (.I0(setpoint[20]), .I1(n47236), .I2(n23533), .I3(GND_net), 
            .O(n42279));   // verilog/coms.v(125[12] 284[6])
    defparam i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1646_3_lut_3_lut (.I0(n2471), .I1(n6939), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10995_3_lut (.I0(setpoint[21]), .I1(n3820), .I2(n23533), 
            .I3(GND_net), .O(n24410));   // verilog/coms.v(125[12] 284[6])
    defparam i10995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10996_3_lut (.I0(setpoint[22]), .I1(n3821), .I2(n23533), 
            .I3(GND_net), .O(n24411));   // verilog/coms.v(125[12] 284[6])
    defparam i10996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1650_3_lut_3_lut (.I0(n2471), .I1(n6943), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1651_3_lut_3_lut (.I0(n2471), .I1(n6944), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1649_3_lut_3_lut (.I0(n2471), .I1(n6942), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_12_unary_minus_4_add_3_23 (.CI(n38003), .I0(GND_net), .I1(n4_adj_4048), 
            .CO(n38004));
    SB_LUT4 i33460_3_lut (.I0(n48961), .I1(n94), .I2(n41_adj_4109), .I3(GND_net), 
            .O(n48962));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33460_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1658_3_lut_3_lut (.I0(n2471), .I1(n6951), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i968_3_lut (.I0(n1418), .I1(n6695), .I2(n1436), .I3(GND_net), 
            .O(n1535));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1659_3_lut_3_lut (.I0(n2471), .I1(n6952), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4049), .I3(n38002), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1653_3_lut_3_lut (.I0(n2471), .I1(n6946), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1654_3_lut_3_lut (.I0(n2471), .I1(n6947), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1652_3_lut_3_lut (.I0(n2471), .I1(n6945), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_12_unary_minus_4_add_3_22 (.CI(n38002), .I0(GND_net), .I1(n5_adj_4049), 
            .CO(n38003));
    SB_LUT4 i10997_3_lut (.I0(setpoint[23]), .I1(n3822), .I2(n23533), 
            .I3(GND_net), .O(n24412));   // verilog/coms.v(125[12] 284[6])
    defparam i10997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1657_3_lut_3_lut (.I0(n2471), .I1(n6950), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1656_3_lut_3_lut (.I0(n2471), .I1(n6949), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4050), .I3(n38001), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_21 (.CI(n38001), .I0(GND_net), .I1(n6_adj_4050), 
            .CO(n38002));
    SB_LUT4 div_12_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4051), .I3(n38000), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_20 (.CI(n38000), .I0(GND_net), .I1(n7_adj_4051), 
            .CO(n38001));
    SB_LUT4 div_12_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4052), .I3(n37999), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_19 (.CI(n37999), .I0(GND_net), .I1(n8_adj_4052), 
            .CO(n38000));
    SB_LUT4 div_12_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4053), .I3(n37998), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_18 (.CI(n37998), .I0(GND_net), .I1(n9_adj_4053), 
            .CO(n37999));
    SB_LUT4 div_12_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4054), .I3(n37997), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1660_3_lut_3_lut (.I0(n2471), .I1(n6953), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_12_unary_minus_4_add_3_17 (.CI(n37997), .I0(GND_net), .I1(n10_adj_4054), 
            .CO(n37998));
    SB_LUT4 div_12_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4055), .I3(n37996), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_16 (.CI(n37996), .I0(GND_net), .I1(n11_adj_4055), 
            .CO(n37997));
    SB_LUT4 i10397_4_lut (.I0(n23714), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n23596), .O(n23812));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10397_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4056), .I3(n37995), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_15 (.CI(n37995), .I0(GND_net), .I1(n12_adj_4056), 
            .CO(n37996));
    SB_LUT4 div_12_i1712_3_lut_3_lut (.I0(n2558), .I1(n6970), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1700_3_lut_3_lut (.I0(n2558), .I1(n6958), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1699_3_lut_3_lut (.I0(n2558), .I1(n6957), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4057), .I3(n37994), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1702_3_lut_3_lut (.I0(n2558), .I1(n6960), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_12_unary_minus_4_add_3_14 (.CI(n37994), .I0(GND_net), .I1(n13_adj_4057), 
            .CO(n37995));
    SB_LUT4 div_12_i1701_3_lut_3_lut (.I0(n2558), .I1(n6959), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1705_3_lut_3_lut (.I0(n2558), .I1(n6963), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4058), .I3(n37993), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_13 (.CI(n37993), .I0(GND_net), .I1(n14_adj_4058), 
            .CO(n37994));
    SB_LUT4 div_12_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4059), .I3(n37992), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_12 (.CI(n37992), .I0(GND_net), .I1(n15_adj_4059), 
            .CO(n37993));
    SB_LUT4 div_12_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4060), .I3(n37991), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_11 (.CI(n37991), .I0(GND_net), .I1(n16_adj_4060), 
            .CO(n37992));
    SB_LUT4 div_12_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4061), .I3(n37990), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_10 (.CI(n37990), .I0(GND_net), .I1(n17_adj_4061), 
            .CO(n37991));
    SB_LUT4 div_12_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4062), .I3(n37989), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_9 (.CI(n37989), .I0(GND_net), .I1(n18_adj_4062), 
            .CO(n37990));
    SB_LUT4 div_12_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4063), .I3(n37988), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_8 (.CI(n37988), .I0(GND_net), .I1(n19_adj_4063), 
            .CO(n37989));
    SB_LUT4 div_12_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4064), .I3(n37987), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_7 (.CI(n37987), .I0(GND_net), .I1(n20_adj_4064), 
            .CO(n37988));
    SB_LUT4 div_12_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4065), .I3(n37986), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_6 (.CI(n37986), .I0(GND_net), .I1(n21_adj_4065), 
            .CO(n37987));
    SB_LUT4 div_12_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4066), .I3(n37985), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1045_3_lut (.I0(n1535), .I1(n6735), .I2(n1553), .I3(GND_net), 
            .O(n1649));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_12_unary_minus_4_add_3_5 (.CI(n37985), .I0(GND_net), .I1(n22_adj_4066), 
            .CO(n37986));
    SB_LUT4 div_12_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4067), .I3(n37984), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_4 (.CI(n37984), .I0(GND_net), .I1(n23_adj_4067), 
            .CO(n37985));
    SB_LUT4 div_12_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4068), .I3(n37983), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_12_unary_minus_4_add_3_3 (.CI(n37983), .I0(GND_net), .I1(n24_adj_4068), 
            .CO(n37984));
    SB_LUT4 div_12_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4069), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_12_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1703_3_lut_3_lut (.I0(n2558), .I1(n6961), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1706_3_lut_3_lut (.I0(n2558), .I1(n6964), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1120_3_lut (.I0(n1649), .I1(n6748), .I2(n1667), .I3(GND_net), 
            .O(n1760));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1120_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY div_12_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4069), 
            .CO(n37983));
    SB_LUT4 i10394_4_lut (.I0(n23714), .I1(r_Bit_Index[2]), .I2(n4015), 
            .I3(n23596), .O(n23809));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10394_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_i1719_3_lut_3_lut (.I0(n2558), .I1(n6977), .I2(n388), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1193_3_lut (.I0(n1760), .I1(n6789), .I2(n1778), .I3(GND_net), 
            .O(n1868));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n380));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32060_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n47157));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32060_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i10391_4_lut (.I0(n23716), .I1(r_Bit_Index_adj_4419[1]), .I2(r_Bit_Index_adj_4419[0]), 
            .I3(n23602), .O(n23806));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10391_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_i1704_3_lut_3_lut (.I0(n2558), .I1(n6962), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1709_3_lut_3_lut (.I0(n2558), .I1(n6967), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1451 (.I0(n47157), .I1(n22467), .I2(n99), .I3(n5_adj_4374), 
            .O(n392));
    defparam i1_4_lut_adj_1451.LUT_INIT = 16'hefce;
    SB_LUT4 div_12_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10388_4_lut (.I0(n23716), .I1(r_Bit_Index_adj_4419[2]), .I2(n4037), 
            .I3(n23602), .O(n23803));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10388_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_12_i1708_3_lut_3_lut (.I0(n2558), .I1(n6966), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10384_2_lut (.I0(n23845), .I1(n23797), .I2(GND_net), .I3(GND_net), 
            .O(n23799));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10384_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1717_3_lut_3_lut (.I0(n2558), .I1(n6975), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10381_2_lut (.I0(n23845), .I1(n23794), .I2(GND_net), .I3(GND_net), 
            .O(n23796));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10381_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10378_2_lut (.I0(n23845), .I1(n23791), .I2(GND_net), .I3(GND_net), 
            .O(n23793));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10378_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10375_2_lut (.I0(n23845), .I1(n23788), .I2(GND_net), .I3(GND_net), 
            .O(n23790));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10372_2_lut (.I0(n23845), .I1(n23785), .I2(GND_net), .I3(GND_net), 
            .O(n23787));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10372_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10369_2_lut (.I0(n23845), .I1(n23782), .I2(GND_net), .I3(GND_net), 
            .O(n23784));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10366_2_lut (.I0(n23845), .I1(n23779), .I2(GND_net), .I3(GND_net), 
            .O(n23781));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10366_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32674_4_lut (.I0(n41_adj_4109), .I1(n39_adj_4108), .I2(n37), 
            .I3(n47529), .O(n48176));
    defparam i32674_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_i1718_3_lut_3_lut (.I0(n2558), .I1(n6976), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10363_2_lut (.I0(n23845), .I1(n23776), .I2(GND_net), .I3(GND_net), 
            .O(n23778));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_12_i1713_3_lut_3_lut (.I0(n2558), .I1(n6971), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1715_3_lut_3_lut (.I0(n2558), .I1(n6973), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1716_3_lut_3_lut (.I0(n2558), .I1(n6974), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1711_3_lut_3_lut (.I0(n2558), .I1(n6969), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1710_3_lut_3_lut (.I0(n2558), .I1(n6968), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2999_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n37385), 
            .O(n6217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2999_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n37384), 
            .O(n6218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_7 (.CI(n37384), .I0(n1044), .I1(n95), .CO(n37385));
    SB_LUT4 add_2999_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n37383), 
            .O(n6219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_6 (.CI(n37383), .I0(n1045), .I1(n96), .CO(n37384));
    SB_LUT4 div_12_i1714_3_lut_3_lut (.I0(n2558), .I1(n6972), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2999_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n37382), 
            .O(n6220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_5 (.CI(n37382), .I0(n1046), .I1(n97), .CO(n37383));
    SB_LUT4 div_12_i1707_3_lut_3_lut (.I0(n2558), .I1(n6965), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1768_3_lut_3_lut (.I0(n2642), .I1(n6994), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2999_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n37381), 
            .O(n6221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_4 (.CI(n37381), .I0(n1047), .I1(n98), .CO(n37382));
    SB_LUT4 add_2999_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n37380), 
            .O(n6222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_3 (.CI(n37380), .I0(n1048), .I1(n99), .CO(n37381));
    SB_LUT4 div_12_i1754_3_lut_3_lut (.I0(n2642), .I1(n6980), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_2999_2_lut (.I0(GND_net), .I1(n374), .I2(n558), .I3(VCC_net), 
            .O(n6223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2999_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2999_2 (.CI(VCC_net), .I0(n374), .I1(n558), .CO(n37380));
    SB_LUT4 div_12_i1755_3_lut_3_lut (.I0(n2642), .I1(n6981), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14660_3_lut (.I0(n20342), .I1(rx_data[7]), .I2(\data_in_frame[7] [7]), 
            .I3(GND_net), .O(n24029));   // verilog/coms.v(88[13:20])
    defparam i14660_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1756_3_lut_3_lut (.I0(n2642), .I1(n6982), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10615_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n20342), 
            .I3(GND_net), .O(n24030));   // verilog/coms.v(125[12] 284[6])
    defparam i10615_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1758_3_lut_3_lut (.I0(n2642), .I1(n6984), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1757_3_lut_3_lut (.I0(n2642), .I1(n6983), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1761_3_lut_3_lut (.I0(n2642), .I1(n6987), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1762_3_lut_3_lut (.I0(n2642), .I1(n6988), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10616_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n20342), 
            .I3(GND_net), .O(n24031));   // verilog/coms.v(125[12] 284[6])
    defparam i10616_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1114_3_lut (.I0(n1643), .I1(n6742), .I2(n1667), .I3(GND_net), 
            .O(n1754));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1187_3_lut (.I0(n1754), .I1(n6783), .I2(n1778), .I3(GND_net), 
            .O(n1862));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i725_3_lut (.I0(n374), .I1(n6223), .I2(n1067), .I3(GND_net), 
            .O(n1175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i808_3_lut (.I0(n1175), .I1(n6584), .I2(n1193), .I3(GND_net), 
            .O(n1298));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i808_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i889_3_lut (.I0(n1298), .I1(n6655), .I2(n1316), .I3(GND_net), 
            .O(n1418));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_297_i46_4_lut (.I0(n370), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1452 (.I0(n46), .I1(n22504), .I2(n98), .I3(n43905), 
            .O(n533));
    defparam i1_4_lut_adj_1452.LUT_INIT = 16'hefce;
    SB_LUT4 i23056_2_lut (.I0(n370), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3963));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23056_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32317_3_lut (.I0(n369), .I1(n558), .I2(n392), .I3(GND_net), 
            .O(n510));
    defparam i32317_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_12_LessThan_390_i44_4_lut (.I0(n371), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33283_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n48785));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33283_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i10617_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n20342), 
            .I3(GND_net), .O(n24032));   // verilog/coms.v(125[12] 284[6])
    defparam i10617_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33078_3_lut (.I0(n34_adj_4107), .I1(n96), .I2(n37), .I3(GND_net), 
            .O(n48580));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33078_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10618_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n20342), 
            .I3(GND_net), .O(n24033));   // verilog/coms.v(125[12] 284[6])
    defparam i10618_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3033_25_lut (.I0(n249), .I1(n49961), .I2(n248), .I3(n37885), 
            .O(displacement_23__N_91[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_25_lut.LUT_INIT = 16'h8BB8;
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_7_c_1)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b011001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i1_4_lut_adj_1453 (.I0(n48785), .I1(n22507), .I2(n97), .I3(n43907), 
            .O(n671));
    defparam i1_4_lut_adj_1453.LUT_INIT = 16'hefce;
    SB_LUT4 div_12_i368_4_lut (.I0(n510), .I1(n2_adj_3963), .I2(n533), 
            .I3(n99), .O(n648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i368_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_481_i42_4_lut (.I0(n372), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33285_3_lut (.I0(n42), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n48787));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33285_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33286_3_lut (.I0(n48787), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n48788));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33286_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1454 (.I0(n48788), .I1(n22510), .I2(n96), .I3(n43909), 
            .O(n806));
    defparam i1_4_lut_adj_1454.LUT_INIT = 16'hefce;
    SB_LUT4 i23128_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4045), .I3(GND_net), 
            .O(n6_adj_4037));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23128_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_12_i459_4_lut (.I0(n648), .I1(n4), .I2(n671), .I3(n98), 
            .O(n783));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i459_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_LessThan_570_i40_4_lut (.I0(n373), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_LessThan_570_i44_3_lut (.I0(n42_adj_4095), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4096));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33287_4_lut (.I0(n44_adj_4096), .I1(n40), .I2(n45), .I3(n47589), 
            .O(n48789));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33287_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1455 (.I0(n48789), .I1(n22513), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1455.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i548_4_lut (.I0(n783), .I1(n6_adj_4037), .I2(n806), 
            .I3(n97), .O(n915));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i548_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_i1759_3_lut_3_lut (.I0(n2642), .I1(n6985), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3033_24_lut (.I0(n393), .I1(n49961), .I2(n392), .I3(n37884), 
            .O(displacement_23__N_91[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_24 (.CI(n37884), .I0(n49961), .I1(n392), .CO(n37885));
    SB_LUT4 i10619_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n20342), 
            .I3(GND_net), .O(n24034));   // verilog/coms.v(125[12] 284[6])
    defparam i10619_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1760_3_lut_3_lut (.I0(n2642), .I1(n6986), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1775_3_lut_3_lut (.I0(n2642), .I1(n7001), .I2(n389), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1765_3_lut_3_lut (.I0(n2642), .I1(n6991), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3033_23_lut (.I0(n534), .I1(n49961), .I2(n533), .I3(n37883), 
            .O(displacement_23__N_91[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_23 (.CI(n37883), .I0(n49961), .I1(n533), .CO(n37884));
    SB_LUT4 div_12_i1764_3_lut_3_lut (.I0(n2642), .I1(n6990), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10620_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n20342), 
            .I3(GND_net), .O(n24035));   // verilog/coms.v(125[12] 284[6])
    defparam i10620_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1773_3_lut_3_lut (.I0(n2642), .I1(n6999), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_657_i38_4_lut (.I0(n374), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3033_22_lut (.I0(n672), .I1(n49961), .I2(n671), .I3(n37882), 
            .O(displacement_23__N_91[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i10835_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24250));   // verilog/coms.v(125[12] 284[6])
    defparam i10835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_657_i42_3_lut (.I0(n40_adj_4097), .I1(n96), 
            .I2(n43), .I3(GND_net), .O(n42_adj_4098));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33465_4_lut (.I0(n42_adj_4098), .I1(n38), .I2(n43), .I3(n47571), 
            .O(n48967));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33465_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33466_3_lut (.I0(n48967), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n48968));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33466_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY add_3033_22 (.CI(n37882), .I0(n49961), .I1(n671), .CO(n37883));
    SB_LUT4 i1_4_lut_adj_1456 (.I0(n48968), .I1(n22516), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1456.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1774_3_lut_3_lut (.I0(n2642), .I1(n7000), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3033_21_lut (.I0(n807), .I1(n49961), .I2(n806), .I3(n37881), 
            .O(displacement_23__N_91[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_21 (.CI(n37881), .I0(n49961), .I1(n806), .CO(n37882));
    SB_LUT4 add_3033_20_lut (.I0(n939), .I1(n49961), .I2(n938), .I3(n37880), 
            .O(displacement_23__N_91[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_20 (.CI(n37880), .I0(n49961), .I1(n938), .CO(n37881));
    SB_LUT4 add_3033_19_lut (.I0(n1068), .I1(n49961), .I2(n1067), .I3(n37879), 
            .O(displacement_23__N_91[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_19 (.CI(n37879), .I0(n49961), .I1(n1067), .CO(n37880));
    SB_LUT4 add_3033_18_lut (.I0(n1194), .I1(n49961), .I2(n1193), .I3(n37878), 
            .O(displacement_23__N_91[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_18 (.CI(n37878), .I0(n49961), .I1(n1193), .CO(n37879));
    SB_LUT4 div_12_i635_3_lut (.I0(n915), .I1(n5826), .I2(n938), .I3(GND_net), 
            .O(n1044));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i635_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3033_17_lut (.I0(n1317), .I1(n49961), .I2(n1316), .I3(n37877), 
            .O(displacement_23__N_91[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_17 (.CI(n37877), .I0(n49961), .I1(n1316), .CO(n37878));
    SB_LUT4 add_3033_16_lut (.I0(n1437), .I1(n49961), .I2(n1436), .I3(n37876), 
            .O(displacement_23__N_91[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_16 (.CI(n37876), .I0(n49961), .I1(n1436), .CO(n37877));
    SB_LUT4 i10920_3_lut (.I0(encoder1_position[5]), .I1(n2260), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24335));   // quad.v(35[10] 41[6])
    defparam i10920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3033_15_lut (.I0(n1554), .I1(n49961), .I2(n1553), .I3(n37875), 
            .O(displacement_23__N_91[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_15 (.CI(n37875), .I0(n49961), .I1(n1553), .CO(n37876));
    SB_LUT4 add_3033_14_lut (.I0(n1668), .I1(n49961), .I2(n1667), .I3(n37874), 
            .O(displacement_23__N_91[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_14 (.CI(n37874), .I0(n49961), .I1(n1667), .CO(n37875));
    SB_LUT4 add_3033_13_lut (.I0(n1779), .I1(n49961), .I2(n1778), .I3(n37873), 
            .O(displacement_23__N_91[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i10836_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24251));   // verilog/coms.v(125[12] 284[6])
    defparam i10836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10621_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n20342), 
            .I3(GND_net), .O(n24036));   // verilog/coms.v(125[12] 284[6])
    defparam i10621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1766_3_lut_3_lut (.I0(n2642), .I1(n6992), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10837_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24252));   // verilog/coms.v(125[12] 284[6])
    defparam i10837_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3033_13 (.CI(n37873), .I0(n49961), .I1(n1778), .CO(n37874));
    SB_LUT4 i10838_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24253));   // verilog/coms.v(125[12] 284[6])
    defparam i10838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3033_12_lut (.I0(n1887), .I1(n49961), .I2(n1886), .I3(n37872), 
            .O(displacement_23__N_91[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_12_i1767_3_lut_3_lut (.I0(n2642), .I1(n6993), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4069));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4068));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1772_3_lut_3_lut (.I0(n2642), .I1(n6998), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_742_i36_4_lut (.I0(n375), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_i1770_3_lut_3_lut (.I0(n2642), .I1(n6996), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4067));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4066));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4065));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1334_3_lut_3_lut (.I0(n1991), .I1(n6847), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4064));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1769_3_lut_3_lut (.I0(n2642), .I1(n6995), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_91[23]), 
            .I2(n3_adj_3999), .I3(n37168), .O(displacement_23__N_1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_742_i40_3_lut (.I0(n38_adj_4099), .I1(n96), 
            .I2(n41), .I3(GND_net), .O(n40_adj_4100));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33646_4_lut (.I0(n40_adj_4100), .I1(n36), .I2(n41), .I3(n47557), 
            .O(n49148));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33646_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33647_3_lut (.I0(n49148), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n49149));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33647_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33600_3_lut (.I0(n49149), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n49102));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33600_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1457 (.I0(n49102), .I1(n22519), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1457.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i720_3_lut (.I0(n1044), .I1(n6218), .I2(n1067), .I3(GND_net), 
            .O(n1170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_825_i34_4_lut (.I0(n376), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY add_3033_12 (.CI(n37872), .I0(n49961), .I1(n1886), .CO(n37873));
    SB_LUT4 i33461_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4103), .I3(GND_net), 
            .O(n48963));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33461_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33462_3_lut (.I0(n48963), .I1(n94), .I2(n43_adj_4104), .I3(GND_net), 
            .O(n48964));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33462_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32684_4_lut (.I0(n43_adj_4104), .I1(n41_adj_4103), .I2(n39), 
            .I3(n47543), .O(n48186));
    defparam i32684_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_91[22]), 
            .I2(n3_adj_3999), .I3(n37167), .O(displacement_23__N_1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_825_i38_3_lut (.I0(n36_adj_4101), .I1(n96), 
            .I2(n39), .I3(GND_net), .O(n38_adj_4102));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3033_11_lut (.I0(n1992), .I1(n49961), .I2(n1991), .I3(n37871), 
            .O(displacement_23__N_91[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i33294_3_lut (.I0(n48964), .I1(n93), .I2(n45_adj_4106), .I3(GND_net), 
            .O(n44_adj_4105));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33294_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n37167), .I0(displacement_23__N_91[22]), 
            .I1(n3_adj_3999), .CO(n37168));
    SB_LUT4 i33076_4_lut (.I0(n44_adj_4105), .I1(n38_adj_4102), .I2(n45_adj_4106), 
            .I3(n48186), .O(n48578));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33076_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1458 (.I0(n48578), .I1(n22522), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1458.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i803_3_lut (.I0(n1170), .I1(n6579), .I2(n1193), .I3(GND_net), 
            .O(n1293));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i803_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3033_11 (.CI(n37871), .I0(n49961), .I1(n1991), .CO(n37872));
    SB_LUT4 add_3033_10_lut (.I0(n2094), .I1(n49961), .I2(n2093), .I3(n37870), 
            .O(displacement_23__N_91[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_12_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4063));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_91[21]), 
            .I2(n3_adj_3999), .I3(n37166), .O(displacement_23__N_1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3033_10 (.CI(n37870), .I0(n49961), .I1(n2093), .CO(n37871));
    SB_LUT4 add_3033_9_lut (.I0(n2193), .I1(n49961), .I2(n2192), .I3(n37869), 
            .O(displacement_23__N_91[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_9 (.CI(n37869), .I0(n49961), .I1(n2192), .CO(n37870));
    SB_LUT4 add_3033_8_lut (.I0(n2289), .I1(n49961), .I2(n2288), .I3(n37868), 
            .O(displacement_23__N_91[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_8 (.CI(n37868), .I0(n49961), .I1(n2288), .CO(n37869));
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n37166), .I0(displacement_23__N_91[21]), 
            .I1(n3_adj_3999), .CO(n37167));
    SB_LUT4 add_3033_7_lut (.I0(n2382), .I1(n49961), .I2(n2381), .I3(n37867), 
            .O(displacement_23__N_91[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_7 (.CI(n37867), .I0(n49961), .I1(n2381), .CO(n37868));
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_91[20]), 
            .I2(n3_adj_3999), .I3(n37165), .O(displacement_23__N_1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3033_6_lut (.I0(n2472), .I1(n49961), .I2(n2471), .I3(n37866), 
            .O(displacement_23__N_91[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_12_i1763_3_lut_3_lut (.I0(n2642), .I1(n6989), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4062));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3033_6 (.CI(n37866), .I0(n49961), .I1(n2471), .CO(n37867));
    SB_LUT4 add_3033_5_lut (.I0(n2559), .I1(n49961), .I2(n2558), .I3(n37865), 
            .O(displacement_23__N_91[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_12_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n379));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3033_5 (.CI(n37865), .I0(n49961), .I1(n2558), .CO(n37866));
    SB_LUT4 div_12_i1125_3_lut (.I0(n379), .I1(n6753), .I2(n1667), .I3(GND_net), 
            .O(n1765));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3033_4_lut (.I0(n2643), .I1(n49961), .I2(n2642), .I3(n37864), 
            .O(displacement_23__N_91[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3033_4 (.CI(n37864), .I0(n49961), .I1(n2642), .CO(n37865));
    SB_LUT4 div_12_i1198_3_lut (.I0(n1765), .I1(n6794), .I2(n1778), .I3(GND_net), 
            .O(n1873));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3033_3_lut (.I0(n2724), .I1(n49961), .I2(n2723), .I3(n37863), 
            .O(displacement_23__N_91[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n37165), .I0(displacement_23__N_91[20]), 
            .I1(n3_adj_3999), .CO(n37166));
    SB_CARRY add_3033_3 (.CI(n37863), .I0(n49961), .I1(n2723), .CO(n37864));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_91[19]), 
            .I2(n6_adj_3985), .I3(n37164), .O(displacement_23__N_1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3033_2_lut (.I0(n2802), .I1(n49961), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_91[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3033_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n37164), .I0(displacement_23__N_91[19]), 
            .I1(n6_adj_3985), .CO(n37165));
    SB_CARRY add_3033_2 (.CI(VCC_net), .I0(n49961), .I1(n2801), .CO(n37863));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_91[18]), 
            .I2(n7_adj_3984), .I3(n37163), .O(displacement_23__N_1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n37862), 
            .O(n7004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n37163), .I0(displacement_23__N_91[18]), 
            .I1(n7_adj_3984), .CO(n37164));
    SB_LUT4 div_12_i1771_3_lut_3_lut (.I0(n2642), .I1(n6997), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4061));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3032_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n37861), 
            .O(n7005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_24 (.CI(n37861), .I0(n2700), .I1(n79), .CO(n37862));
    SB_LUT4 add_3032_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n37860), 
            .O(n7006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n378));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3032_23 (.CI(n37860), .I0(n2701), .I1(n80), .CO(n37861));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_91[17]), 
            .I2(n8_adj_3983), .I3(n37162), .O(displacement_23__N_1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n37859), 
            .O(n7007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n37162), .I0(displacement_23__N_91[17]), 
            .I1(n8_adj_3983), .CO(n37163));
    SB_CARRY add_3032_22 (.CI(n37859), .I0(n2702), .I1(n81), .CO(n37860));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_91[16]), 
            .I2(n9_adj_3982), .I3(n37161), .O(displacement_23__N_1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1049_3_lut (.I0(n378), .I1(n6739), .I2(n1553), .I3(GND_net), 
            .O(n1653));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n37161), .I0(displacement_23__N_91[16]), 
            .I1(n9_adj_3982), .CO(n37162));
    SB_LUT4 add_3032_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n37858), 
            .O(n7008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_91[15]), 
            .I2(n10_adj_3981), .I3(n37160), .O(displacement_23__N_1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_21 (.CI(n37858), .I0(n2703), .I1(n82), .CO(n37859));
    SB_LUT4 add_3032_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n37857), 
            .O(n7009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_1[23]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n37160), .I0(displacement_23__N_91[15]), 
            .I1(n10_adj_3981), .CO(n37161));
    SB_CARRY add_3032_20 (.CI(n37857), .I0(n2704), .I1(n83), .CO(n37858));
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_91[14]), 
            .I2(n11_adj_3980), .I3(n37159), .O(displacement_23__N_1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n37856), 
            .O(n7010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_19 (.CI(n37856), .I0(n2705), .I1(n84), .CO(n37857));
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n37159), .I0(displacement_23__N_91[14]), 
            .I1(n11_adj_3980), .CO(n37160));
    SB_LUT4 add_3032_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n37855), 
            .O(n7011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_18 (.CI(n37855), .I0(n2706), .I1(n85), .CO(n37856));
    SB_LUT4 add_3032_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n37854), 
            .O(n7012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_17 (.CI(n37854), .I0(n2707), .I1(n86), .CO(n37855));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_91[13]), 
            .I2(n12_adj_3979), .I3(n37158), .O(displacement_23__N_1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n37853), 
            .O(n7013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n37158), .I0(displacement_23__N_91[13]), 
            .I1(n12_adj_3979), .CO(n37159));
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_91[12]), 
            .I2(n13_adj_3978), .I3(n37157), .O(displacement_23__N_1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n37157), .I0(displacement_23__N_91[12]), 
            .I1(n13_adj_3978), .CO(n37158));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_91[11]), 
            .I2(n14_adj_3977), .I3(n37156), .O(displacement_23__N_1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n37156), .I0(displacement_23__N_91[11]), 
            .I1(n14_adj_3977), .CO(n37157));
    SB_CARRY add_3032_16 (.CI(n37853), .I0(n2708), .I1(n87), .CO(n37854));
    SB_LUT4 add_3032_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n37852), 
            .O(n7014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_15 (.CI(n37852), .I0(n2709), .I1(n88), .CO(n37853));
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_91[10]), 
            .I2(n15_adj_3976), .I3(n37155), .O(displacement_23__N_1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n37155), .I0(displacement_23__N_91[10]), 
            .I1(n15_adj_3976), .CO(n37156));
    SB_LUT4 div_12_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4060));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1124_3_lut (.I0(n1653), .I1(n6752), .I2(n1667), .I3(GND_net), 
            .O(n1764));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n22459), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_3992));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_12_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4059));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1197_3_lut (.I0(n1764), .I1(n6793), .I2(n1778), .I3(GND_net), 
            .O(n1872));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1459 (.I0(control_mode[0]), .I1(n22459), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_3965));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i1_2_lut_3_lut_adj_1459.LUT_INIT = 16'hefef;
    SB_LUT4 div_12_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4058));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_91[9]), 
            .I2(n16_adj_3975), .I3(n37154), .O(displacement_23__N_1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n37154), .I0(displacement_23__N_91[9]), 
            .I1(n16_adj_3975), .CO(n37155));
    SB_LUT4 div_12_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4057));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3032_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n37851), 
            .O(n7015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_91[8]), 
            .I2(n17_adj_3974), .I3(n37153), .O(displacement_23__N_1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n37153), .I0(displacement_23__N_91[8]), 
            .I1(n17_adj_3974), .CO(n37154));
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_91[7]), 
            .I2(n18_adj_3973), .I3(n37152), .O(displacement_23__N_1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n37152), .I0(displacement_23__N_91[7]), 
            .I1(n18_adj_3973), .CO(n37153));
    SB_CARRY add_3032_14 (.CI(n37851), .I0(n2710), .I1(n89), .CO(n37852));
    SB_LUT4 div_12_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n377));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4056));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i971_3_lut (.I0(n377), .I1(n6698), .I2(n1436), .I3(GND_net), 
            .O(n1538));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3032_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n37850), 
            .O(n7016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_91[6]), 
            .I2(n19_adj_3972), .I3(n37151), .O(displacement_23__N_1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n37151), .I0(displacement_23__N_91[6]), 
            .I1(n19_adj_3972), .CO(n37152));
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_91[5]), 
            .I2(n20_adj_3971), .I3(n37150), .O(displacement_23__N_1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_1[22]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_LUT4 div_12_i1048_3_lut (.I0(n1538), .I1(n6738), .I2(n1553), .I3(GND_net), 
            .O(n1652));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n37150), .I0(displacement_23__N_91[5]), 
            .I1(n20_adj_3971), .CO(n37151));
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_91[4]), 
            .I2(n21_adj_3970), .I3(n37149), .O(displacement_23__N_1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_13 (.CI(n37850), .I0(n2711), .I1(n90), .CO(n37851));
    SB_LUT4 add_3032_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n37849), 
            .O(n7017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_12 (.CI(n37849), .I0(n2712), .I1(n91), .CO(n37850));
    SB_LUT4 add_3032_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n37848), 
            .O(n7018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_11 (.CI(n37848), .I0(n2713), .I1(n92), .CO(n37849));
    SB_LUT4 add_3032_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n37847), 
            .O(n7019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n37149), .I0(displacement_23__N_91[4]), 
            .I1(n21_adj_3970), .CO(n37150));
    SB_CARRY add_3032_10 (.CI(n37847), .I0(n2714), .I1(n93), .CO(n37848));
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_91[3]), 
            .I2(n22_adj_3969), .I3(n37148), .O(displacement_23__N_1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n37846), 
            .O(n7020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n37148), .I0(displacement_23__N_91[3]), 
            .I1(n22_adj_3969), .CO(n37149));
    SB_CARRY add_3032_9 (.CI(n37846), .I0(n2715), .I1(n94), .CO(n37847));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_91[2]), 
            .I2(n23_adj_3968), .I3(n37147), .O(displacement_23__N_1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3032_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n37845), 
            .O(n7021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_8 (.CI(n37845), .I0(n2716), .I1(n95), .CO(n37846));
    SB_LUT4 add_3032_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n37844), 
            .O(n7022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_7 (.CI(n37844), .I0(n2717), .I1(n96), .CO(n37845));
    SB_LUT4 add_3032_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n37843), 
            .O(n7023)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n37147), .I0(displacement_23__N_91[2]), 
            .I1(n23_adj_3968), .CO(n37148));
    SB_CARRY add_3032_6 (.CI(n37843), .I0(n2718), .I1(n97), .CO(n37844));
    SB_LUT4 add_3032_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n37842), 
            .O(n7024)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_91[1]), 
            .I2(n24_adj_3967), .I3(n37146), .O(displacement_23__N_1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_5 (.CI(n37842), .I0(n2719), .I1(n98), .CO(n37843));
    SB_LUT4 add_3032_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n37841), 
            .O(n7025)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3032_4 (.CI(n37841), .I0(n2720), .I1(n99), .CO(n37842));
    SB_LUT4 add_3032_3_lut (.I0(GND_net), .I1(n390), .I2(n558), .I3(n37840), 
            .O(n7026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3032_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n37146), .I0(displacement_23__N_91[1]), 
            .I1(n24_adj_3967), .CO(n37147));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_91[0]), 
            .I2(n25_adj_3966), .I3(VCC_net), .O(displacement_23__N_1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_91[0]), 
            .I1(n25_adj_3966), .CO(n37146));
    SB_CARRY add_3032_3 (.CI(n37840), .I0(n390), .I1(n558), .CO(n37841));
    SB_LUT4 div_12_i1123_3_lut (.I0(n1652), .I1(n6751), .I2(n1667), .I3(GND_net), 
            .O(n1763));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1123_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_1[21]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_1[20]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_1[19]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_1[18]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_1[17]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_1[16]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_1[15]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_1[14]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_1[13]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_1[12]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_1[11]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_1[10]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_1[9]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_1[8]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_1[7]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_1[6]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_1[5]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_1[4]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_1[3]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_1[2]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_1[1]));   // verilog/TinyFPGA_B.v(161[10] 163[6])
    SB_LUT4 div_12_LessThan_1137_i38_3_lut (.I0(n30_adj_4133), .I1(n91), 
            .I2(n41_adj_4140), .I3(GND_net), .O(n38_adj_4138));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33296_3_lut (.I0(n48962), .I1(n93), .I2(n43_adj_4110), .I3(GND_net), 
            .O(n48798));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33296_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1137_i26_4_lut (.I0(n380), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33449_3_lut (.I0(n26), .I1(n95), .I2(n33_adj_4135), .I3(GND_net), 
            .O(n48951));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33449_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33450_3_lut (.I0(n48951), .I1(n94), .I2(n35_adj_4136), .I3(GND_net), 
            .O(n48952));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33450_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31927_4_lut (.I0(n39_adj_4139), .I1(n37_adj_4137), .I2(n35_adj_4136), 
            .I3(n47434), .O(n47427));
    defparam i31927_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3032_2 (.CI(VCC_net), .I0(n391), .I1(VCC_net), .CO(n37840));
    SB_LUT4 div_12_i1196_3_lut (.I0(n1763), .I1(n6792), .I2(n1778), .I3(GND_net), 
            .O(n1871));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33457_4_lut (.I0(n48798), .I1(n48580), .I2(n43_adj_4110), 
            .I3(n48176), .O(n48959));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33457_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33458_3_lut (.I0(n48959), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n48960));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33458_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1460 (.I0(n48960), .I1(n22525), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1460.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i884_3_lut (.I0(n1293), .I1(n6650), .I2(n1316), .I3(GND_net), 
            .O(n1413));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31984_4_lut (.I0(n37_adj_4114), .I1(n35), .I2(n33), .I3(n31), 
            .O(n47484));
    defparam i31984_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3031_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n37839), 
            .O(n6980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4055));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n376));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3031_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n37838), 
            .O(n6981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i891_3_lut (.I0(n376), .I1(n6657), .I2(n1316), .I3(GND_net), 
            .O(n1420));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i891_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_22 (.CI(n37838), .I0(n2619), .I1(n80), .CO(n37839));
    SB_LUT4 div_12_i970_3_lut (.I0(n1420), .I1(n6697), .I2(n1436), .I3(GND_net), 
            .O(n1537));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4054));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3031_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n37837), 
            .O(n6982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1047_3_lut (.I0(n1537), .I1(n6737), .I2(n1553), .I3(GND_net), 
            .O(n1651));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_21 (.CI(n37837), .I0(n2620), .I1(n81), .CO(n37838));
    SB_LUT4 div_12_i1122_3_lut (.I0(n1651), .I1(n6750), .I2(n1667), .I3(GND_net), 
            .O(n1762));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4053));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1195_3_lut (.I0(n1762), .I1(n6791), .I2(n1778), .I3(GND_net), 
            .O(n1870));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n375));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3031_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n37836), 
            .O(n6983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4052));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i809_3_lut (.I0(n375), .I1(n6585), .I2(n1193), .I3(GND_net), 
            .O(n1299));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i809_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i890_3_lut (.I0(n1299), .I1(n6656), .I2(n1316), .I3(GND_net), 
            .O(n1419));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i890_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_20 (.CI(n37836), .I0(n2621), .I1(n82), .CO(n37837));
    SB_LUT4 div_12_i969_3_lut (.I0(n1419), .I1(n6696), .I2(n1436), .I3(GND_net), 
            .O(n1536));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1046_3_lut (.I0(n1536), .I1(n6736), .I2(n1553), .I3(GND_net), 
            .O(n1650));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n37835), 
            .O(n6984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_19 (.CI(n37835), .I0(n2622), .I1(n83), .CO(n37836));
    SB_LUT4 div_12_i1121_3_lut (.I0(n1650), .I1(n6749), .I2(n1667), .I3(GND_net), 
            .O(n1761));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n37834), 
            .O(n6985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_18 (.CI(n37834), .I0(n2623), .I1(n84), .CO(n37835));
    SB_LUT4 div_12_i1194_3_lut (.I0(n1761), .I1(n6790), .I2(n1778), .I3(GND_net), 
            .O(n1869));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4051));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3031_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n37833), 
            .O(n6986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_17 (.CI(n37833), .I0(n2624), .I1(n85), .CO(n37834));
    SB_LUT4 add_3031_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n37832), 
            .O(n6987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_16 (.CI(n37832), .I0(n2625), .I1(n86), .CO(n37833));
    SB_LUT4 add_3031_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n37831), 
            .O(n6988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_15 (.CI(n37831), .I0(n2626), .I1(n87), .CO(n37832));
    SB_LUT4 add_3031_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n37830), 
            .O(n6989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10630_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n43231), 
            .I3(GND_net), .O(n24045));   // verilog/coms.v(125[12] 284[6])
    defparam i10630_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_14 (.CI(n37830), .I0(n2627), .I1(n88), .CO(n37831));
    SB_LUT4 i10631_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n43231), 
            .I3(GND_net), .O(n24046));   // verilog/coms.v(125[12] 284[6])
    defparam i10631_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n37829), 
            .O(n6990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n373));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3031_13 (.CI(n37829), .I0(n2628), .I1(n89), .CO(n37830));
    SB_LUT4 add_3031_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n37828), 
            .O(n6991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_12 (.CI(n37828), .I0(n2629), .I1(n90), .CO(n37829));
    SB_LUT4 add_3031_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n37827), 
            .O(n6992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_11_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_6_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b011001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_24_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b000001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i33648_4_lut (.I0(n38_adj_4138), .I1(n28_adj_4131), .I2(n41_adj_4140), 
            .I3(n47425), .O(n49150));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33648_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_12_i639_3_lut (.I0(n373), .I1(n5830), .I2(n938), .I3(GND_net), 
            .O(n1048));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i639_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10632_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n43231), 
            .I3(GND_net), .O(n24047));   // verilog/coms.v(125[12] 284[6])
    defparam i10632_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_985_i42_3_lut (.I0(n34_adj_4113), .I1(n91), 
            .I2(n45_adj_4119), .I3(GND_net), .O(n42_adj_4117));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i724_3_lut (.I0(n1048), .I1(n6222), .I2(n1067), .I3(GND_net), 
            .O(n1174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i724_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_11 (.CI(n37827), .I0(n2630), .I1(n91), .CO(n37828));
    SB_LUT4 i10633_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n43231), 
            .I3(GND_net), .O(n24048));   // verilog/coms.v(125[12] 284[6])
    defparam i10633_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4050));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i807_3_lut (.I0(n1174), .I1(n6583), .I2(n1193), .I3(GND_net), 
            .O(n1297));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i807_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10634_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n43231), 
            .I3(GND_net), .O(n24049));   // verilog/coms.v(125[12] 284[6])
    defparam i10634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10635_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n43231), 
            .I3(GND_net), .O(n24050));   // verilog/coms.v(125[12] 284[6])
    defparam i10635_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n37826), 
            .O(n6993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i888_3_lut (.I0(n1297), .I1(n6654), .I2(n1316), .I3(GND_net), 
            .O(n1417));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i967_3_lut (.I0(n1417), .I1(n6694), .I2(n1436), .I3(GND_net), 
            .O(n1534));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i967_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_10 (.CI(n37826), .I0(n2631), .I1(n92), .CO(n37827));
    SB_LUT4 div_12_i1044_3_lut (.I0(n1534), .I1(n6734), .I2(n1553), .I3(GND_net), 
            .O(n1648));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n37825), 
            .O(n6994)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_9 (.CI(n37825), .I0(n2632), .I1(n93), .CO(n37826));
    SB_LUT4 div_12_i1119_3_lut (.I0(n1648), .I1(n6747), .I2(n1667), .I3(GND_net), 
            .O(n1759));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10636_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n43231), 
            .I3(GND_net), .O(n24051));   // verilog/coms.v(125[12] 284[6])
    defparam i10636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n37824), 
            .O(n6995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1192_3_lut (.I0(n1759), .I1(n6788), .I2(n1778), .I3(GND_net), 
            .O(n1867));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1192_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_8 (.CI(n37824), .I0(n2633), .I1(n94), .CO(n37825));
    SB_LUT4 add_3031_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n37823), 
            .O(n6996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32299_3_lut (.I0(n372), .I1(n558), .I2(n806), .I3(GND_net), 
            .O(n918));
    defparam i32299_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_12_i638_3_lut (.I0(n918), .I1(n5829), .I2(n938), .I3(GND_net), 
            .O(n1047));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i638_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10637_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n43231), 
            .I3(GND_net), .O(n24052));   // verilog/coms.v(125[12] 284[6])
    defparam i10637_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_7 (.CI(n37823), .I0(n2634), .I1(n95), .CO(n37824));
    SB_LUT4 div_12_i723_3_lut (.I0(n1047), .I1(n6221), .I2(n1067), .I3(GND_net), 
            .O(n1173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n37822), 
            .O(n6997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i806_3_lut (.I0(n1173), .I1(n6582), .I2(n1193), .I3(GND_net), 
            .O(n1296));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i806_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i887_3_lut (.I0(n1296), .I1(n6653), .I2(n1316), .I3(GND_net), 
            .O(n1416));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i887_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_6 (.CI(n37822), .I0(n2635), .I1(n96), .CO(n37823));
    SB_LUT4 add_3031_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n37821), 
            .O(n6998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_5 (.CI(n37821), .I0(n2636), .I1(n97), .CO(n37822));
    SB_LUT4 add_3031_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n37820), 
            .O(n6999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i966_3_lut (.I0(n1416), .I1(n6693), .I2(n1436), .I3(GND_net), 
            .O(n1533));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i966_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1043_3_lut (.I0(n1533), .I1(n6733), .I2(n1553), .I3(GND_net), 
            .O(n1647));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3031_4 (.CI(n37820), .I0(n2637), .I1(n98), .CO(n37821));
    SB_LUT4 div_12_i1118_3_lut (.I0(n1647), .I1(n6746), .I2(n1667), .I3(GND_net), 
            .O(n1758));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1191_3_lut (.I0(n1758), .I1(n6787), .I2(n1778), .I3(GND_net), 
            .O(n1866));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3031_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n37819), 
            .O(n7000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_985_i30_4_lut (.I0(n378), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30_adj_4111));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY add_3031_3 (.CI(n37819), .I0(n2638), .I1(n99), .CO(n37820));
    SB_LUT4 add_3031_2_lut (.I0(GND_net), .I1(n389), .I2(n558), .I3(VCC_net), 
            .O(n7001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3031_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3031_2 (.CI(VCC_net), .I0(n389), .I1(n558), .CO(n37819));
    SB_LUT4 add_3030_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n37818), 
            .O(n6957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4049));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3030_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n37817), 
            .O(n6958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i550_4_lut (.I0(n785), .I1(n2_adj_4094), .I2(n806), 
            .I3(n99), .O(n917));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i550_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_i637_3_lut (.I0(n917), .I1(n5828), .I2(n938), .I3(GND_net), 
            .O(n1046));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i637_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i722_3_lut (.I0(n1046), .I1(n6220), .I2(n1067), .I3(GND_net), 
            .O(n1172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i722_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3030_21 (.CI(n37817), .I0(n2535), .I1(n81), .CO(n37818));
    SB_LUT4 add_3030_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n37816), 
            .O(n6959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_20 (.CI(n37816), .I0(n2536), .I1(n82), .CO(n37817));
    SB_LUT4 add_3030_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n37815), 
            .O(n6960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i805_3_lut (.I0(n1172), .I1(n6581), .I2(n1193), .I3(GND_net), 
            .O(n1295));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i805_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i886_3_lut (.I0(n1295), .I1(n6652), .I2(n1316), .I3(GND_net), 
            .O(n1415));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i965_3_lut (.I0(n1415), .I1(n6692), .I2(n1436), .I3(GND_net), 
            .O(n1532));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i965_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3030_19 (.CI(n37815), .I0(n2537), .I1(n83), .CO(n37816));
    SB_LUT4 add_3030_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n37814), 
            .O(n6961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1042_3_lut (.I0(n1532), .I1(n6732), .I2(n1553), .I3(GND_net), 
            .O(n1646));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1117_3_lut (.I0(n1646), .I1(n6745), .I2(n1667), .I3(GND_net), 
            .O(n1757));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_3030_18 (.CI(n37814), .I0(n2538), .I1(n84), .CO(n37815));
    SB_LUT4 add_3030_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n37813), 
            .O(n6962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_i1190_3_lut (.I0(n1757), .I1(n6786), .I2(n1778), .I3(GND_net), 
            .O(n1865));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1190_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3030_17 (.CI(n37813), .I0(n2539), .I1(n85), .CO(n37814));
    SB_LUT4 add_3030_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n37812), 
            .O(n6963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_16 (.CI(n37812), .I0(n2540), .I1(n86), .CO(n37813));
    SB_LUT4 add_3030_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n37811), 
            .O(n6964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_15 (.CI(n37811), .I0(n2541), .I1(n87), .CO(n37812));
    SB_LUT4 add_3030_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n37810), 
            .O(n6965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_14 (.CI(n37810), .I0(n2542), .I1(n88), .CO(n37811));
    SB_LUT4 add_3030_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n37809), 
            .O(n6966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_13 (.CI(n37809), .I0(n2543), .I1(n89), .CO(n37810));
    SB_LUT4 add_3030_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n37808), 
            .O(n6967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_12 (.CI(n37808), .I0(n2544), .I1(n90), .CO(n37809));
    SB_LUT4 add_3030_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n37807), 
            .O(n6968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_11 (.CI(n37807), .I0(n2545), .I1(n91), .CO(n37808));
    SB_LUT4 add_3030_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n37806), 
            .O(n6969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_10_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_19_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b000001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_3030_10 (.CI(n37806), .I0(n2546), .I1(n92), .CO(n37807));
    SB_LUT4 add_3030_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n37805), 
            .O(n6970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_9 (.CI(n37805), .I0(n2547), .I1(n93), .CO(n37806));
    SB_LUT4 add_3030_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n37804), 
            .O(n6971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_8 (.CI(n37804), .I0(n2548), .I1(n94), .CO(n37805));
    SB_LUT4 add_3030_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n37803), 
            .O(n6972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_7 (.CI(n37803), .I0(n2549), .I1(n95), .CO(n37804));
    SB_LUT4 add_3030_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n37802), 
            .O(n6973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_6 (.CI(n37802), .I0(n2550), .I1(n96), .CO(n37803));
    SB_LUT4 add_3030_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n37801), 
            .O(n6974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_5 (.CI(n37801), .I0(n2551), .I1(n97), .CO(n37802));
    SB_LUT4 add_3030_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n37800), 
            .O(n6975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_4 (.CI(n37800), .I0(n2552), .I1(n98), .CO(n37801));
    SB_LUT4 add_3030_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n37799), 
            .O(n6976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_3 (.CI(n37799), .I0(n2553), .I1(n99), .CO(n37800));
    SB_LUT4 add_3030_2_lut (.I0(GND_net), .I1(n388), .I2(n558), .I3(VCC_net), 
            .O(n6977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3030_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3030_2 (.CI(VCC_net), .I0(n388), .I1(n558), .CO(n37799));
    SB_LUT4 add_3029_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n37798), 
            .O(n6935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3029_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n37797), 
            .O(n6936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_20 (.CI(n37797), .I0(n2448), .I1(n82), .CO(n37798));
    SB_LUT4 add_3029_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n37796), 
            .O(n6937)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_19 (.CI(n37796), .I0(n2449), .I1(n83), .CO(n37797));
    SB_LUT4 add_3029_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n37795), 
            .O(n6938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_18 (.CI(n37795), .I0(n2450), .I1(n84), .CO(n37796));
    SB_LUT4 add_3029_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n37794), 
            .O(n6939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_17 (.CI(n37794), .I0(n2451), .I1(n85), .CO(n37795));
    SB_LUT4 add_3029_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n37793), 
            .O(n6940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_16 (.CI(n37793), .I0(n2452), .I1(n86), .CO(n37794));
    SB_LUT4 add_3029_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n37792), 
            .O(n6941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_15 (.CI(n37792), .I0(n2453), .I1(n87), .CO(n37793));
    SB_LUT4 add_3029_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n37791), 
            .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_14 (.CI(n37791), .I0(n2454), .I1(n88), .CO(n37792));
    SB_LUT4 add_3029_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n37790), 
            .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_13 (.CI(n37790), .I0(n2455), .I1(n89), .CO(n37791));
    SB_LUT4 add_3029_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n37789), 
            .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_12 (.CI(n37789), .I0(n2456), .I1(n90), .CO(n37790));
    SB_LUT4 add_3029_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n37788), 
            .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_11 (.CI(n37788), .I0(n2457), .I1(n91), .CO(n37789));
    SB_LUT4 add_3029_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n37787), 
            .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10828_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24243));   // verilog/coms.v(125[12] 284[6])
    defparam i10828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4048));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3029_10 (.CI(n37787), .I0(n2458), .I1(n92), .CO(n37788));
    SB_LUT4 add_3029_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n37786), 
            .O(n6947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_9 (.CI(n37786), .I0(n2459), .I1(n93), .CO(n37787));
    SB_LUT4 add_3029_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n37785), 
            .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_2_lut (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_515));   // verilog/coms.v(93[12:25])
    defparam i7_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3029_8 (.CI(n37785), .I0(n2460), .I1(n94), .CO(n37786));
    SB_LUT4 add_3029_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n37784), 
            .O(n6949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_7 (.CI(n37784), .I0(n2461), .I1(n95), .CO(n37785));
    SB_LUT4 add_3029_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n37783), 
            .O(n6950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33306_3_lut (.I0(n48952), .I1(n93), .I2(n37_adj_4137), .I3(GND_net), 
            .O(n48808));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33306_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10646_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n43229), 
            .I3(GND_net), .O(n24061));   // verilog/coms.v(125[12] 284[6])
    defparam i10646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10647_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n43229), 
            .I3(GND_net), .O(n24062));   // verilog/coms.v(125[12] 284[6])
    defparam i10647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33455_3_lut (.I0(n30_adj_4111), .I1(n95), .I2(n37_adj_4114), 
            .I3(GND_net), .O(n48957));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33455_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10648_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n43229), 
            .I3(GND_net), .O(n24063));   // verilog/coms.v(125[12] 284[6])
    defparam i10648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4047));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10649_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n43229), 
            .I3(GND_net), .O(n24064));   // verilog/coms.v(125[12] 284[6])
    defparam i10649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4046));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3029_6 (.CI(n37783), .I0(n2462), .I1(n96), .CO(n37784));
    SB_LUT4 add_3029_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n37782), 
            .O(n6951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10650_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n43229), 
            .I3(GND_net), .O(n24065));   // verilog/coms.v(125[12] 284[6])
    defparam i10650_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3029_5 (.CI(n37782), .I0(n2463), .I1(n97), .CO(n37783));
    SB_LUT4 add_3029_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n37781), 
            .O(n6952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_4 (.CI(n37781), .I0(n2464), .I1(n98), .CO(n37782));
    SB_LUT4 add_3029_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n37780), 
            .O(n6953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_3 (.CI(n37780), .I0(n2465), .I1(n99), .CO(n37781));
    SB_LUT4 add_3029_2_lut (.I0(GND_net), .I1(n387_adj_4000), .I2(n558), 
            .I3(VCC_net), .O(n6954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3029_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3029_2 (.CI(VCC_net), .I0(n387_adj_4000), .I1(n558), 
            .CO(n37780));
    SB_LUT4 add_3028_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n37779), 
            .O(n6914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3028_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n37778), 
            .O(n6915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_19 (.CI(n37778), .I0(n2358), .I1(n83), .CO(n37779));
    SB_LUT4 add_3028_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n37777), 
            .O(n6916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_18 (.CI(n37777), .I0(n2359), .I1(n84), .CO(n37778));
    SB_LUT4 add_3028_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n37776), 
            .O(n6917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_17 (.CI(n37776), .I0(n2360), .I1(n85), .CO(n37777));
    SB_LUT4 add_3028_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n37775), 
            .O(n6918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_16 (.CI(n37775), .I0(n2361), .I1(n86), .CO(n37776));
    SB_LUT4 i10651_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n43229), 
            .I3(GND_net), .O(n24066));   // verilog/coms.v(125[12] 284[6])
    defparam i10651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3028_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n37774), 
            .O(n6919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10652_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n43229), 
            .I3(GND_net), .O(n24067));   // verilog/coms.v(125[12] 284[6])
    defparam i10652_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_3028_15 (.CI(n37774), .I0(n2362), .I1(n87), .CO(n37775));
    SB_LUT4 add_3028_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n37773), 
            .O(n6920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_14 (.CI(n37773), .I0(n2363), .I1(n88), .CO(n37774));
    SB_LUT4 add_3028_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n37772), 
            .O(n6921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_13 (.CI(n37772), .I0(n2364), .I1(n89), .CO(n37773));
    SB_LUT4 add_3028_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n37771), 
            .O(n6922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_12 (.CI(n37771), .I0(n2365), .I1(n90), .CO(n37772));
    SB_LUT4 add_3028_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n37770), 
            .O(n6923)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_11 (.CI(n37770), .I0(n2366), .I1(n91), .CO(n37771));
    SB_LUT4 add_3028_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n37769), 
            .O(n6924)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_10 (.CI(n37769), .I0(n2367), .I1(n92), .CO(n37770));
    SB_LUT4 add_3028_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n37768), 
            .O(n6925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_9 (.CI(n37768), .I0(n2368), .I1(n93), .CO(n37769));
    SB_LUT4 add_3028_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n37767), 
            .O(n6926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_8 (.CI(n37767), .I0(n2369), .I1(n94), .CO(n37768));
    SB_LUT4 i10653_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n43229), 
            .I3(GND_net), .O(n24068));   // verilog/coms.v(125[12] 284[6])
    defparam i10653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3028_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n37766), 
            .O(n6927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_7 (.CI(n37766), .I0(n2370), .I1(n95), .CO(n37767));
    SB_LUT4 add_3028_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n37765), 
            .O(n6928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_6 (.CI(n37765), .I0(n2371), .I1(n96), .CO(n37766));
    SB_LUT4 add_3028_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n37764), 
            .O(n6929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\data_in_frame[15] [6]), .I1(n43441), .I2(\data_in_frame[13] [5]), 
            .I3(n22833), .O(n43709));   // verilog/coms.v(93[12:25])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3028_5 (.CI(n37764), .I0(n2372), .I1(n97), .CO(n37765));
    SB_LUT4 add_3028_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n37763), 
            .O(n6930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_4 (.CI(n37763), .I0(n2373), .I1(n98), .CO(n37764));
    SB_LUT4 div_12_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4093));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3028_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n37762), 
            .O(n6931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33456_3_lut (.I0(n48957), .I1(n94), .I2(n39_adj_4115), .I3(GND_net), 
            .O(n48958));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33456_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3028_3 (.CI(n37762), .I0(n2374), .I1(n99), .CO(n37763));
    SB_LUT4 add_3028_2_lut (.I0(GND_net), .I1(n386), .I2(n558), .I3(VCC_net), 
            .O(n6932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3028_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3028_2 (.CI(VCC_net), .I0(n386), .I1(n558), .CO(n37762));
    SB_LUT4 add_3027_19_lut (.I0(GND_net), .I1(n2264_adj_4009), .I2(n83), 
            .I3(n37761), .O(n6894)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4092));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4091));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3027_18_lut (.I0(GND_net), .I1(n2265_adj_4010), .I2(n84), 
            .I3(n37760), .O(n6895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_18 (.CI(n37760), .I0(n2265_adj_4010), .I1(n84), 
            .CO(n37761));
    SB_LUT4 div_12_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4090));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4089));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4088));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33745_4_lut (.I0(n48808), .I1(n49150), .I2(n41_adj_4140), 
            .I3(n47427), .O(n49247));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33745_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33746_3_lut (.I0(n49247), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n49248));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33746_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33718_3_lut (.I0(n49248), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n49220));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33718_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1461 (.I0(n49220), .I1(n22534), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1461.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1115_3_lut (.I0(n1644), .I1(n6743), .I2(n1667), .I3(GND_net), 
            .O(n1755));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3027_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n37759), 
            .O(n6896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4087));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3027_17 (.CI(n37759), .I0(n2266), .I1(n85), .CO(n37760));
    SB_LUT4 div_12_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1188_3_lut (.I0(n1755), .I1(n6784), .I2(n1778), .I3(GND_net), 
            .O(n1863));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1210_i45_2_lut (.I0(n1863), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4158));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31978_4_lut (.I0(n43_adj_4118), .I1(n41_adj_4116), .I2(n39_adj_4115), 
            .I3(n47484), .O(n47478));
    defparam i31978_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4151));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3027_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n37758), 
            .O(n6897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4142));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31907_4_lut (.I0(n31_adj_4148), .I1(n29_adj_4146), .I2(n27_adj_4144), 
            .I3(n25_adj_4142), .O(n47407));
    defparam i31907_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31892_4_lut (.I0(n37_adj_4153), .I1(n35_adj_4151), .I2(n33_adj_4150), 
            .I3(n47407), .O(n47392));
    defparam i31892_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33080_4_lut (.I0(n42_adj_4117), .I1(n32_adj_4112), .I2(n45_adj_4119), 
            .I3(n47471), .O(n48582));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33080_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33300_3_lut (.I0(n48958), .I1(n93), .I2(n41_adj_4116), .I3(GND_net), 
            .O(n48802));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33300_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1210_i24_4_lut (.I0(n381), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4141));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY add_3027_16 (.CI(n37758), .I0(n2267), .I1(n86), .CO(n37759));
    SB_LUT4 div_12_LessThan_1210_i32_3_lut (.I0(n30_adj_4147), .I1(n93), 
            .I2(n35_adj_4151), .I3(GND_net), .O(n32_adj_4149));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33517_4_lut (.I0(n48802), .I1(n48582), .I2(n45_adj_4119), 
            .I3(n47478), .O(n49019));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33517_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_3027_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n37757), 
            .O(n6898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_12_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4086));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1462 (.I0(n49019), .I1(n22528), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1462.LUT_INIT = 16'hceef;
    SB_CARRY add_3027_15 (.CI(n37757), .I0(n2268), .I1(n87), .CO(n37758));
    SB_LUT4 div_12_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4085));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4084));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1210_i36_3_lut (.I0(n28_adj_4145), .I1(n91), 
            .I2(n39_adj_4154), .I3(GND_net), .O(n36_adj_4152));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i963_3_lut (.I0(n1413), .I1(n6690), .I2(n1436), .I3(GND_net), 
            .O(n1530));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i963_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_3027_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n37756), 
            .O(n6899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_14 (.CI(n37756), .I0(n2269), .I1(n88), .CO(n37757));
    SB_LUT4 add_3027_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n37755), 
            .O(n6900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_13 (.CI(n37755), .I0(n2270), .I1(n89), .CO(n37756));
    SB_LUT4 add_3027_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n37754), 
            .O(n6901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_12 (.CI(n37754), .I0(n2271), .I1(n90), .CO(n37755));
    SB_LUT4 add_3027_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n37753), 
            .O(n6902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_11 (.CI(n37753), .I0(n2272), .I1(n91), .CO(n37754));
    SB_LUT4 add_3027_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n37752), 
            .O(n6903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_10 (.CI(n37752), .I0(n2273), .I1(n92), .CO(n37753));
    SB_LUT4 add_3027_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n37751), 
            .O(n6904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_9 (.CI(n37751), .I0(n2274), .I1(n93), .CO(n37752));
    SB_LUT4 add_3027_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n37750), 
            .O(n6905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33650_4_lut (.I0(n36_adj_4152), .I1(n26_adj_4143), .I2(n39_adj_4154), 
            .I3(n47386), .O(n49152));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33650_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3027_8 (.CI(n37750), .I0(n2275), .I1(n94), .CO(n37751));
    SB_LUT4 add_3027_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n37749), 
            .O(n6906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[18] [2]), .I1(n43709), .I2(\data_in_frame[14] [0]), 
            .I3(\data_in_frame[16] [1]), .O(n10_adj_4035));   // verilog/coms.v(93[12:25])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    GND i1 (.Y(GND_net));
    SB_CARRY add_3027_7 (.CI(n37749), .I0(n2276), .I1(n95), .CO(n37750));
    SB_LUT4 div_12_i1341_3_lut_3_lut (.I0(n1991), .I1(n6854), .I2(n382), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3027_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n37748), 
            .O(n6907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_6 (.CI(n37748), .I0(n2277), .I1(n96), .CO(n37749));
    SB_LUT4 add_3027_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n37747), 
            .O(n6908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_5 (.CI(n37747), .I0(n2278), .I1(n97), .CO(n37748));
    SB_LUT4 add_3027_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n37746), 
            .O(n6909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_4 (.CI(n37746), .I0(n2279), .I1(n98), .CO(n37747));
    SB_LUT4 add_3027_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n37745), 
            .O(n6910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_3 (.CI(n37745), .I0(n2280), .I1(n99), .CO(n37746));
    SB_LUT4 add_3027_2_lut (.I0(GND_net), .I1(n385), .I2(n558), .I3(VCC_net), 
            .O(n6911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3027_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3027_2 (.CI(VCC_net), .I0(n385), .I1(n558), .CO(n37745));
    SB_LUT4 add_3026_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n37744), 
            .O(n6875)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3026_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n37743), 
            .O(n6876)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_17 (.CI(n37743), .I0(n2169), .I1(n85), .CO(n37744));
    SB_LUT4 add_3026_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n37742), 
            .O(n6877)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_16 (.CI(n37742), .I0(n2170), .I1(n86), .CO(n37743));
    SB_LUT4 add_3026_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n37741), 
            .O(n6878)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_15 (.CI(n37741), .I0(n2171), .I1(n87), .CO(n37742));
    SB_LUT4 add_3026_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n37740), 
            .O(n6879)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_14 (.CI(n37740), .I0(n2172), .I1(n88), .CO(n37741));
    SB_LUT4 add_3026_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n37739), 
            .O(n6880)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_13 (.CI(n37739), .I0(n2173), .I1(n89), .CO(n37740));
    SB_LUT4 add_3026_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n37738), 
            .O(n6881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_12 (.CI(n37738), .I0(n2174), .I1(n90), .CO(n37739));
    SB_LUT4 add_3026_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n37737), 
            .O(n6882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_11 (.CI(n37737), .I0(n2175), .I1(n91), .CO(n37738));
    SB_LUT4 add_3026_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n37736), 
            .O(n6883)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_10 (.CI(n37736), .I0(n2176), .I1(n92), .CO(n37737));
    SB_LUT4 add_3026_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n37735), 
            .O(n6884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_9 (.CI(n37735), .I0(n2177), .I1(n93), .CO(n37736));
    SB_LUT4 add_3026_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n37734), 
            .O(n6885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_8 (.CI(n37734), .I0(n2178), .I1(n94), .CO(n37735));
    SB_LUT4 add_3026_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n37733), 
            .O(n6886)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_7 (.CI(n37733), .I0(n2179), .I1(n95), .CO(n37734));
    SB_LUT4 add_3026_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n37732), 
            .O(n6887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_6 (.CI(n37732), .I0(n2180), .I1(n96), .CO(n37733));
    SB_LUT4 add_3026_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n37731), 
            .O(n6888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_5 (.CI(n37731), .I0(n2181), .I1(n97), .CO(n37732));
    SB_LUT4 add_3026_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n37730), 
            .O(n6889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_4 (.CI(n37730), .I0(n2182), .I1(n98), .CO(n37731));
    SB_LUT4 add_3026_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n37729), 
            .O(n6890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_3 (.CI(n37729), .I0(n2183), .I1(n99), .CO(n37730));
    SB_LUT4 add_3026_2_lut (.I0(GND_net), .I1(n384), .I2(n558), .I3(VCC_net), 
            .O(n6891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3026_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3026_2 (.CI(VCC_net), .I0(n384), .I1(n558), .CO(n37729));
    SB_LUT4 add_3025_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n37728), 
            .O(n6857)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3025_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n37727), 
            .O(n6858)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_16 (.CI(n37727), .I0(n2070), .I1(n86), .CO(n37728));
    SB_LUT4 add_3025_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n37726), 
            .O(n6859)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_15 (.CI(n37726), .I0(n2071), .I1(n87), .CO(n37727));
    SB_LUT4 add_3025_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n37725), 
            .O(n6860)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_14 (.CI(n37725), .I0(n2072), .I1(n88), .CO(n37726));
    SB_LUT4 add_3025_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n37724), 
            .O(n6861)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_13 (.CI(n37724), .I0(n2073), .I1(n89), .CO(n37725));
    SB_LUT4 add_3025_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n37723), 
            .O(n6862)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_12 (.CI(n37723), .I0(n2074), .I1(n90), .CO(n37724));
    SB_LUT4 add_3025_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n37722), 
            .O(n6863)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_11 (.CI(n37722), .I0(n2075), .I1(n91), .CO(n37723));
    SB_LUT4 add_3025_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n37721), 
            .O(n6864)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_10 (.CI(n37721), .I0(n2076), .I1(n92), .CO(n37722));
    SB_LUT4 add_3025_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n37720), 
            .O(n6865)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_9 (.CI(n37720), .I0(n2077), .I1(n93), .CO(n37721));
    SB_LUT4 add_3025_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n37719), 
            .O(n6866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_8 (.CI(n37719), .I0(n2078), .I1(n94), .CO(n37720));
    SB_LUT4 add_3025_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n37718), 
            .O(n6867)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_7 (.CI(n37718), .I0(n2079), .I1(n95), .CO(n37719));
    SB_LUT4 add_3025_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n37717), 
            .O(n6868)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_6 (.CI(n37717), .I0(n2080), .I1(n96), .CO(n37718));
    SB_LUT4 add_3025_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n37716), 
            .O(n6869)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_5 (.CI(n37716), .I0(n2081), .I1(n97), .CO(n37717));
    SB_LUT4 add_3025_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n37715), 
            .O(n6870)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_4 (.CI(n37715), .I0(n2082), .I1(n98), .CO(n37716));
    SB_LUT4 add_3025_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n37714), 
            .O(n6871)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_3 (.CI(n37714), .I0(n2083), .I1(n99), .CO(n37715));
    SB_LUT4 add_3025_2_lut (.I0(GND_net), .I1(n383), .I2(n558), .I3(VCC_net), 
            .O(n6872)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3025_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3025_2 (.CI(VCC_net), .I0(n383), .I1(n558), .CO(n37714));
    SB_LUT4 add_3024_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n37713), 
            .O(n6840)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3024_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n37712), 
            .O(n6841)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_15 (.CI(n37712), .I0(n1968), .I1(n87), .CO(n37713));
    SB_LUT4 add_3024_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n37711), 
            .O(n6842)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_14 (.CI(n37711), .I0(n1969), .I1(n88), .CO(n37712));
    SB_LUT4 add_3024_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n37710), 
            .O(n6843)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_13 (.CI(n37710), .I0(n1970), .I1(n89), .CO(n37711));
    SB_LUT4 add_3024_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n37709), 
            .O(n6844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_12 (.CI(n37709), .I0(n1971), .I1(n90), .CO(n37710));
    SB_LUT4 add_3024_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n37708), 
            .O(n6845)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_11 (.CI(n37708), .I0(n1972), .I1(n91), .CO(n37709));
    SB_LUT4 add_3024_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n37707), 
            .O(n6846)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_10 (.CI(n37707), .I0(n1973), .I1(n92), .CO(n37708));
    SB_LUT4 add_3024_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n37706), 
            .O(n6847)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_9 (.CI(n37706), .I0(n1974), .I1(n93), .CO(n37707));
    SB_LUT4 add_3024_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n37705), 
            .O(n6848)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_8 (.CI(n37705), .I0(n1975), .I1(n94), .CO(n37706));
    SB_LUT4 add_3024_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n37704), 
            .O(n6849)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_7 (.CI(n37704), .I0(n1976), .I1(n95), .CO(n37705));
    SB_LUT4 add_3024_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n37703), 
            .O(n6850)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_6 (.CI(n37703), .I0(n1977), .I1(n96), .CO(n37704));
    SB_LUT4 add_3024_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n37702), 
            .O(n6851)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3024_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3024_5 (.CI(n37702), .I0(n1978), .I1(n97), .CO(n37703));
    SB_LUT4 i1_2_lut_adj_1463 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4027));   // verilog/coms.v(93[12:25])
    defparam i1_2_lut_adj_1463.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4083));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4082));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4081));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4080));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4079));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4078));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4077));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4076));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4075));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4074));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4073));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4072));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4071));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4070));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[13] [4]), .I3(GND_net), .O(n43459));
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1464 (.I0(n40155), .I1(n43459), .I2(\data_in_frame[18] [0]), 
            .I3(Kp_23__N_865), .O(n44311));
    defparam i3_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 div_12_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4120));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_3961), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n372));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23112_2_lut (.I0(n372), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4094));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23112_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32302_3_lut (.I0(n371), .I1(n558), .I2(n671), .I3(GND_net), 
            .O(n785));
    defparam i32302_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_12_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_3962), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i23080_2_lut (.I0(n371), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23080_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32314_3_lut (.I0(n370), .I1(n558), .I2(n533), .I3(GND_net), 
            .O(n649));
    defparam i32314_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 div_12_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4103));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4104));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4106));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4108));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i460_4_lut (.I0(n649), .I1(n2), .I2(n671), .I3(n99), 
            .O(n784));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i460_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4109));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4110));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i549_4_lut (.I0(n784), .I1(n4_adj_4045), .I2(n806), 
            .I3(n98), .O(n916));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i549_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4114));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4115));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i636_3_lut (.I0(n916), .I1(n5827), .I2(n938), .I3(GND_net), 
            .O(n1045));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i636_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4118));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i721_3_lut (.I0(n1045), .I1(n6219), .I2(n1067), .I3(GND_net), 
            .O(n1171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4116));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4119));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4124));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i804_3_lut (.I0(n1171), .I1(n6580), .I2(n1193), .I3(GND_net), 
            .O(n1294));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i804_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4122));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4125));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4126));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4129));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4127));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4130));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i885_3_lut (.I0(n1294), .I1(n6651), .I2(n1316), .I3(GND_net), 
            .O(n1414));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4134));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4132));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4135));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4136));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4139));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4137));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i964_3_lut (.I0(n1414), .I1(n6691), .I2(n1436), .I3(GND_net), 
            .O(n1531));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4140));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1465 (.I0(n87), .I1(n22537), .I2(GND_net), .I3(GND_net), 
            .O(n22534));
    defparam i1_2_lut_adj_1465.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_i1041_3_lut (.I0(n1531), .I1(n6731), .I2(n1553), .I3(GND_net), 
            .O(n1645));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4148));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4150));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4146));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4153));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4144));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4154));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i41_2_lut (.I0(n1865), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4155));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1116_3_lut (.I0(n1645), .I1(n6744), .I2(n1667), .I3(GND_net), 
            .O(n1756));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1210_i43_2_lut (.I0(n1864), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4156));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1189_3_lut (.I0(n1756), .I1(n6785), .I2(n1778), .I3(GND_net), 
            .O(n1864));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1189_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10924_3_lut (.I0(encoder1_position[9]), .I1(n2256), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24339));   // quad.v(35[10] 41[6])
    defparam i10924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10925_3_lut (.I0(encoder1_position[10]), .I1(n2255), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24340));   // quad.v(35[10] 41[6])
    defparam i10925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10926_3_lut (.I0(encoder1_position[11]), .I1(n2254), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24341));   // quad.v(35[10] 41[6])
    defparam i10926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10829_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24244));   // verilog/coms.v(125[12] 284[6])
    defparam i10829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(LED_c));   // verilog/TinyFPGA_B.v(64[16:21])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10921_3_lut (.I0(encoder1_position[6]), .I1(n2259), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24336));   // quad.v(35[10] 41[6])
    defparam i10921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10830_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24245));   // verilog/coms.v(125[12] 284[6])
    defparam i10830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32114_3_lut_4_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(pwm_count[2]), .O(n47615));   // verilog/motorControl.v(77[28:44])
    defparam i32114_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_558_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(n873), .I2(n874), 
            .I3(GND_net), .O(n6_adj_4039));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_558_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i10922_3_lut (.I0(encoder1_position[7]), .I1(n2258), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24337));   // quad.v(35[10] 41[6])
    defparam i10922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10923_3_lut (.I0(encoder1_position[8]), .I1(n2257), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24338));   // quad.v(35[10] 41[6])
    defparam i10923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n382));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_555_i15_2_lut (.I0(pwm_count[7]), .I1(pwm[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4034));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_555_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n381));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_555_i9_2_lut (.I0(pwm_count[4]), .I1(pwm[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4031));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_555_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 div_12_i1271_3_lut (.I0(n381), .I1(n6837), .I2(n1886), .I3(GND_net), 
            .O(n1980));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_555_i13_2_lut (.I0(pwm_count[6]), .I1(pwm[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4033));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_555_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_555_i11_2_lut (.I0(pwm_count[5]), .I1(pwm[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4032));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_555_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut (.I0(n21_adj_4004), .I1(n23_adj_4002), .I2(n22_adj_4003), 
            .I3(n24_adj_4001), .O(n30));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n17_adj_4008), .I1(n19_adj_4006), .I2(n18_adj_4007), 
            .I3(n20_adj_4005), .O(n29));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31960_4_lut (.I0(n35_adj_4125), .I1(n33_adj_4124), .I2(n31_adj_4122), 
            .I3(n29_adj_4120), .O(n47460));
    defparam i31960_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10328_3_lut (.I0(\PID_CONTROLLER.err_prev [0]), .I1(\PID_CONTROLLER.err [0]), 
            .I2(n44626), .I3(GND_net), .O(n23743));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28513_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44009));
    defparam i28513_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_555_i4_4_lut (.I0(pwm_count[0]), .I1(pwm[1]), .I2(pwm_count[1]), 
            .I3(pwm[0]), .O(n4_adj_4028));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_555_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\FRAME_MATCHER.state [0]), .I1(n20136), 
            .I2(GND_net), .I3(GND_net), .O(n40_adj_4377));   // verilog/coms.v(125[12] 284[6])
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_1467 (.I0(n44019), .I1(n40_adj_4377), .I2(n45225), 
            .I3(n5_adj_4375), .O(n41_adj_4376));   // verilog/coms.v(125[12] 284[6])
    defparam i1_4_lut_adj_1467.LUT_INIT = 16'hcc4c;
    SB_LUT4 i33217_3_lut (.I0(n4_adj_4028), .I1(pwm[5]), .I2(n11_adj_4032), 
            .I3(GND_net), .O(n48719));   // verilog/motorControl.v(58[19:32])
    defparam i33217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1468 (.I0(n44238), .I1(n41_adj_4376), .I2(n22456), 
            .I3(\FRAME_MATCHER.state [3]), .O(n42561));   // verilog/coms.v(125[12] 284[6])
    defparam i1_4_lut_adj_1468.LUT_INIT = 16'hcdcc;
    SB_LUT4 i10330_3_lut (.I0(encoder0_position[0]), .I1(n2315), .I2(count_enable), 
            .I3(GND_net), .O(n23745));   // quad.v(35[10] 41[6])
    defparam i10330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33218_3_lut (.I0(n48719), .I1(pwm[6]), .I2(n13_adj_4033), 
            .I3(GND_net), .O(n48720));   // verilog/motorControl.v(58[19:32])
    defparam i33218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32771_4_lut (.I0(n13_adj_4033), .I1(n11_adj_4032), .I2(n9_adj_4031), 
            .I3(n47623), .O(n48273));
    defparam i32771_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 LessThan_555_i8_3_lut (.I0(n6_adj_4029), .I1(pwm[4]), .I2(n9_adj_4031), 
            .I3(GND_net), .O(n8_adj_4030));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_555_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10331_3_lut (.I0(encoder1_position[0]), .I1(n2265), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n23746));   // quad.v(35[10] 41[6])
    defparam i10331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32669_3_lut (.I0(n48720), .I1(pwm[7]), .I2(n15_adj_4034), 
            .I3(GND_net), .O(n48171));   // verilog/motorControl.v(58[19:32])
    defparam i32669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10335_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n44902), 
            .I3(GND_net), .O(n23750));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10335_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33275_4_lut (.I0(n48171), .I1(n8_adj_4030), .I2(n15_adj_4034), 
            .I3(n48273), .O(n48777));   // verilog/motorControl.v(58[19:32])
    defparam i33275_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33276_3_lut (.I0(n48777), .I1(pwm[8]), .I2(pwm_count[8]), 
            .I3(GND_net), .O(n48778));   // verilog/motorControl.v(58[19:32])
    defparam i33276_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i10336_4_lut (.I0(r_SM_Main[2]), .I1(n1_adj_4372), .I2(n28760), 
            .I3(r_SM_Main[1]), .O(n23751));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10336_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i10337_3_lut (.I0(quadB_debounced_adj_3990), .I1(reg_B_adj_4426[0]), 
            .I2(n44576), .I3(GND_net), .O(n23752));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10337_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10341_3_lut (.I0(setpoint[0]), .I1(n3799), .I2(n23533), .I3(GND_net), 
            .O(n23756));   // verilog/coms.v(125[12] 284[6])
    defparam i10341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33651_3_lut (.I0(n49152), .I1(n90), .I2(n41_adj_4155), .I3(GND_net), 
            .O(n49153));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33651_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33596_3_lut (.I0(n49153), .I1(n89), .I2(n43_adj_4156), .I3(GND_net), 
            .O(n49098));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33596_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33247_4_lut (.I0(n43_adj_4156), .I1(n41_adj_4155), .I2(n39_adj_4154), 
            .I3(n47392), .O(n48749));
    defparam i33247_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_12_LessThan_1062_i40_3_lut (.I0(n32_adj_4123), .I1(n91), 
            .I2(n43_adj_4130), .I3(GND_net), .O(n40_adj_4128));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33311_4_lut (.I0(n32_adj_4149), .I1(n24_adj_4141), .I2(n35_adj_4151), 
            .I3(n47396), .O(n48813));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33311_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_12_LessThan_1062_i28_4_lut (.I0(n379), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_12_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(n91), .I1(n22525), .I2(GND_net), .I3(GND_net), 
            .O(n22522));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'hdddd;
    SB_LUT4 i10398_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n28350), 
            .I3(n22470), .O(n23813));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10398_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 div_12_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i33522_3_lut (.I0(n49098), .I1(n88), .I2(n45_adj_4158), .I3(GND_net), 
            .O(n44_adj_4157));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33522_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1470 (.I0(n94), .I1(n22516), .I2(GND_net), .I3(GND_net), 
            .O(n22513));
    defparam i1_2_lut_adj_1470.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i33313_4_lut (.I0(n44_adj_4157), .I1(n48813), .I2(n45_adj_4158), 
            .I3(n48749), .O(n48815));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33313_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1471 (.I0(n48815), .I1(n22537), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1471.LUT_INIT = 16'hceef;
    SB_LUT4 i10399_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n28350), 
            .I3(n22462), .O(n23814));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10399_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i10400_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_3993), 
            .I3(n22470), .O(n23815));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10400_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33453_3_lut (.I0(n28), .I1(n95), .I2(n35_adj_4125), .I3(GND_net), 
            .O(n48955));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33453_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10906_3_lut (.I0(encoder1_position[1]), .I1(n2264), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24321));   // quad.v(35[10] 41[6])
    defparam i10906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1199_3_lut (.I0(n380), .I1(n6795), .I2(n1778), .I3(GND_net), 
            .O(n1874));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10438_3_lut (.I0(n23714), .I1(r_Bit_Index[0]), .I2(n23596), 
            .I3(GND_net), .O(n23853));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10438_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i10434_3_lut (.I0(n23716), .I1(r_Bit_Index_adj_4419[0]), .I2(n23602), 
            .I3(GND_net), .O(n23849));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10434_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_2_lut_adj_1472 (.I0(n97), .I1(n22507), .I2(GND_net), .I3(GND_net), 
            .O(n22504));
    defparam i1_2_lut_adj_1472.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_1473 (.I0(n224), .I1(n99), .I2(n22467), .I3(n558), 
            .O(n5_adj_4374));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i1_4_lut_adj_1473.LUT_INIT = 16'h555d;
    SB_LUT4 i23040_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_3988));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23040_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_i274_4_lut (.I0(n5_adj_4374), .I1(n2_adj_3988), .I2(n392), 
            .I3(n99), .O(n43905));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i274_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_i367_4_lut (.I0(n43905), .I1(n4_adj_3960), .I2(n533), 
            .I3(n98), .O(n43907));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i367_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 div_12_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i23096_3_lut (.I0(n648), .I1(n98), .I2(n4), .I3(GND_net), 
            .O(n6));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23096_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_12_i458_4_lut (.I0(n43907), .I1(n6), .I2(n671), .I3(n97), 
            .O(n43909));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i458_4_lut.LUT_INIT = 16'ha9a6;
    SB_LUT4 i23136_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4037), .I3(GND_net), 
            .O(n8_adj_4036));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23136_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i10833_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24248));   // verilog/coms.v(125[12] 284[6])
    defparam i10833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i547_4_lut (.I0(n43909), .I1(n8_adj_4036), .I2(n806), 
            .I3(n96), .O(n914));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i547_4_lut.LUT_INIT = 16'h5659;
    SB_LUT4 div_12_i634_3_lut (.I0(n914), .I1(n5825), .I2(n938), .I3(GND_net), 
            .O(n1043));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i634_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10834_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24249));   // verilog/coms.v(125[12] 284[6])
    defparam i10834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i719_3_lut (.I0(n1043), .I1(n6217), .I2(n1067), .I3(GND_net), 
            .O(n1169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i802_3_lut (.I0(n1169), .I1(n6578), .I2(n1193), .I3(GND_net), 
            .O(n1292));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i802_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i883_3_lut (.I0(n1292), .I1(n6649), .I2(n1316), .I3(GND_net), 
            .O(n1412));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i883_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i962_3_lut (.I0(n1412), .I1(n6689), .I2(n1436), .I3(GND_net), 
            .O(n1529));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_i1039_3_lut (.I0(n1529), .I1(n6729), .I2(n1553), .I3(GND_net), 
            .O(n1643));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10401_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_3993), 
            .I3(n22462), .O(n23816));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10401_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10431_2_lut (.I0(n23845), .I1(n23844), .I2(GND_net), .I3(GND_net), 
            .O(n23846));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10431_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10402_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_3987), 
            .I3(n22470), .O(n23817));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10402_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10403_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_3987), 
            .I3(n22462), .O(n23818));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10403_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10404_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_3986), 
            .I3(n22470), .O(n23819));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10404_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10825_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24240));   // verilog/coms.v(125[12] 284[6])
    defparam i10825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10802_4_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n5022), .I3(n22429), .O(n24217));   // verilog/coms.v(125[12] 284[6])
    defparam i10802_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i10425_2_lut (.I0(n29726), .I1(n23838), .I2(GND_net), .I3(GND_net), 
            .O(n23840));   // verilog/coms.v(125[12] 284[6])
    defparam i10425_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10422_2_lut (.I0(n29726), .I1(n23835), .I2(GND_net), .I3(GND_net), 
            .O(n23837));   // verilog/coms.v(125[12] 284[6])
    defparam i10422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10805_3_lut (.I0(\data_out_frame[0] [4]), .I1(n5022), .I2(n23563), 
            .I3(GND_net), .O(n24220));   // verilog/coms.v(125[12] 284[6])
    defparam i10805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10419_2_lut (.I0(n29726), .I1(n23832), .I2(GND_net), .I3(GND_net), 
            .O(n23834));   // verilog/coms.v(125[12] 284[6])
    defparam i10419_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10806_3_lut (.I0(\data_out_frame[0] [3]), .I1(n5022), .I2(n23563), 
            .I3(GND_net), .O(n24221));   // verilog/coms.v(125[12] 284[6])
    defparam i10806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10807_3_lut (.I0(\data_out_frame[0] [2]), .I1(n5022), .I2(n23563), 
            .I3(GND_net), .O(n24222));   // verilog/coms.v(125[12] 284[6])
    defparam i10807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10808_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24223));   // verilog/coms.v(125[12] 284[6])
    defparam i10808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10810_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24225));   // verilog/coms.v(125[12] 284[6])
    defparam i10810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10811_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24226));   // verilog/coms.v(125[12] 284[6])
    defparam i10811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10812_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24227));   // verilog/coms.v(125[12] 284[6])
    defparam i10812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10813_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24228));   // verilog/coms.v(125[12] 284[6])
    defparam i10813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_558_i15_2_lut (.I0(pwm_count[7]), .I1(n869), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4044));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_558_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i9_2_lut (.I0(pwm_count[4]), .I1(n872), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4041));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_558_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i13_2_lut (.I0(pwm_count[6]), .I1(n870), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4043));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_558_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_558_i11_2_lut (.I0(pwm_count[5]), .I1(n871), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4042));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_558_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10818_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24233));   // verilog/coms.v(125[12] 284[6])
    defparam i10818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_558_i4_3_lut (.I0(n47156), .I1(n875), .I2(pwm_count[1]), 
            .I3(GND_net), .O(n4_adj_4038));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_558_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33211_3_lut (.I0(n4_adj_4038), .I1(n871), .I2(n11_adj_4042), 
            .I3(GND_net), .O(n48713));   // verilog/motorControl.v(77[28:44])
    defparam i33211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33212_3_lut (.I0(n48713), .I1(n870), .I2(n13_adj_4043), .I3(GND_net), 
            .O(n48714));   // verilog/motorControl.v(77[28:44])
    defparam i33212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32763_4_lut (.I0(n13_adj_4043), .I1(n11_adj_4042), .I2(n9_adj_4041), 
            .I3(n47615), .O(n48265));
    defparam i32763_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i10819_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24234));   // verilog/coms.v(125[12] 284[6])
    defparam i10819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_558_i8_3_lut (.I0(n6_adj_4039), .I1(n872), .I2(n9_adj_4041), 
            .I3(GND_net), .O(n8_adj_4040));   // verilog/motorControl.v(77[28:44])
    defparam LessThan_558_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32695_3_lut (.I0(n48714), .I1(n869), .I2(n15_adj_4044), .I3(GND_net), 
            .O(n48197));   // verilog/motorControl.v(77[28:44])
    defparam i32695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33279_4_lut (.I0(n48197), .I1(n8_adj_4040), .I2(n15_adj_4044), 
            .I3(n48265), .O(n48781));   // verilog/motorControl.v(77[28:44])
    defparam i33279_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33280_3_lut (.I0(n48781), .I1(n868), .I2(pwm_count[8]), .I3(GND_net), 
            .O(n48782));   // verilog/motorControl.v(77[28:44])
    defparam i33280_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33454_3_lut (.I0(n48955), .I1(n94), .I2(n37_adj_4126), .I3(GND_net), 
            .O(n48956));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33454_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10821_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24236));   // verilog/coms.v(125[12] 284[6])
    defparam i10821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10435_3_lut (.I0(encoder0_position[23]), .I1(n2292), .I2(count_enable), 
            .I3(GND_net), .O(n23850));   // quad.v(35[10] 41[6])
    defparam i10435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10439_3_lut (.I0(encoder0_position[22]), .I1(n2293), .I2(count_enable), 
            .I3(GND_net), .O(n23854));   // quad.v(35[10] 41[6])
    defparam i10439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10440_3_lut (.I0(encoder0_position[21]), .I1(n2294), .I2(count_enable), 
            .I3(GND_net), .O(n23855));   // quad.v(35[10] 41[6])
    defparam i10440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31950_4_lut (.I0(n41_adj_4129), .I1(n39_adj_4127), .I2(n37_adj_4126), 
            .I3(n47460), .O(n47450));
    defparam i31950_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i10441_3_lut (.I0(encoder0_position[20]), .I1(n2295), .I2(count_enable), 
            .I3(GND_net), .O(n23856));   // quad.v(35[10] 41[6])
    defparam i10441_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10927_3_lut (.I0(encoder1_position[12]), .I1(n2253), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24342));   // quad.v(35[10] 41[6])
    defparam i10927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10442_3_lut (.I0(encoder0_position[19]), .I1(n2296), .I2(count_enable), 
            .I3(GND_net), .O(n23857));   // quad.v(35[10] 41[6])
    defparam i10442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10443_3_lut (.I0(encoder0_position[18]), .I1(n2297), .I2(count_enable), 
            .I3(GND_net), .O(n23858));   // quad.v(35[10] 41[6])
    defparam i10443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10928_3_lut (.I0(encoder1_position[13]), .I1(n2252), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24343));   // quad.v(35[10] 41[6])
    defparam i10928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10444_3_lut (.I0(encoder0_position[17]), .I1(n2298), .I2(count_enable), 
            .I3(GND_net), .O(n23859));   // quad.v(35[10] 41[6])
    defparam i10444_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10445_3_lut (.I0(encoder0_position[16]), .I1(n2299), .I2(count_enable), 
            .I3(GND_net), .O(n23860));   // quad.v(35[10] 41[6])
    defparam i10445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10446_3_lut (.I0(encoder0_position[15]), .I1(n2300), .I2(count_enable), 
            .I3(GND_net), .O(n23861));   // quad.v(35[10] 41[6])
    defparam i10446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10447_3_lut (.I0(encoder0_position[14]), .I1(n2301), .I2(count_enable), 
            .I3(GND_net), .O(n23862));   // quad.v(35[10] 41[6])
    defparam i10447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33451_4_lut (.I0(n40_adj_4128), .I1(n30_adj_4121), .I2(n43_adj_4130), 
            .I3(n47446), .O(n48953));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33451_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i10929_3_lut (.I0(encoder1_position[14]), .I1(n2251), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24344));   // quad.v(35[10] 41[6])
    defparam i10929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10448_3_lut (.I0(encoder0_position[13]), .I1(n2302), .I2(count_enable), 
            .I3(GND_net), .O(n23863));   // quad.v(35[10] 41[6])
    defparam i10448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10930_3_lut (.I0(encoder1_position[15]), .I1(n2250), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24345));   // quad.v(35[10] 41[6])
    defparam i10930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10931_3_lut (.I0(encoder1_position[16]), .I1(n2249), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24346));   // quad.v(35[10] 41[6])
    defparam i10931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10449_3_lut (.I0(encoder0_position[12]), .I1(n2303), .I2(count_enable), 
            .I3(GND_net), .O(n23864));   // quad.v(35[10] 41[6])
    defparam i10449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10450_3_lut (.I0(encoder0_position[11]), .I1(n2304), .I2(count_enable), 
            .I3(GND_net), .O(n23865));   // quad.v(35[10] 41[6])
    defparam i10450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10451_3_lut (.I0(encoder0_position[10]), .I1(n2305), .I2(count_enable), 
            .I3(GND_net), .O(n23866));   // quad.v(35[10] 41[6])
    defparam i10451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10452_3_lut (.I0(encoder0_position[9]), .I1(n2306), .I2(count_enable), 
            .I3(GND_net), .O(n23867));   // quad.v(35[10] 41[6])
    defparam i10452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10932_3_lut (.I0(encoder1_position[17]), .I1(n2248), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24347));   // quad.v(35[10] 41[6])
    defparam i10932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33302_3_lut (.I0(n48956), .I1(n93), .I2(n39_adj_4127), .I3(GND_net), 
            .O(n48804));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33302_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i10453_3_lut (.I0(encoder0_position[8]), .I1(n2307), .I2(count_enable), 
            .I3(GND_net), .O(n23868));   // quad.v(35[10] 41[6])
    defparam i10453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10933_3_lut (.I0(encoder1_position[18]), .I1(n2247), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24348));   // quad.v(35[10] 41[6])
    defparam i10933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10454_3_lut (.I0(encoder0_position[7]), .I1(n2308), .I2(count_enable), 
            .I3(GND_net), .O(n23869));   // quad.v(35[10] 41[6])
    defparam i10454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10934_3_lut (.I0(encoder1_position[19]), .I1(n2246), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24349));   // quad.v(35[10] 41[6])
    defparam i10934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10455_3_lut (.I0(encoder0_position[6]), .I1(n2309), .I2(count_enable), 
            .I3(GND_net), .O(n23870));   // quad.v(35[10] 41[6])
    defparam i10455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10456_3_lut (.I0(encoder0_position[5]), .I1(n2310), .I2(count_enable), 
            .I3(GND_net), .O(n23871));   // quad.v(35[10] 41[6])
    defparam i10456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10457_3_lut (.I0(encoder0_position[4]), .I1(n2311), .I2(count_enable), 
            .I3(GND_net), .O(n23872));   // quad.v(35[10] 41[6])
    defparam i10457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10458_3_lut (.I0(encoder0_position[3]), .I1(n2312), .I2(count_enable), 
            .I3(GND_net), .O(n23873));   // quad.v(35[10] 41[6])
    defparam i10458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10935_3_lut (.I0(encoder1_position[20]), .I1(n2245), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24350));   // quad.v(35[10] 41[6])
    defparam i10935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10459_3_lut (.I0(encoder0_position[2]), .I1(n2313), .I2(count_enable), 
            .I3(GND_net), .O(n23874));   // quad.v(35[10] 41[6])
    defparam i10459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10936_3_lut (.I0(encoder1_position[21]), .I1(n2244), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24351));   // quad.v(35[10] 41[6])
    defparam i10936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10937_3_lut (.I0(encoder1_position[22]), .I1(n2243), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24352));   // quad.v(35[10] 41[6])
    defparam i10937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10460_3_lut (.I0(encoder0_position[1]), .I1(n2314), .I2(count_enable), 
            .I3(GND_net), .O(n23875));   // quad.v(35[10] 41[6])
    defparam i10460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10938_3_lut (.I0(encoder1_position[23]), .I1(n2242), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24353));   // quad.v(35[10] 41[6])
    defparam i10938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1474 (.I0(n103), .I1(n22458), .I2(n5_adj_4375), 
            .I3(n122), .O(n7_adj_4373));   // verilog/coms.v(125[12] 284[6])
    defparam i2_4_lut_adj_1474.LUT_INIT = 16'hb333;
    SB_LUT4 i4_4_lut_adj_1475 (.I0(n7_adj_4373), .I1(n44586), .I2(n5_adj_4011), 
            .I3(n7_adj_4012), .O(n50101));   // verilog/coms.v(125[12] 284[6])
    defparam i4_4_lut_adj_1475.LUT_INIT = 16'hfffe;
    SB_LUT4 i10462_3_lut (.I0(\PID_CONTROLLER.err_prev [31]), .I1(\PID_CONTROLLER.err [31]), 
            .I2(n44626), .I3(GND_net), .O(n23877));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10462_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10463_3_lut (.I0(\PID_CONTROLLER.err_prev [23]), .I1(\PID_CONTROLLER.err [23]), 
            .I2(n44626), .I3(GND_net), .O(n23878));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10464_3_lut (.I0(\PID_CONTROLLER.err_prev [22]), .I1(\PID_CONTROLLER.err [22]), 
            .I2(n44626), .I3(GND_net), .O(n23879));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10465_3_lut (.I0(\PID_CONTROLLER.err_prev [21]), .I1(\PID_CONTROLLER.err [21]), 
            .I2(n44626), .I3(GND_net), .O(n23880));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10466_3_lut (.I0(\PID_CONTROLLER.err_prev [20]), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n44626), .I3(GND_net), .O(n23881));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10942_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_3986), 
            .I3(n22462), .O(n24357));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10942_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10467_3_lut (.I0(\PID_CONTROLLER.err_prev [19]), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n44626), .I3(GND_net), .O(n23882));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10943_4_lut (.I0(pwm_23__N_2948), .I1(n471), .I2(PWMLimit[0]), 
            .I3(n387), .O(n24358));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10943_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10468_3_lut (.I0(\PID_CONTROLLER.err_prev [18]), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n44626), .I3(GND_net), .O(n23883));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10944_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n44902), 
            .I3(GND_net), .O(n24359));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i10944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34444_4_lut (.I0(r_SM_Main[2]), .I1(n47206), .I2(n47207), 
            .I3(r_SM_Main[1]), .O(n28794));
    defparam i34444_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 i10407_2_lut (.I0(n29726), .I1(n23820), .I2(GND_net), .I3(GND_net), 
            .O(n23822));   // verilog/coms.v(125[12] 284[6])
    defparam i10407_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10469_3_lut (.I0(\PID_CONTROLLER.err_prev [17]), .I1(\PID_CONTROLLER.err [17]), 
            .I2(n44626), .I3(GND_net), .O(n23884));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10469_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10470_3_lut (.I0(\PID_CONTROLLER.err_prev [16]), .I1(\PID_CONTROLLER.err [16]), 
            .I2(n44626), .I3(GND_net), .O(n23885));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10470_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10947_4_lut (.I0(pwm_23__N_2948), .I1(n470), .I2(PWMLimit[1]), 
            .I3(n387), .O(n24362));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10947_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10471_3_lut (.I0(\PID_CONTROLLER.err_prev [15]), .I1(\PID_CONTROLLER.err [15]), 
            .I2(n44626), .I3(GND_net), .O(n23886));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10948_4_lut (.I0(pwm_23__N_2948), .I1(n469), .I2(PWMLimit[2]), 
            .I3(n387), .O(n24363));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10948_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10472_3_lut (.I0(\PID_CONTROLLER.err_prev [14]), .I1(\PID_CONTROLLER.err [14]), 
            .I2(n44626), .I3(GND_net), .O(n23887));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10472_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10473_3_lut (.I0(\PID_CONTROLLER.err_prev [13]), .I1(\PID_CONTROLLER.err [13]), 
            .I2(n44626), .I3(GND_net), .O(n23888));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10473_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10474_3_lut (.I0(\PID_CONTROLLER.err_prev [12]), .I1(\PID_CONTROLLER.err [12]), 
            .I2(n44626), .I3(GND_net), .O(n23889));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10474_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10949_4_lut (.I0(pwm_23__N_2948), .I1(n468), .I2(PWMLimit[3]), 
            .I3(n387), .O(n24364));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10949_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10475_3_lut (.I0(\PID_CONTROLLER.err_prev [11]), .I1(\PID_CONTROLLER.err [11]), 
            .I2(n44626), .I3(GND_net), .O(n23890));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10475_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10476_3_lut (.I0(\PID_CONTROLLER.err_prev [10]), .I1(\PID_CONTROLLER.err [10]), 
            .I2(n44626), .I3(GND_net), .O(n23891));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10476_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10477_3_lut (.I0(\PID_CONTROLLER.err_prev [9]), .I1(\PID_CONTROLLER.err [9]), 
            .I2(n44626), .I3(GND_net), .O(n23892));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10477_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10950_4_lut (.I0(pwm_23__N_2948), .I1(n467), .I2(PWMLimit[4]), 
            .I3(n387), .O(n24365));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10950_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i5_3_lut (.I0(\PID_CONTROLLER.result [5]), .I1(n415), .I2(n421), 
            .I3(GND_net), .O(n1_adj_4026));
    defparam i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10478_3_lut (.I0(\PID_CONTROLLER.err_prev [8]), .I1(\PID_CONTROLLER.err [8]), 
            .I2(n44626), .I3(GND_net), .O(n23893));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10478_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10479_3_lut (.I0(\PID_CONTROLLER.err_prev [7]), .I1(\PID_CONTROLLER.err [7]), 
            .I2(n44626), .I3(GND_net), .O(n23894));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10479_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10480_3_lut (.I0(\PID_CONTROLLER.err_prev [6]), .I1(\PID_CONTROLLER.err [6]), 
            .I2(n44626), .I3(GND_net), .O(n23895));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10480_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14653_3_lut (.I0(\PID_CONTROLLER.result [6]), .I1(n414), .I2(n421), 
            .I3(GND_net), .O(n28052));
    defparam i14653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10481_3_lut (.I0(\PID_CONTROLLER.err_prev [5]), .I1(\PID_CONTROLLER.err [5]), 
            .I2(n44626), .I3(GND_net), .O(n23896));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10481_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10482_3_lut (.I0(\PID_CONTROLLER.err_prev [4]), .I1(\PID_CONTROLLER.err [4]), 
            .I2(n44626), .I3(GND_net), .O(n23897));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10482_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_3_lut_adj_1476 (.I0(\PID_CONTROLLER.result [7]), .I1(n413), 
            .I2(n421), .I3(GND_net), .O(n1));
    defparam i5_3_lut_adj_1476.LUT_INIT = 16'hcaca;
    SB_LUT4 i10483_3_lut (.I0(\PID_CONTROLLER.err_prev [3]), .I1(\PID_CONTROLLER.err [3]), 
            .I2(n44626), .I3(GND_net), .O(n23898));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10483_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10484_3_lut (.I0(\PID_CONTROLLER.err_prev [2]), .I1(\PID_CONTROLLER.err [2]), 
            .I2(n44626), .I3(GND_net), .O(n23899));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10484_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10954_4_lut (.I0(pwm_23__N_2948), .I1(n463), .I2(PWMLimit[8]), 
            .I3(n387), .O(n24369));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10954_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10485_3_lut (.I0(\PID_CONTROLLER.err_prev [1]), .I1(\PID_CONTROLLER.err [1]), 
            .I2(n44626), .I3(GND_net), .O(n23900));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10485_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10955_4_lut (.I0(pwm_23__N_2948), .I1(n462), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24370));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10955_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10956_4_lut (.I0(pwm_23__N_2948), .I1(n461), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24371));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10956_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10957_4_lut (.I0(pwm_23__N_2948), .I1(n460), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24372));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10957_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10958_4_lut (.I0(pwm_23__N_2948), .I1(n459), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24373));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10958_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10959_4_lut (.I0(pwm_23__N_2948), .I1(n458), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24374));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10959_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10502_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n43238), .I3(GND_net), .O(n23917));   // verilog/coms.v(125[12] 284[6])
    defparam i10502_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10503_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n43238), .I3(GND_net), .O(n23918));   // verilog/coms.v(125[12] 284[6])
    defparam i10503_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10960_4_lut (.I0(pwm_23__N_2948), .I1(n457), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24375));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10960_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10504_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n43238), .I3(GND_net), .O(n23919));   // verilog/coms.v(125[12] 284[6])
    defparam i10504_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10961_4_lut (.I0(pwm_23__N_2948), .I1(n456), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24376));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10961_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10505_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n43238), .I3(GND_net), .O(n23920));   // verilog/coms.v(125[12] 284[6])
    defparam i10505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10962_4_lut (.I0(pwm_23__N_2948), .I1(n455), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24377));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10962_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1477 (.I0(pwm_23__N_2948), .I1(n47225), .I2(PWMLimit[9]), 
            .I3(n387), .O(n42011));   // verilog/motorControl.v(31[14] 52[8])
    defparam i1_4_lut_adj_1477.LUT_INIT = 16'ha088;
    SB_LUT4 i10506_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n43238), .I3(GND_net), .O(n23921));   // verilog/coms.v(125[12] 284[6])
    defparam i10506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10965_4_lut (.I0(pwm_23__N_2948), .I1(n47180), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24380));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10965_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10507_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n43238), .I3(GND_net), .O(n23922));   // verilog/coms.v(125[12] 284[6])
    defparam i10507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10508_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n43238), .I3(GND_net), .O(n23923));   // verilog/coms.v(125[12] 284[6])
    defparam i10508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10966_4_lut (.I0(pwm_23__N_2948), .I1(n47182), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24381));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10966_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10509_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n43238), .I3(GND_net), .O(n23924));   // verilog/coms.v(125[12] 284[6])
    defparam i10509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10967_4_lut (.I0(pwm_23__N_2948), .I1(n47184), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24382));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10967_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i10968_4_lut (.I0(pwm_23__N_2948), .I1(n47186), .I2(PWMLimit[9]), 
            .I3(n387), .O(n24383));   // verilog/motorControl.v(31[14] 52[8])
    defparam i10968_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i15_2_lut (.I0(pwm_23__N_2951[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4019));   // verilog/motorControl.v(25[23:29])
    defparam i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i20_2_lut (.I0(deadband[5]), .I1(\PID_CONTROLLER.result [5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4014));   // verilog/motorControl.v(25[23:29])
    defparam i20_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_2_lut (.I0(deadband[6]), .I1(\PID_CONTROLLER.result [6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4015));   // verilog/motorControl.v(25[23:29])
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10518_3_lut (.I0(\data_in_frame[19] [7]), .I1(rx_data[7]), 
            .I2(n43236), .I3(GND_net), .O(n23933));   // verilog/coms.v(125[12] 284[6])
    defparam i10518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20_2_lut_adj_1478 (.I0(deadband[7]), .I1(\PID_CONTROLLER.result [7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4016));   // verilog/motorControl.v(25[23:29])
    defparam i20_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i10519_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n43236), .I3(GND_net), .O(n23934));   // verilog/coms.v(125[12] 284[6])
    defparam i10519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10520_3_lut (.I0(\data_in_frame[19] [5]), .I1(rx_data[5]), 
            .I2(n43236), .I3(GND_net), .O(n23935));   // verilog/coms.v(125[12] 284[6])
    defparam i10520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10521_3_lut (.I0(\data_in_frame[19] [4]), .I1(rx_data[4]), 
            .I2(n43236), .I3(GND_net), .O(n23936));   // verilog/coms.v(125[12] 284[6])
    defparam i10521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10522_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n43236), .I3(GND_net), .O(n23937));   // verilog/coms.v(125[12] 284[6])
    defparam i10522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10523_3_lut (.I0(\data_in_frame[19] [2]), .I1(rx_data[2]), 
            .I2(n43236), .I3(GND_net), .O(n23938));   // verilog/coms.v(125[12] 284[6])
    defparam i10523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10524_3_lut (.I0(\data_in_frame[19] [1]), .I1(rx_data[1]), 
            .I2(n43236), .I3(GND_net), .O(n23939));   // verilog/coms.v(125[12] 284[6])
    defparam i10524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10525_3_lut (.I0(\data_in_frame[19] [0]), .I1(rx_data[0]), 
            .I2(n43236), .I3(GND_net), .O(n23940));   // verilog/coms.v(125[12] 284[6])
    defparam i10525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10550_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n43255), .I3(GND_net), .O(n23965));   // verilog/coms.v(125[12] 284[6])
    defparam i10550_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33688_4_lut (.I0(n48804), .I1(n48953), .I2(n43_adj_4130), 
            .I3(n47450), .O(n49190));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33688_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33689_3_lut (.I0(n49190), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n49191));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33689_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_12_i1332_3_lut_3_lut (.I0(n1991), .I1(n6845), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_23_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[0]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_25[0]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_555_i6_3_lut_3_lut (.I0(pwm_count[3]), .I1(pwm[3]), 
            .I2(pwm[2]), .I3(GND_net), .O(n6_adj_4029));   // verilog/motorControl.v(58[19:32])
    defparam LessThan_555_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i32122_3_lut_4_lut (.I0(pwm_count[3]), .I1(pwm[3]), .I2(pwm[2]), 
            .I3(pwm_count[2]), .O(n47623));   // verilog/motorControl.v(58[19:32])
    defparam i32122_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i32028_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n47529));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32028_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4107));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 mux_23_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[1]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_25[1]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32042_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n47543));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32042_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 mux_23_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[2]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_25[2]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4101));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 mux_23_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[3]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_25[3]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4099));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32056_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n47557));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32056_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4097));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32070_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n47571));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32070_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4095));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32088_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n47589));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32088_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i1_4_lut_adj_1479 (.I0(n49191), .I1(n22531), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1479.LUT_INIT = 16'hceef;
    SB_LUT4 i10551_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n43255), .I3(GND_net), .O(n23966));   // verilog/coms.v(125[12] 284[6])
    defparam i10551_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10552_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n43255), .I3(GND_net), .O(n23967));   // verilog/coms.v(125[12] 284[6])
    defparam i10552_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10553_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n43255), .I3(GND_net), .O(n23968));   // verilog/coms.v(125[12] 284[6])
    defparam i10553_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10554_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n43255), .I3(GND_net), .O(n23969));   // verilog/coms.v(125[12] 284[6])
    defparam i10554_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10555_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n43255), .I3(GND_net), .O(n23970));   // verilog/coms.v(125[12] 284[6])
    defparam i10555_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10556_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n43255), .I3(GND_net), .O(n23971));   // verilog/coms.v(125[12] 284[6])
    defparam i10556_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10557_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n43255), .I3(GND_net), .O(n23972));   // verilog/coms.v(125[12] 284[6])
    defparam i10557_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_23_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[4]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_25[4]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[5]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_25[5]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[6]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_25[6]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4196));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31782_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n47282));
    defparam i31782_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i1333_3_lut_3_lut (.I0(n1991), .I1(n6846), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4198));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_4200));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31788_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n47288));
    defparam i31788_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4217));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32336_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n47838));
    defparam i32336_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4219));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_4221));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31752_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n47252));
    defparam i31752_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4235));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32293_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n47795));
    defparam i32293_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4237));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_4239));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32271_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n47773));
    defparam i32271_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_i1040_3_lut (.I0(n1530), .I1(n6730), .I2(n1553), .I3(GND_net), 
            .O(n1644));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4241));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_4_lut (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n22555));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1480 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n22558));
    defparam i1_2_lut_3_lut_adj_1480.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4257));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32253_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n47755));
    defparam i32253_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4259));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_4261));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32216_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n47718));
    defparam i32216_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4263));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n89), .I1(n88), .I2(n87), .I3(n22537), 
            .O(n22528));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 div_12_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4279));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32188_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n47690));
    defparam i32188_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4281));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 mux_23_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[7]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_25[7]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10826_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24241));   // verilog/coms.v(125[12] 284[6])
    defparam i10826_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[8]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_25[8]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[9]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_25[9]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[10]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_25[10]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[11]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_25[11]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_4283));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    SB_LUT4 i32127_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n47628));
    defparam i32127_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4285));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 mux_23_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[12]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_25[12]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[13]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_25[13]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[14]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_25[14]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[15]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_25[15]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[16]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_25[16]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[17]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_25[17]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10566_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n43253), .I3(GND_net), .O(n23981));   // verilog/coms.v(125[12] 284[6])
    defparam i10566_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_23_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[18]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_25[18]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[19]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_25[19]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_23_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[20]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_25[20]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10567_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n43253), .I3(GND_net), .O(n23982));   // verilog/coms.v(125[12] 284[6])
    defparam i10567_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10568_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n43253), .I3(GND_net), .O(n23983));   // verilog/coms.v(125[12] 284[6])
    defparam i10568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_23_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[21]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_25[21]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10569_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n43253), .I3(GND_net), .O(n23984));   // verilog/coms.v(125[12] 284[6])
    defparam i10569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10570_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n43253), .I3(GND_net), .O(n23985));   // verilog/coms.v(125[12] 284[6])
    defparam i10570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10571_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n43253), .I3(GND_net), .O(n23986));   // verilog/coms.v(125[12] 284[6])
    defparam i10571_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10572_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n43253), .I3(GND_net), .O(n23987));   // verilog/coms.v(125[12] 284[6])
    defparam i10572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4301));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10573_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n43253), .I3(GND_net), .O(n23988));   // verilog/coms.v(125[12] 284[6])
    defparam i10573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_4305));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31994_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n47494));
    defparam i31994_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4307));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4303));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i32080_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n47581));
    defparam i32080_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4323));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_4327));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31894_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n47394));
    defparam i31894_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i10582_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n43251), .I3(GND_net), .O(n23997));   // verilog/coms.v(125[12] 284[6])
    defparam i10582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10583_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n43251), .I3(GND_net), .O(n23998));   // verilog/coms.v(125[12] 284[6])
    defparam i10583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10584_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n43251), .I3(GND_net), .O(n23999));   // verilog/coms.v(125[12] 284[6])
    defparam i10584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10585_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n43251), .I3(GND_net), .O(n24000));   // verilog/coms.v(125[12] 284[6])
    defparam i10585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10586_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n43251), .I3(GND_net), .O(n24001));   // verilog/coms.v(125[12] 284[6])
    defparam i10586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10587_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n43251), .I3(GND_net), .O(n24002));   // verilog/coms.v(125[12] 284[6])
    defparam i10587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10588_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n43251), .I3(GND_net), .O(n24003));   // verilog/coms.v(125[12] 284[6])
    defparam i10588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_12_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4329));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4325));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i10589_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n43251), .I3(GND_net), .O(n24004));   // verilog/coms.v(125[12] 284[6])
    defparam i10589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31942_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n47442));
    defparam i31942_2_lut_4_lut.LUT_INIT = 16'hf99f;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n24341(n24341), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n24340(n24340), .n24339(n24339), .n24353(n24353), 
            .n24352(n24352), .n24351(n24351), .n24350(n24350), .n24349(n24349), 
            .n24348(n24348), .n24347(n24347), .n24346(n24346), .n24345(n24345), 
            .n24344(n24344), .n24343(n24343), .n24342(n24342), .n24338(n24338), 
            .n24337(n24337), .data_o({quadA_debounced_adj_3989, quadB_debounced_adj_3990}), 
            .n24336(n24336), .n24335(n24335), .n24334(n24334), .n24333(n24333), 
            .n24332(n24332), .n2241({n2242, n2243, n2244, n2245, n2246, 
            n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, 
            n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
            n2263, n2264, n2265}), .GND_net(GND_net), .n24321(n24321), 
            .n23746(n23746), .count_enable(count_enable_adj_3991), .n24385(n24385), 
            .n44576(n44576), .reg_B({reg_B_adj_4426}), .PIN_18_c_1(PIN_18_c_1), 
            .PIN_19_c_0(PIN_19_c_0), .n23752(n23752)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(174[15] 179[4])
    SB_LUT4 mux_23_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[22]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_25[22]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1481 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4013));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i4_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1482 (.I0(control_mode[6]), .I1(n10_adj_4013), 
            .I2(control_mode[2]), .I3(GND_net), .O(n22459));   // verilog/TinyFPGA_B.v(137[5:22])
    defparam i5_3_lut_adj_1482.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1483 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n22459), .I3(GND_net), .O(n15_adj_3964));   // verilog/TinyFPGA_B.v(138[5:22])
    defparam i2_3_lut_adj_1483.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_23_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_3964), .I3(n15_adj_3965), .O(motor_state_23__N_25[23]));   // verilog/TinyFPGA_B.v(138[5] 141[10])
    defparam mux_23_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_22_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_25[23]), 
            .I2(n15_adj_3992), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(137[5] 141[10])
    defparam mux_22_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_3966));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_3967));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_3968));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_3969));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_3970));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_3971));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_3972));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_3973));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_3974));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_3975));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_3976));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_3977));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_3978));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_3979));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_3980));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10410_2_lut (.I0(n29726), .I1(n23823), .I2(GND_net), .I3(GND_net), 
            .O(n23825));   // verilog/coms.v(125[12] 284[6])
    defparam i10410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10917_3_lut (.I0(encoder1_position[2]), .I1(n2263), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24332));   // quad.v(35[10] 41[6])
    defparam i10917_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10918_3_lut (.I0(encoder1_position[3]), .I1(n2262), .I2(count_enable_adj_3991), 
            .I3(GND_net), .O(n24333));   // quad.v(35[10] 41[6])
    defparam i10918_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_3981));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_3982));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_3983));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_3984));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n7007), 
            .I3(n2724), .O(n41_adj_4369));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n7008), 
            .I3(n2724), .O(n39_adj_4367));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n391));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n7005), 
            .I3(n2724), .O(n45_adj_4371));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n7006), 
            .I3(n2724), .O(n43_adj_4370));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n7009), 
            .I3(n2724), .O(n37_adj_4366));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n7013), 
            .I3(n2724), .O(n29_adj_4361));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n7012), 
            .I3(n2724), .O(n31_adj_4363));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n7017), 
            .I3(n2724), .O(n21_adj_4356));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n7016), 
            .I3(n2724), .O(n23_adj_4357));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n7015), 
            .I3(n2724), .O(n25_adj_4359));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n7019), 
            .I3(n2724), .O(n17_adj_4354));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n7018), 
            .I3(n2724), .O(n19_adj_4355));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n7023), 
            .I3(n2724), .O(n9_adj_4347));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n7024), 
            .I3(n2724), .O(n7_adj_4345));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n7011), 
            .I3(n2724), .O(n33_adj_4364));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n7022), 
            .I3(n2724), .O(n11_adj_4349));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n7021), 
            .I3(n2724), .O(n13_adj_4351));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n7020), 
            .I3(n2724), .O(n15_adj_4352));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n7014), 
            .I3(n2724), .O(n27_adj_4360));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n7010), 
            .I3(n2724), .O(n35_adj_4365));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_12_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31818_4_lut (.I0(n27_adj_4360), .I1(n15_adj_4352), .I2(n13_adj_4351), 
            .I3(n11_adj_4349), .O(n47318));
    defparam i31818_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4364), 
            .I3(GND_net), .O(n12_adj_4350));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i31804_2_lut (.I0(n33_adj_4364), .I1(n15_adj_4352), .I2(GND_net), 
            .I3(GND_net), .O(n47304));
    defparam i31804_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_4351), 
            .I3(GND_net), .O(n10_adj_4348));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1830_i30_3_lut (.I0(n12_adj_4350), .I1(n83), 
            .I2(n35_adj_4365), .I3(GND_net), .O(n30_adj_4362));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1828_3_lut (.I0(n2720), .I1(n7025), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31857_3_lut (.I0(n7_adj_4345), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n47357));
    defparam i31857_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i32538_4_lut (.I0(n13_adj_4351), .I1(n11_adj_4349), .I2(n9_adj_4347), 
            .I3(n47357), .O(n48040));
    defparam i32538_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32530_4_lut (.I0(n19_adj_4355), .I1(n17_adj_4354), .I2(n15_adj_4352), 
            .I3(n48040), .O(n48032));
    defparam i32530_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33491_4_lut (.I0(n25_adj_4359), .I1(n23_adj_4357), .I2(n21_adj_4356), 
            .I3(n48032), .O(n48993));
    defparam i33491_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33006_4_lut (.I0(n31_adj_4363), .I1(n29_adj_4361), .I2(n27_adj_4360), 
            .I3(n48993), .O(n48508));
    defparam i33006_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33619_4_lut (.I0(n37_adj_4366), .I1(n35_adj_4365), .I2(n33_adj_4364), 
            .I3(n48508), .O(n49121));
    defparam i33619_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_12_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4370), 
            .I3(GND_net), .O(n16_adj_4353));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4345), 
            .I3(GND_net), .O(n6_adj_4344));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i33417_3_lut (.I0(n6_adj_4344), .I1(n90), .I2(n21_adj_4356), 
            .I3(GND_net), .O(n48919));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33417_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33418_3_lut (.I0(n48919), .I1(n89), .I2(n23_adj_4357), .I3(GND_net), 
            .O(n48920));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33418_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31835_4_lut (.I0(n21_adj_4356), .I1(n19_adj_4355), .I2(n17_adj_4354), 
            .I3(n9_adj_4347), .O(n47335));
    defparam i31835_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31766_2_lut (.I0(n43_adj_4370), .I1(n19_adj_4355), .I2(GND_net), 
            .I3(GND_net), .O(n47266));
    defparam i31766_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_12_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4354), 
            .I3(GND_net), .O(n8_adj_4346));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_LessThan_1830_i24_3_lut (.I0(n16_adj_4353), .I1(n78), 
            .I2(n45_adj_4371), .I3(GND_net), .O(n24_adj_4358));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31774_4_lut (.I0(n43_adj_4370), .I1(n25_adj_4359), .I2(n23_adj_4357), 
            .I3(n47335), .O(n47274));
    defparam i31774_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33365_4_lut (.I0(n24_adj_4358), .I1(n8_adj_4346), .I2(n45_adj_4371), 
            .I3(n47266), .O(n48867));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33365_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_12_i1270_3_lut (.I0(n1874), .I1(n6836), .I2(n1886), .I3(GND_net), 
            .O(n1979));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33360_3_lut (.I0(n48920), .I1(n88), .I2(n25_adj_4359), .I3(GND_net), 
            .O(n48862));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33360_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1829_3_lut (.I0(n390), .I1(n7026), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1830_i4_4_lut (.I0(n391), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4343));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33415_3_lut (.I0(n4_adj_4343), .I1(n87), .I2(n27_adj_4360), 
            .I3(GND_net), .O(n48917));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33415_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33416_3_lut (.I0(n48917), .I1(n86), .I2(n29_adj_4361), .I3(GND_net), 
            .O(n48918));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33416_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31808_4_lut (.I0(n33_adj_4364), .I1(n31_adj_4363), .I2(n29_adj_4361), 
            .I3(n47318), .O(n47308));
    defparam i31808_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33664_4_lut (.I0(n30_adj_4362), .I1(n10_adj_4348), .I2(n35_adj_4365), 
            .I3(n47304), .O(n49166));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33664_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33362_3_lut (.I0(n48918), .I1(n85), .I2(n31_adj_4363), .I3(GND_net), 
            .O(n48864));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33362_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33751_4_lut (.I0(n48864), .I1(n49166), .I2(n35_adj_4365), 
            .I3(n47308), .O(n49253));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33751_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33752_3_lut (.I0(n49253), .I1(n82), .I2(n37_adj_4366), .I3(GND_net), 
            .O(n49254));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33752_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33710_3_lut (.I0(n49254), .I1(n81), .I2(n39_adj_4367), .I3(GND_net), 
            .O(n49212));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33710_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31776_4_lut (.I0(n43_adj_4370), .I1(n41_adj_4369), .I2(n39_adj_4367), 
            .I3(n49121), .O(n47276));
    defparam i31776_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33541_4_lut (.I0(n48862), .I1(n48867), .I2(n45_adj_4371), 
            .I3(n47274), .O(n49043));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33541_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33700_3_lut (.I0(n49212), .I1(n80), .I2(n41_adj_4369), .I3(GND_net), 
            .O(n40_adj_4368));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33700_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1807_3_lut (.I0(n2699), .I1(n7004), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33543_4_lut (.I0(n40_adj_4368), .I1(n49043), .I2(n45_adj_4371), 
            .I3(n47276), .O(n49045));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33543_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33544_3_lut (.I0(n49045), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33544_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_3985));   // verilog/TinyFPGA_B.v(162[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_i1269_3_lut_3_lut (.I0(n1886), .I1(n6835), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1265_3_lut_3_lut (.I0(n1886), .I1(n6831), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4340));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4338));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4342));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4341));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n390));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4335));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4336));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4324));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4333));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4334));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4328));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4330));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4331));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4337));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4326));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1264_3_lut_3_lut (.I0(n1886), .I1(n6830), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4332));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31919_4_lut (.I0(n29_adj_4337), .I1(n17_adj_4331), .I2(n15_adj_4330), 
            .I3(n13_adj_4328), .O(n47419));
    defparam i31919_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32614_4_lut (.I0(n11_adj_4326), .I1(n9_adj_4324), .I2(n2719), 
            .I3(n98), .O(n48116));
    defparam i32614_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i33046_4_lut (.I0(n17_adj_4331), .I1(n15_adj_4330), .I2(n13_adj_4328), 
            .I3(n48116), .O(n48548));
    defparam i33046_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33042_4_lut (.I0(n23_adj_4334), .I1(n21_adj_4333), .I2(n19_adj_4332), 
            .I3(n48548), .O(n48544));
    defparam i33042_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i31923_4_lut (.I0(n29_adj_4337), .I1(n27_adj_4336), .I2(n25_adj_4335), 
            .I3(n48544), .O(n47423));
    defparam i31923_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1777_i6_4_lut (.I0(n390), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4322));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33423_3_lut (.I0(n6_adj_4322), .I1(n87), .I2(n29_adj_4337), 
            .I3(GND_net), .O(n48925));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33423_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1777_i32_3_lut (.I0(n14_adj_4329), .I1(n83), 
            .I2(n37_adj_4342), .I3(GND_net), .O(n32_adj_4339));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33424_3_lut (.I0(n48925), .I1(n86), .I2(n31_adj_4338), .I3(GND_net), 
            .O(n48926));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33424_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31911_4_lut (.I0(n35_adj_4341), .I1(n33_adj_4340), .I2(n31_adj_4338), 
            .I3(n47419), .O(n47411));
    defparam i31911_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33662_4_lut (.I0(n32_adj_4339), .I1(n12_adj_4327), .I2(n37_adj_4342), 
            .I3(n47394), .O(n49164));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33662_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33352_3_lut (.I0(n48926), .I1(n85), .I2(n33_adj_4340), .I3(GND_net), 
            .O(n48854));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33352_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33425_3_lut (.I0(n8_adj_4323), .I1(n90), .I2(n23_adj_4334), 
            .I3(GND_net), .O(n48927));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33425_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33426_3_lut (.I0(n48927), .I1(n89), .I2(n25_adj_4335), .I3(GND_net), 
            .O(n48928));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33426_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32594_4_lut (.I0(n25_adj_4335), .I1(n23_adj_4334), .I2(n21_adj_4333), 
            .I3(n47442), .O(n48096));
    defparam i32594_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33349_3_lut (.I0(n10_adj_4325), .I1(n91), .I2(n21_adj_4333), 
            .I3(GND_net), .O(n48851));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33349_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33348_3_lut (.I0(n48928), .I1(n88), .I2(n27_adj_4336), .I3(GND_net), 
            .O(n48850));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33348_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1268_3_lut_3_lut (.I0(n1886), .I1(n6834), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33251_4_lut (.I0(n35_adj_4341), .I1(n33_adj_4340), .I2(n31_adj_4338), 
            .I3(n47423), .O(n48753));
    defparam i33251_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33749_4_lut (.I0(n48854), .I1(n49164), .I2(n37_adj_4342), 
            .I3(n47411), .O(n49251));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33749_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33419_4_lut (.I0(n48850), .I1(n48851), .I2(n27_adj_4336), 
            .I3(n48096), .O(n48921));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33419_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33763_4_lut (.I0(n48921), .I1(n49251), .I2(n37_adj_4342), 
            .I3(n48753), .O(n49265));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33763_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33764_3_lut (.I0(n49265), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n49266));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33764_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33758_3_lut (.I0(n49266), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n49260));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33758_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33613_3_lut (.I0(n49260), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n49115));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33613_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33614_3_lut (.I0(n49115), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n49116));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33614_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1834_4_lut (.I0(n49116), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1834_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4319));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4321));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4317));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n389));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4320));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4314));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4315));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4302));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4312));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4313));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4304));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1267_3_lut_3_lut (.I0(n1886), .I1(n6833), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i23064_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n370), .I3(n558), 
            .O(n4_adj_3960));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23064_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i1_2_lut_3_lut_adj_1484 (.I0(n98), .I1(n97), .I2(n22507), 
            .I3(GND_net), .O(n22467));
    defparam i1_2_lut_3_lut_adj_1484.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4306));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4308));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4309));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4316));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4311));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32038_4_lut (.I0(n31_adj_4316), .I1(n19_adj_4309), .I2(n17_adj_4308), 
            .I3(n15_adj_4306), .O(n47539));
    defparam i32038_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32757_4_lut (.I0(n13_adj_4304), .I1(n11_adj_4302), .I2(n2637), 
            .I3(n98), .O(n48259));
    defparam i32757_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i33087_4_lut (.I0(n19_adj_4309), .I1(n17_adj_4308), .I2(n15_adj_4306), 
            .I3(n48259), .O(n48589));
    defparam i33087_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33072_4_lut (.I0(n25_adj_4313), .I1(n23_adj_4312), .I2(n21_adj_4311), 
            .I3(n48589), .O(n48574));
    defparam i33072_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32040_4_lut (.I0(n31_adj_4316), .I1(n29_adj_4315), .I2(n27_adj_4314), 
            .I3(n48574), .O(n47541));
    defparam i32040_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1722_i8_4_lut (.I0(n389), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4300));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33429_3_lut (.I0(n8_adj_4300), .I1(n87), .I2(n31_adj_4316), 
            .I3(GND_net), .O(n48931));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33429_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33430_3_lut (.I0(n48931), .I1(n86), .I2(n33_adj_4317), .I3(GND_net), 
            .O(n48932));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33430_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1722_i34_3_lut (.I0(n16_adj_4307), .I1(n83), 
            .I2(n39_adj_4321), .I3(GND_net), .O(n34_adj_4318));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31998_4_lut (.I0(n37_adj_4320), .I1(n35_adj_4319), .I2(n33_adj_4317), 
            .I3(n47539), .O(n47498));
    defparam i31998_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33660_4_lut (.I0(n34_adj_4318), .I1(n14_adj_4305), .I2(n39_adj_4321), 
            .I3(n47494), .O(n49162));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33660_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33340_3_lut (.I0(n48932), .I1(n85), .I2(n35_adj_4319), .I3(GND_net), 
            .O(n48842));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33340_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33431_3_lut (.I0(n10_adj_4301), .I1(n90), .I2(n25_adj_4313), 
            .I3(GND_net), .O(n48933));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33431_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33432_3_lut (.I0(n48933), .I1(n89), .I2(n27_adj_4314), .I3(GND_net), 
            .O(n48934));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33432_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32698_4_lut (.I0(n27_adj_4314), .I1(n25_adj_4313), .I2(n23_adj_4312), 
            .I3(n47581), .O(n48200));
    defparam i32698_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_LessThan_1722_i20_3_lut (.I0(n12_adj_4303), .I1(n91), 
            .I2(n23_adj_4312), .I3(GND_net), .O(n20_adj_4310));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33338_3_lut (.I0(n48934), .I1(n88), .I2(n29_adj_4315), .I3(GND_net), 
            .O(n48840));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33338_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33277_4_lut (.I0(n37_adj_4320), .I1(n35_adj_4319), .I2(n33_adj_4317), 
            .I3(n47541), .O(n48779));
    defparam i33277_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33747_4_lut (.I0(n48842), .I1(n49162), .I2(n39_adj_4321), 
            .I3(n47498), .O(n49249));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33747_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33343_4_lut (.I0(n48840), .I1(n20_adj_4310), .I2(n29_adj_4315), 
            .I3(n48200), .O(n48845));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33343_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33765_4_lut (.I0(n48845), .I1(n49249), .I2(n39_adj_4321), 
            .I3(n48779), .O(n49267));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33765_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33766_3_lut (.I0(n49267), .I1(n82), .I2(n2621), .I3(GND_net), 
            .O(n49268));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33766_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33756_3_lut (.I0(n49268), .I1(n81), .I2(n2620), .I3(GND_net), 
            .O(n49258));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33756_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33345_3_lut (.I0(n49258), .I1(n80), .I2(n2619), .I3(GND_net), 
            .O(n48847));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33345_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1485 (.I0(n48847), .I1(n22561), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1485.LUT_INIT = 16'hceef;
    SB_LUT4 i1_2_lut_4_lut_adj_1486 (.I0(n96), .I1(n95), .I2(n94), .I3(n22516), 
            .O(n22507));
    defparam i1_2_lut_4_lut_adj_1486.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1487 (.I0(n95), .I1(n94), .I2(n22516), 
            .I3(GND_net), .O(n22510));
    defparam i1_2_lut_3_lut_adj_1487.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4297));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4299));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1488 (.I0(n93), .I1(n92), .I2(n91), .I3(n22525), 
            .O(n22516));
    defparam i1_2_lut_4_lut_adj_1488.LUT_INIT = 16'hff7f;
    SB_LUT4 div_12_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4295));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n388));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1489 (.I0(n92), .I1(n91), .I2(n22525), 
            .I3(GND_net), .O(n22519));
    defparam i1_2_lut_3_lut_adj_1489.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4298));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4292));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4293));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1490 (.I0(n90), .I1(n89), .I2(n88), .I3(n22534), 
            .O(n22525));
    defparam i1_2_lut_4_lut_adj_1490.LUT_INIT = 16'hff7f;
    SB_LUT4 div_12_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4289));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1263_3_lut_3_lut (.I0(n1886), .I1(n6829), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4290));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4291));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4121));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31946_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n47446));
    defparam i31946_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4123));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4280));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4282));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4284));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4286));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4287));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4294));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32138_4_lut (.I0(n33_adj_4294), .I1(n21_adj_4287), .I2(n19_adj_4286), 
            .I3(n17_adj_4284), .O(n47639));
    defparam i32138_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32815_4_lut (.I0(n15_adj_4282), .I1(n13_adj_4280), .I2(n2552), 
            .I3(n98), .O(n48317));
    defparam i32815_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i33111_4_lut (.I0(n21_adj_4287), .I1(n19_adj_4286), .I2(n17_adj_4284), 
            .I3(n48317), .O(n48613));
    defparam i33111_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33109_4_lut (.I0(n27_adj_4291), .I1(n25_adj_4290), .I2(n23_adj_4289), 
            .I3(n48613), .O(n48611));
    defparam i33109_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32146_4_lut (.I0(n33_adj_4294), .I1(n31_adj_4293), .I2(n29_adj_4292), 
            .I3(n48611), .O(n47647));
    defparam i32146_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1665_i10_4_lut (.I0(n388), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4278));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33191_3_lut (.I0(n10_adj_4278), .I1(n87), .I2(n33_adj_4294), 
            .I3(GND_net), .O(n48693));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33191_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33192_3_lut (.I0(n48693), .I1(n86), .I2(n35_adj_4295), .I3(GND_net), 
            .O(n48694));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33192_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1665_i36_3_lut (.I0(n18_adj_4285), .I1(n83), 
            .I2(n41_adj_4299), .I3(GND_net), .O(n36_adj_4296));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32130_4_lut (.I0(n39_adj_4298), .I1(n37_adj_4297), .I2(n35_adj_4295), 
            .I3(n47639), .O(n47631));
    defparam i32130_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33611_4_lut (.I0(n36_adj_4296), .I1(n16_adj_4283), .I2(n41_adj_4299), 
            .I3(n47628), .O(n49113));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33611_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32740_3_lut (.I0(n48694), .I1(n85), .I2(n37_adj_4297), .I3(GND_net), 
            .O(n48242));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32740_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i31934_4_lut (.I0(n33_adj_4135), .I1(n31_adj_4134), .I2(n29_adj_4132), 
            .I3(n27), .O(n47434));
    defparam i31934_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1665_i22_3_lut (.I0(n14_adj_4281), .I1(n91), 
            .I2(n25_adj_4290), .I3(GND_net), .O(n22_adj_4288));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33609_4_lut (.I0(n22_adj_4288), .I1(n12_adj_4279), .I2(n25_adj_4290), 
            .I3(n47690), .O(n49111));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33609_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33610_3_lut (.I0(n49111), .I1(n90), .I2(n27_adj_4291), .I3(GND_net), 
            .O(n49112));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33610_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33470_3_lut (.I0(n49112), .I1(n89), .I2(n29_adj_4292), .I3(GND_net), 
            .O(n48972));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33470_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33373_4_lut (.I0(n39_adj_4298), .I1(n37_adj_4297), .I2(n35_adj_4295), 
            .I3(n47647), .O(n48875));
    defparam i33373_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33727_4_lut (.I0(n48242), .I1(n49113), .I2(n41_adj_4299), 
            .I3(n47631), .O(n49229));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33727_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32738_3_lut (.I0(n48972), .I1(n88), .I2(n31_adj_4293), .I3(GND_net), 
            .O(n48240));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32738_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33761_4_lut (.I0(n48240), .I1(n49229), .I2(n41_adj_4299), 
            .I3(n48875), .O(n49263));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33761_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33762_3_lut (.I0(n49263), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n49264));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33762_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i33760_3_lut (.I0(n49264), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n49262));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33760_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_12_i1262_3_lut_3_lut (.I0(n1886), .I1(n6828), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1491 (.I0(n49262), .I1(n22558), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1491.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4275));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4273));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4277));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4276));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n387_adj_4000));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4270));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4271));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1492 (.I0(n88), .I1(n87), .I2(n22537), 
            .I3(GND_net), .O(n22531));
    defparam i1_2_lut_3_lut_adj_1492.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4267));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4268));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4269));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i23120_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n372), .I3(n558), 
            .O(n4_adj_4045));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23120_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_12_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4258));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4260));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4262));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4264));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4265));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4272));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32241_4_lut (.I0(n35_adj_4272), .I1(n23_adj_4265), .I2(n21_adj_4264), 
            .I3(n19_adj_4262), .O(n47743));
    defparam i32241_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32863_4_lut (.I0(n17_adj_4260), .I1(n15_adj_4258), .I2(n2464), 
            .I3(n98), .O(n48365));
    defparam i32863_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i33131_4_lut (.I0(n23_adj_4265), .I1(n21_adj_4264), .I2(n19_adj_4262), 
            .I3(n48365), .O(n48633));
    defparam i33131_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33127_4_lut (.I0(n29_adj_4269), .I1(n27_adj_4268), .I2(n25_adj_4267), 
            .I3(n48633), .O(n48629));
    defparam i33127_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32245_4_lut (.I0(n35_adj_4272), .I1(n33_adj_4271), .I2(n31_adj_4270), 
            .I3(n48629), .O(n47747));
    defparam i32245_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_i1261_3_lut_3_lut (.I0(n1886), .I1(n6827), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1260_3_lut_3_lut (.I0(n1886), .I1(n6826), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1259_3_lut_3_lut (.I0(n1886), .I1(n6825), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1606_i12_4_lut (.I0(n387_adj_4000), .I1(n99), 
            .I2(n2465), .I3(n558), .O(n12_adj_4256));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33197_3_lut (.I0(n12_adj_4256), .I1(n87), .I2(n35_adj_4272), 
            .I3(GND_net), .O(n48699));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33197_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1606_i38_3_lut (.I0(n20_adj_4263), .I1(n83), 
            .I2(n43_adj_4277), .I3(GND_net), .O(n38_adj_4274));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33198_3_lut (.I0(n48699), .I1(n86), .I2(n37_adj_4273), .I3(GND_net), 
            .O(n48700));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33198_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32220_4_lut (.I0(n41_adj_4276), .I1(n39_adj_4275), .I2(n37_adj_4273), 
            .I3(n47743), .O(n47722));
    defparam i32220_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33585_4_lut (.I0(n38_adj_4274), .I1(n18_adj_4261), .I2(n43_adj_4277), 
            .I3(n47718), .O(n49087));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33585_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32734_3_lut (.I0(n48700), .I1(n85), .I2(n39_adj_4275), .I3(GND_net), 
            .O(n48236));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32734_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1258_3_lut_3_lut (.I0(n1886), .I1(n6824), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1606_i24_3_lut (.I0(n16_adj_4259), .I1(n91), 
            .I2(n27_adj_4268), .I3(GND_net), .O(n24_adj_4266));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1266_3_lut_3_lut (.I0(n1886), .I1(n6832), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33617_4_lut (.I0(n24_adj_4266), .I1(n14_adj_4257), .I2(n27_adj_4268), 
            .I3(n47755), .O(n49119));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33617_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33618_3_lut (.I0(n49119), .I1(n90), .I2(n29_adj_4269), .I3(GND_net), 
            .O(n49120));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33618_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33472_3_lut (.I0(n49120), .I1(n89), .I2(n31_adj_4270), .I3(GND_net), 
            .O(n48974));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33472_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33385_4_lut (.I0(n41_adj_4276), .I1(n39_adj_4275), .I2(n37_adj_4273), 
            .I3(n47747), .O(n48887));
    defparam i33385_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33715_4_lut (.I0(n48236), .I1(n49087), .I2(n43_adj_4277), 
            .I3(n47722), .O(n49217));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33715_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32732_3_lut (.I0(n48974), .I1(n88), .I2(n33_adj_4271), .I3(GND_net), 
            .O(n48234));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32732_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33753_4_lut (.I0(n48234), .I1(n49217), .I2(n43_adj_4277), 
            .I3(n48887), .O(n49255));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33753_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33754_3_lut (.I0(n49255), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n49256));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33754_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1493 (.I0(n49256), .I1(n22555), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1493.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1340_3_lut_3_lut (.I0(n1991), .I1(n6853), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n22561));
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_i1331_3_lut_3_lut (.I0(n1991), .I1(n6844), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_12_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1495 (.I0(n81), .I1(n22555), .I2(GND_net), .I3(GND_net), 
            .O(n22552));
    defparam i1_2_lut_adj_1495.LUT_INIT = 16'hdddd;
    SB_LUT4 div_12_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4253));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4255));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4251));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n386));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_i1330_3_lut_3_lut (.I0(n1991), .I1(n6843), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4254));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1329_3_lut_3_lut (.I0(n1991), .I1(n6842), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4248));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4249));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4143));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1328_3_lut_3_lut (.I0(n1991), .I1(n6841), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4245));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4246));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4247));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31886_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n47386));
    defparam i31886_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4145));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4236));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4238));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31896_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n47396));
    defparam i31896_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_4147));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4240));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4242));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4243));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4250));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32279_4_lut (.I0(n37_adj_4250), .I1(n25_adj_4243), .I2(n23_adj_4242), 
            .I3(n21_adj_4240), .O(n47781));
    defparam i32279_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32899_4_lut (.I0(n19_adj_4238), .I1(n17_adj_4236), .I2(n2373), 
            .I3(n98), .O(n48401));
    defparam i32899_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i33151_4_lut (.I0(n25_adj_4243), .I1(n23_adj_4242), .I2(n21_adj_4240), 
            .I3(n48401), .O(n48653));
    defparam i33151_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33147_4_lut (.I0(n31_adj_4247), .I1(n29_adj_4246), .I2(n27_adj_4245), 
            .I3(n48653), .O(n48649));
    defparam i33147_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32281_4_lut (.I0(n37_adj_4250), .I1(n35_adj_4249), .I2(n33_adj_4248), 
            .I3(n48649), .O(n47783));
    defparam i32281_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_12_LessThan_1545_i14_4_lut (.I0(n386), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4234));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33201_3_lut (.I0(n14_adj_4234), .I1(n87), .I2(n37_adj_4250), 
            .I3(GND_net), .O(n48703));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33201_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33202_3_lut (.I0(n48703), .I1(n86), .I2(n39_adj_4251), .I3(GND_net), 
            .O(n48704));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33202_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1545_i40_3_lut (.I0(n22_adj_4241), .I1(n83), 
            .I2(n45_adj_4255), .I3(GND_net), .O(n40_adj_4252));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32273_4_lut (.I0(n43_adj_4254), .I1(n41_adj_4253), .I2(n39_adj_4251), 
            .I3(n47781), .O(n47775));
    defparam i32273_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33333_4_lut (.I0(n40_adj_4252), .I1(n20_adj_4239), .I2(n45_adj_4255), 
            .I3(n47773), .O(n48835));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33333_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32726_3_lut (.I0(n48704), .I1(n85), .I2(n41_adj_4253), .I3(GND_net), 
            .O(n48228));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32726_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1545_i26_3_lut (.I0(n18_adj_4237), .I1(n91), 
            .I2(n29_adj_4246), .I3(GND_net), .O(n26_adj_4244));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33607_4_lut (.I0(n26_adj_4244), .I1(n16_adj_4235), .I2(n29_adj_4246), 
            .I3(n47795), .O(n49109));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33607_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33608_3_lut (.I0(n49109), .I1(n90), .I2(n31_adj_4247), .I3(GND_net), 
            .O(n49110));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33608_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33474_3_lut (.I0(n49110), .I1(n89), .I2(n33_adj_4248), .I3(GND_net), 
            .O(n48976));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33474_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33393_4_lut (.I0(n43_adj_4254), .I1(n41_adj_4253), .I2(n39_adj_4251), 
            .I3(n47783), .O(n48895));
    defparam i33393_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33633_4_lut (.I0(n48228), .I1(n48835), .I2(n45_adj_4255), 
            .I3(n47775), .O(n49135));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33633_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32724_3_lut (.I0(n48976), .I1(n88), .I2(n35_adj_4249), .I3(GND_net), 
            .O(n48226));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32724_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33635_4_lut (.I0(n48226), .I1(n49135), .I2(n45_adj_4255), 
            .I3(n48895), .O(n49137));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33635_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1496 (.I0(n49137), .I1(n22552), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1496.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4230));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4233));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4232));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4231));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n385));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4227));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4228));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4229));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4224));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4226));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4223));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4218));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4220));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4222));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4216));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31758_4_lut (.I0(n23_adj_4222), .I1(n21_adj_4220), .I2(n19_adj_4218), 
            .I3(n17_adj_4216), .O(n47258));
    defparam i31758_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32338_4_lut (.I0(n29_adj_4226), .I1(n27_adj_4224), .I2(n25_adj_4223), 
            .I3(n47258), .O(n47840));
    defparam i32338_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33403_4_lut (.I0(n35_adj_4229), .I1(n33_adj_4228), .I2(n31_adj_4227), 
            .I3(n47840), .O(n48905));
    defparam i33403_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_12_LessThan_1482_i16_4_lut (.I0(n385), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4215));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33207_3_lut (.I0(n16_adj_4215), .I1(n87), .I2(n39_adj_4231), 
            .I3(GND_net), .O(n48709));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33207_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33208_3_lut (.I0(n48709), .I1(n86), .I2(n41_adj_4232), .I3(GND_net), 
            .O(n48710));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33208_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32909_4_lut (.I0(n41_adj_4232), .I1(n39_adj_4231), .I2(n27_adj_4224), 
            .I3(n47252), .O(n48411));
    defparam i32909_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33331_3_lut (.I0(n22_adj_4221), .I1(n93), .I2(n27_adj_4224), 
            .I3(GND_net), .O(n48833));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33331_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32716_3_lut (.I0(n48710), .I1(n85), .I2(n43_adj_4233), .I3(GND_net), 
            .O(n48218));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32716_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_LessThan_1482_i28_3_lut (.I0(n20_adj_4219), .I1(n91), 
            .I2(n31_adj_4227), .I3(GND_net), .O(n28_adj_4225));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1327_3_lut_3_lut (.I0(n1991), .I1(n6840), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33605_4_lut (.I0(n28_adj_4225), .I1(n18_adj_4217), .I2(n31_adj_4227), 
            .I3(n47838), .O(n49107));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33605_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33606_3_lut (.I0(n49107), .I1(n90), .I2(n33_adj_4228), .I3(GND_net), 
            .O(n49108));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33606_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33478_3_lut (.I0(n49108), .I1(n89), .I2(n35_adj_4229), .I3(GND_net), 
            .O(n48980));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33478_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1339_3_lut_3_lut (.I0(n1991), .I1(n6852), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i32913_4_lut (.I0(n41_adj_4232), .I1(n39_adj_4231), .I2(n37_adj_4230), 
            .I3(n48905), .O(n48415));
    defparam i32913_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i33475_4_lut (.I0(n48218), .I1(n48833), .I2(n43_adj_4233), 
            .I3(n48411), .O(n48977));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33475_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32714_3_lut (.I0(n48980), .I1(n88), .I2(n37_adj_4230), .I3(GND_net), 
            .O(n48216));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i32714_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33670_4_lut (.I0(n48216), .I1(n48977), .I2(n43_adj_4233), 
            .I3(n48415), .O(n49172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33670_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33671_3_lut (.I0(n49172), .I1(n84), .I2(n2265_adj_4010), 
            .I3(GND_net), .O(n49173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33671_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1497 (.I0(n49173), .I1(n22549), .I2(n83), .I3(n2264_adj_4009), 
            .O(n2288));
    defparam i1_4_lut_adj_1497.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4112));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4210));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31971_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n47471));
    defparam i31971_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4214));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4113));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4213));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i23088_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n371), .I3(n558), 
            .O(n4));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i23088_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_12_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4211));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1498 (.I0(n86), .I1(n85), .I2(n84), .I3(n22546), 
            .O(n22537));
    defparam i1_2_lut_4_lut_adj_1498.LUT_INIT = 16'hff7f;
    SB_LUT4 div_12_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n384));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_12_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4131));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4207));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4208));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4209));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31925_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n47425));
    defparam i31925_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4204));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4206));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4197));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4199));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n22467), 
            .O(n249));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 div_12_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4201));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4203));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4195));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31790_4_lut (.I0(n25_adj_4201), .I1(n23_adj_4199), .I2(n21_adj_4197), 
            .I3(n19_adj_4195), .O(n47290));
    defparam i31790_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31784_4_lut (.I0(n31_adj_4206), .I1(n29_adj_4204), .I2(n27_adj_4203), 
            .I3(n47290), .O(n47284));
    defparam i31784_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33213_4_lut (.I0(n37_adj_4209), .I1(n35_adj_4208), .I2(n33_adj_4207), 
            .I3(n47284), .O(n48715));
    defparam i33213_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_12_LessThan_1417_i18_4_lut (.I0(n384), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4194));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i33433_3_lut (.I0(n18_adj_4194), .I1(n87), .I2(n41_adj_4211), 
            .I3(GND_net), .O(n48935));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33433_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33434_3_lut (.I0(n48935), .I1(n86), .I2(n43_adj_4213), .I3(GND_net), 
            .O(n48936));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33434_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32466_4_lut (.I0(n43_adj_4213), .I1(n41_adj_4211), .I2(n29_adj_4204), 
            .I3(n47288), .O(n47968));
    defparam i32466_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_LessThan_1417_i26_3_lut (.I0(n24_adj_4200), .I1(n93), 
            .I2(n29_adj_4204), .I3(GND_net), .O(n26_adj_4202));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33330_3_lut (.I0(n48936), .I1(n85), .I2(n45_adj_4214), .I3(GND_net), 
            .O(n42_adj_4212));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33330_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1404_3_lut_3_lut (.I0(n2093), .I1(n6867), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1417_i30_3_lut (.I0(n22_adj_4198), .I1(n91), 
            .I2(n33_adj_4207), .I3(GND_net), .O(n30_adj_4205));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33658_4_lut (.I0(n30_adj_4205), .I1(n20_adj_4196), .I2(n33_adj_4207), 
            .I3(n47282), .O(n49160));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33658_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_12_i1399_3_lut_3_lut (.I0(n2093), .I1(n6862), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1409_3_lut_3_lut (.I0(n2093), .I1(n6872), .I2(n383), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33659_3_lut (.I0(n49160), .I1(n90), .I2(n35_adj_4208), .I3(GND_net), 
            .O(n49161));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33659_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_12_i1397_3_lut_3_lut (.I0(n2093), .I1(n6860), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1396_3_lut_3_lut (.I0(n2093), .I1(n6859), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33588_3_lut (.I0(n49161), .I1(n89), .I2(n37_adj_4209), .I3(GND_net), 
            .O(n49090));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33588_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i32470_4_lut (.I0(n43_adj_4213), .I1(n41_adj_4211), .I2(n39_adj_4210), 
            .I3(n48715), .O(n47972));
    defparam i32470_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_12_i1395_3_lut_3_lut (.I0(n2093), .I1(n6858), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33084_4_lut (.I0(n42_adj_4212), .I1(n26_adj_4202), .I2(n45_adj_4214), 
            .I3(n47968), .O(n48586));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33084_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33532_3_lut (.I0(n49090), .I1(n88), .I2(n39_adj_4210), .I3(GND_net), 
            .O(n49034));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33532_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33086_4_lut (.I0(n49034), .I1(n48586), .I2(n45_adj_4214), 
            .I3(n47972), .O(n48588));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam i33086_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1499 (.I0(n48588), .I1(n22546), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1499.LUT_INIT = 16'hceef;
    SB_LUT4 div_12_i1398_3_lut_3_lut (.I0(n2093), .I1(n6861), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1394_3_lut_3_lut (.I0(n2093), .I1(n6857), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1405_3_lut_3_lut (.I0(n2093), .I1(n6868), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1408_3_lut_3_lut (.I0(n2093), .I1(n6871), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1406_3_lut_3_lut (.I0(n2093), .I1(n6869), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1337_3_lut_3_lut (.I0(n1991), .I1(n6850), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1407_3_lut_3_lut (.I0(n2093), .I1(n6870), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1403_3_lut_3_lut (.I0(n2093), .I1(n6866), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1402_3_lut_3_lut (.I0(n2093), .I1(n6865), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1400_3_lut_3_lut (.I0(n2093), .I1(n6863), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1401_3_lut_3_lut (.I0(n2093), .I1(n6864), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_i1459_3_lut_3_lut (.I0(n2192), .I1(n6875), .I2(n2168), 
            .I3(GND_net), .O(n2264_adj_4009));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4133));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_adj_1500 (.I0(n85), .I1(n84), .I2(n22546), 
            .I3(GND_net), .O(n22540));
    defparam i1_2_lut_3_lut_adj_1500.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1501 (.I0(n83), .I1(n82), .I2(n81), .I3(n22555), 
            .O(n22546));
    defparam i1_2_lut_4_lut_adj_1501.LUT_INIT = 16'hff7f;
    SB_LUT4 div_12_i1460_3_lut_3_lut (.I0(n2192), .I1(n6876), .I2(n2169), 
            .I3(GND_net), .O(n2265_adj_4010));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4161));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1474_3_lut_3_lut (.I0(n2192), .I1(n6890), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31849_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n47349));
    defparam i31849_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4193));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4163));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1466_3_lut_3_lut (.I0(n2192), .I1(n6882), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_12_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4192));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1467_3_lut_3_lut (.I0(n2192), .I1(n6883), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31855_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n47355));
    defparam i31855_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4190));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_4165));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4191));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_i1465_3_lut_3_lut (.I0(n2192), .I1(n6881), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    coms c0 (.clk32MHz(clk32MHz), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .GND_net(GND_net), 
         .gearBoxRatio({gearBoxRatio}), .n10(n10_adj_4035), .n24253(n24253), 
         .\data_in[0] ({Open_0, \data_in[0] [6:1], Open_1}), .n24252(n24252), 
         .n24251(n24251), .\data_in_frame[14] ({Open_2, Open_3, Open_4, 
         \data_in_frame[14] [4], Open_5, Open_6, Open_7, Open_8}), 
         .\data_in_frame[19] ({\data_in_frame[19] }), .n24250(n24250), .rx_data({rx_data}), 
         .\deadband[9] (deadband[9]), .\deadband[8] (deadband[8]), .\deadband[7] (deadband[7]), 
         .\deadband[6] (deadband[6]), .\deadband[5] (deadband[5]), .\deadband[4] (deadband[4]), 
         .\deadband[3] (deadband[3]), .\deadband[2] (deadband[2]), .\deadband[1] (deadband[1]), 
         .n24412(n24412), .setpoint({setpoint}), .n24411(n24411), .n24410(n24410), 
         .n42279(n42279), .n24408(n24408), .n24407(n24407), .n24406(n24406), 
         .n24405(n24405), .n24404(n24404), .n24403(n24403), .n24402(n24402), 
         .n24401(n24401), .n24400(n24400), .n24399(n24399), .n24398(n24398), 
         .n24397(n24397), .n24396(n24396), .n24395(n24395), .n24394(n24394), 
         .n24393(n24393), .n24392(n24392), .n24391(n24391), .n24390(n24390), 
         .n24388(n24388), .VCC_net(VCC_net), .byte_transmit_counter({Open_9, 
         Open_10, Open_11, Open_12, Open_13, Open_14, Open_15, byte_transmit_counter[0]}), 
         .n23822(n23822), .n24236(n24236), .\data_in[2] ({Open_16, \data_in[2] [6:2], 
         Open_17, Open_18}), .n24234(n24234), .n24233(n24233), .n24228(n24228), 
         .\data_in[3][2] (\data_in[3] [2]), .n24227(n24227), .\data_in[3][3] (\data_in[3] [3]), 
         .n24226(n24226), .\data_in[3][4] (\data_in[3] [4]), .n24225(n24225), 
         .\data_in[3][5] (\data_in[3] [5]), .n24223(n24223), .\data_in[3][7] (\data_in[3] [7]), 
         .n24222(n24222), .\data_out_frame[0][2] (\data_out_frame[0] [2]), 
         .n24221(n24221), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n24220(n24220), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .n24217(n24217), .\data_out_frame[5][2] (\data_out_frame[5] [2]), 
         .IntegralLimit({IntegralLimit}), .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), 
         .n24249(n24249), .n24248(n24248), .rx_data_ready(rx_data_ready), 
         .n24245(n24245), .\data_in[1][1] (\data_in[1] [1]), .n24244(n24244), 
         .\data_in[1][2] (\data_in[1] [2]), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), 
         .\FRAME_MATCHER.state ({Open_19, Open_20, Open_21, Open_22, 
         Open_23, Open_24, Open_25, Open_26, Open_27, Open_28, Open_29, 
         Open_30, Open_31, Open_32, Open_33, Open_34, Open_35, Open_36, 
         Open_37, Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, 
         Open_44, Open_45, Open_46, \FRAME_MATCHER.state [3:0]}), .n47(n47), 
         .n3839(n3839), .n29726(n29726), .\Kp[5] (Kp[5]), .n43231(n43231), 
         .n43238(n43238), .n43253(n43253), .\data_in_frame[1][4] (\data_in_frame[1] [4]), 
         .n24068(n24068), .\data_in_frame[3] ({\data_in_frame[3] }), .n24067(n24067), 
         .n24066(n24066), .n24065(n24065), .n24064(n24064), .n24063(n24063), 
         .n24062(n24062), .n24061(n24061), .n24243(n24243), .\data_in[1][3] (\data_in[1] [3]), 
         .\data_in_frame[5] ({\data_in_frame[5] }), .n24052(n24052), .n24051(n24051), 
         .n24050(n24050), .n24049(n24049), .n23533(n23533), .n24048(n24048), 
         .n24047(n24047), .n24046(n24046), .n24045(n24045), .\Kp[6] (Kp[6]), 
         .\Kp[7] (Kp[7]), .\Ki[1] (Ki[1]), .n24036(n24036), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .n24035(n24035), .n24034(n24034), .n24033(n24033), .n24032(n24032), 
         .n24031(n24031), .n24030(n24030), .n24029(n24029), .n24242(n24242), 
         .\data_in[1][4] (\data_in[1] [4]), .n23825(n23825), .\data_in_frame[10][6] (\data_in_frame[10] [6]), 
         .n24004(n24004), .n24003(n24003), .n24002(n24002), .n24001(n24001), 
         .n24000(n24000), .n23999(n23999), .n23998(n23998), .n23997(n23997), 
         .n23988(n23988), .n23987(n23987), .n23986(n23986), .n23985(n23985), 
         .n23984(n23984), .n23983(n23983), .n23982(n23982), .n20342(n20342), 
         .n23981(n23981), .\data_in_frame[14][0] (\data_in_frame[14] [0]), 
         .n24241(n24241), .\data_in[1][5] (\data_in[1] [5]), .n23972(n23972), 
         .\data_in_frame[15] ({\data_in_frame[15] }), .n23971(n23971), .n23970(n23970), 
         .n23969(n23969), .n23968(n23968), .n23967(n23967), .n23966(n23966), 
         .n23965(n23965), .n23838(n23838), .n22456(n22456), .n43255(n43255), 
         .\data_in_frame[16][1] (\data_in_frame[16] [1]), .n23835(n23835), 
         .n23832(n23832), .n23823(n23823), .n23820(n23820), .n2241(n2241), 
         .\data_in_frame[18][0] (\data_in_frame[18] [0]), .\data_in_frame[18][2] (\data_in_frame[18] [2]), 
         .Kp_23__N_865(Kp_23__N_865), .n43441(n43441), .n23940(n23940), 
         .n23939(n23939), .n23938(n23938), .n103(n103), .n23937(n23937), 
         .n23936(n23936), .n23935(n23935), .n23934(n23934), .n23933(n23933), 
         .Kp_23__N_515(Kp_23__N_515), .n45225(n45225), .n122(n122), .n44586(n44586), 
         .n23924(n23924), .\data_in_frame[21] ({\data_in_frame[21] }), .n23923(n23923), 
         .n23922(n23922), .n23921(n23921), .n23920(n23920), .n23919(n23919), 
         .n23918(n23918), .n23917(n23917), .control_mode({control_mode}), 
         .\PWMLimit[1] (PWMLimit[1]), .\PWMLimit[2] (PWMLimit[2]), .\PWMLimit[3] (PWMLimit[3]), 
         .\PWMLimit[4] (PWMLimit[4]), .\PWMLimit[5] (PWMLimit[5]), .\PWMLimit[6] (PWMLimit[6]), 
         .\PWMLimit[7] (PWMLimit[7]), .\PWMLimit[8] (PWMLimit[8]), .\PWMLimit[9] (PWMLimit[9]), 
         .n50101(n50101), .n23834(n23834), .n23837(n23837), .n23840(n23840), 
         .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .n24240(n24240), 
         .\data_in[1][6] (\data_in[1] [6]), .\Ki[5] (Ki[5]), .\data_in[2][1] (\data_in[2] [1]), 
         .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .\Kd[1] (Kd[1]), .\Kd[2] (Kd[2]), 
         .\Kd[3] (Kd[3]), .n43459(n43459), .\Kd[4] (Kd[4]), .\Kd[5] (Kd[5]), 
         .\Kd[6] (Kd[6]), .\Kd[7] (Kd[7]), .\deadband[0] (deadband[0]), 
         .n23756(n23756), .n42561(n42561), .\PWMLimit[0] (PWMLimit[0]), 
         .\Kd[0] (Kd[0]), .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .n22(n22_adj_4027), 
         .n22833(n22833), .n40155(n40155), .n44311(n44311), .n43709(n43709), 
         .n3799(n3799), .n3800(n3800), .n3801(n3801), .n3802(n3802), 
         .n3803(n3803), .n3804(n3804), .n3805(n3805), .n22429(n22429), 
         .encoder0_position({encoder0_position}), .n3806(n3806), .n3807(n3807), 
         .displacement({displacement}), .n3808(n3808), .encoder1_position({encoder1_position}), 
         .n3809(n3809), .n3810(n3810), .n3811(n3811), .n3812(n3812), 
         .n3813(n3813), .pwm({pwm}), .n3814(n3814), .n44238(n44238), 
         .n3815(n3815), .n5022(n5022), .n23563(n23563), .n3817(n3817), 
         .n3818(n3818), .n3822(n3822), .n3816(n3816), .n3820(n3820), 
         .n3821(n3821), .n7(n7_adj_4012), .n5(n5_adj_4011), .n5_adj_3(n5_adj_4375), 
         .n44019(n44019), .n22458(n22458), .n20136(n20136), .n44009(n44009), 
         .n43229(n43229), .n43236(n43236), .n43251(n43251), .n23776(n23776), 
         .n23779(n23779), .n23778(n23778), .n23781(n23781), .n23784(n23784), 
         .n23787(n23787), .n23790(n23790), .n23793(n23793), .n23796(n23796), 
         .n23799(n23799), .n23803(n23803), .r_Bit_Index({r_Bit_Index_adj_4419}), 
         .n23806(n23806), .n23782(n23782), .n23785(n23785), .n23788(n23788), 
         .n23602(n23602), .n23716(n23716), .n4037(n4037), .n23845(n23845), 
         .n23791(n23791), .n23794(n23794), .n23797(n23797), .n23844(n23844), 
         .n23846(n23846), .n23849(n23849), .tx_o(tx_o), .tx_enable(tx_enable), 
         .n23809(n23809), .r_Bit_Index_adj_9({r_Bit_Index}), .n23812(n23812), 
         .n28794(n28794), .\r_SM_Main[1] (r_SM_Main[1]), .n24357(n24357), 
         .r_Rx_Data(r_Rx_Data), .LED_c(LED_c), .\r_SM_Main[2] (r_SM_Main[2]), 
         .n23596(n23596), .n23714(n23714), .n4015(n4015), .n23819(n23819), 
         .n23818(n23818), .n23817(n23817), .n23816(n23816), .n23853(n23853), 
         .n23815(n23815), .n23814(n23814), .n23813(n23813), .n23751(n23751), 
         .n28760(n28760), .n1(n1_adj_4372), .n28350(n28350), .n4(n4_adj_3993), 
         .n4_adj_7(n4_adj_3987), .n22470(n22470), .n22462(n22462), .n4_adj_8(n4_adj_3986), 
         .n47207(n47207), .n47206(n47206)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(79[8] 98[4])
    SB_LUT4 div_12_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n383));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1502 (.I0(n82), .I1(n81), .I2(n22555), 
            .I3(GND_net), .O(n22549));
    defparam i1_2_lut_3_lut_adj_1502.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_12_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4179));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i31810_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n47310));
    defparam i31810_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4186));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4187));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4189));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4181));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1475_3_lut_3_lut (.I0(n2192), .I1(n6891), .I2(n384), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i31816_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n47316));
    defparam i31816_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_12_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4180));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4182));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4184));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_12_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_4183));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_12_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_12_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4178));   // verilog/TinyFPGA_B.v(162[21:53])
    defparam div_12_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i31820_4_lut (.I0(n27_adj_4184), .I1(n25_adj_4182), .I2(n23_adj_4180), 
            .I3(n21_adj_4178), .O(n47320));
    defparam i31820_4_lut.LUT_INIT = 16'haaab;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n2291, encoder0_position, GND_net, 
            data_o, clk32MHz, n23875, n23874, n23873, n23872, n23871, 
            n23870, n23869, n23868, n23867, n23866, n23865, n23864, 
            n23863, n23862, n23861, n23860, n23859, n23858, n23857, 
            n23856, n23855, n23854, n23850, n23745, count_enable, 
            n24359, reg_B, PIN_23_c_1, PIN_24_c_0, n23750, n44902) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]n2291;
    output [23:0]encoder0_position;
    input GND_net;
    output [1:0]data_o;
    input clk32MHz;
    input n23875;
    input n23874;
    input n23873;
    input n23872;
    input n23871;
    input n23870;
    input n23869;
    input n23868;
    input n23867;
    input n23866;
    input n23865;
    input n23864;
    input n23863;
    input n23862;
    input n23861;
    input n23860;
    input n23859;
    input n23858;
    input n23857;
    input n23856;
    input n23855;
    input n23854;
    input n23850;
    input n23745;
    output count_enable;
    input n24359;
    output [1:0]reg_B;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n23750;
    output n44902;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n2287, n36987, n36988, n36986, n36985, n36984, count_direction, 
        n36983, B_delayed, A_delayed, n37006, n37005, n37004, n37003, 
        n37002, n37001, n37000, n36999, n36998, n36997, n36996, 
        n36995, n36994, n36993, n36992, n36991, n36989, n36990;
    
    SB_LUT4 add_549_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2287), 
            .I3(n36987), .O(n2291[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_6 (.CI(n36987), .I0(encoder0_position[4]), .I1(n2287), 
            .CO(n36988));
    SB_LUT4 add_549_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2287), 
            .I3(n36986), .O(n2291[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_5 (.CI(n36986), .I0(encoder0_position[3]), .I1(n2287), 
            .CO(n36987));
    SB_LUT4 add_549_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2287), 
            .I3(n36985), .O(n2291[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_4 (.CI(n36985), .I0(encoder0_position[2]), .I1(n2287), 
            .CO(n36986));
    SB_LUT4 add_549_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2287), 
            .I3(n36984), .O(n2291[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_3 (.CI(n36984), .I0(encoder0_position[1]), .I1(n2287), 
            .CO(n36985));
    SB_LUT4 add_549_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n36983), .O(n2291[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_2 (.CI(n36983), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n36984));
    SB_CARRY add_549_1 (.CI(GND_net), .I0(n2287), .I1(n2287), .CO(n36983));
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_549_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2287), 
            .I3(n37006), .O(n2291[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_549_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2287), 
            .I3(n37005), .O(n2291[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_24 (.CI(n37005), .I0(encoder0_position[22]), .I1(n2287), 
            .CO(n37006));
    SB_LUT4 add_549_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2287), 
            .I3(n37004), .O(n2291[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_23 (.CI(n37004), .I0(encoder0_position[21]), .I1(n2287), 
            .CO(n37005));
    SB_LUT4 add_549_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2287), 
            .I3(n37003), .O(n2291[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_22 (.CI(n37003), .I0(encoder0_position[20]), .I1(n2287), 
            .CO(n37004));
    SB_LUT4 add_549_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2287), 
            .I3(n37002), .O(n2291[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_21 (.CI(n37002), .I0(encoder0_position[19]), .I1(n2287), 
            .CO(n37003));
    SB_LUT4 add_549_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2287), 
            .I3(n37001), .O(n2291[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_20 (.CI(n37001), .I0(encoder0_position[18]), .I1(n2287), 
            .CO(n37002));
    SB_LUT4 add_549_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2287), 
            .I3(n37000), .O(n2291[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_19 (.CI(n37000), .I0(encoder0_position[17]), .I1(n2287), 
            .CO(n37001));
    SB_LUT4 add_549_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2287), 
            .I3(n36999), .O(n2291[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_18 (.CI(n36999), .I0(encoder0_position[16]), .I1(n2287), 
            .CO(n37000));
    SB_LUT4 add_549_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2287), 
            .I3(n36998), .O(n2291[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_17 (.CI(n36998), .I0(encoder0_position[15]), .I1(n2287), 
            .CO(n36999));
    SB_LUT4 add_549_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2287), 
            .I3(n36997), .O(n2291[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_16 (.CI(n36997), .I0(encoder0_position[14]), .I1(n2287), 
            .CO(n36998));
    SB_LUT4 add_549_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2287), 
            .I3(n36996), .O(n2291[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_15 (.CI(n36996), .I0(encoder0_position[13]), .I1(n2287), 
            .CO(n36997));
    SB_LUT4 add_549_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2287), 
            .I3(n36995), .O(n2291[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_14 (.CI(n36995), .I0(encoder0_position[12]), .I1(n2287), 
            .CO(n36996));
    SB_LUT4 add_549_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2287), 
            .I3(n36994), .O(n2291[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_13 (.CI(n36994), .I0(encoder0_position[11]), .I1(n2287), 
            .CO(n36995));
    SB_LUT4 add_549_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2287), 
            .I3(n36993), .O(n2291[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_12 (.CI(n36993), .I0(encoder0_position[10]), .I1(n2287), 
            .CO(n36994));
    SB_LUT4 add_549_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2287), 
            .I3(n36992), .O(n2291[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_11 (.CI(n36992), .I0(encoder0_position[9]), .I1(n2287), 
            .CO(n36993));
    SB_LUT4 add_549_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2287), 
            .I3(n36991), .O(n2291[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_10 (.CI(n36991), .I0(encoder0_position[8]), .I1(n2287), 
            .CO(n36992));
    SB_LUT4 add_549_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2287), 
            .I3(n36988), .O(n2291[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_8 (.CI(n36989), .I0(encoder0_position[6]), .I1(n2287), 
            .CO(n36990));
    SB_LUT4 add_549_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2287), 
            .I3(n36989), .O(n2291[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_9 (.CI(n36990), .I0(encoder0_position[7]), .I1(n2287), 
            .CO(n36991));
    SB_LUT4 add_549_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2287), 
            .I3(n36990), .O(n2291[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_549_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_549_7 (.CI(n36988), .I0(encoder0_position[5]), .I1(n2287), 
            .CO(n36989));
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n23875));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n23874));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n23873));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n23872));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n23871));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n23870));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n23869));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n23868));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n23867));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n23866));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n23865));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n23864));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n23863));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n23862));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n23861));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n23860));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n23859));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n23858));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n23857));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n23856));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n23855));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n23854));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n23850));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n23745));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i774_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2287));   // quad.v(37[5] 40[8])
    defparam i774_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n24359(n24359), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .PIN_23_c_1(PIN_23_c_1), 
            .PIN_24_c_0(PIN_24_c_0), .n23750(n23750), .GND_net(GND_net), 
            .n44902(n44902)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n24359, data_o, clk32MHz, reg_B, PIN_23_c_1, 
            PIN_24_c_0, n23750, GND_net, n44902) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24359;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input PIN_23_c_1;
    input PIN_24_c_0;
    input n23750;
    input GND_net;
    output n44902;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3104, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24359));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_23_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1049__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_24_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1049__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1049__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23750));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i23349_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23349_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i23342_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n44902));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n44902), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i23340_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23340_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \PWMLimit[4] , \PWMLimit[0] , \PWMLimit[1] , 
            \PID_CONTROLLER.result[5] , n11, \PID_CONTROLLER.result[6] , 
            n13, \PID_CONTROLLER.result[7] , n15, \PWMLimit[8] , \PWMLimit[9] , 
            \PID_CONTROLLER.err[31] , n387, n11_adj_10, n24384, pwm, 
            clk32MHz, n24383, n24382, n24381, n24380, n42011, n24377, 
            n24376, n24375, n24374, n24373, n24372, n24371, n24370, 
            n24369, n24365, n24364, n24363, n24362, n24358, \deadband[9] , 
            \pwm_23__N_2951[5] , \pwm_23__N_2951[6] , n13_adj_11, n15_adj_12, 
            \pwm_23__N_2951[7] , pwm_23__N_2948, \Ki[7] , \Ki[3] , \Kp[1] , 
            \PID_CONTROLLER.err[7] , \Kp[0] , \PID_CONTROLLER.err[8] , 
            \Kp[2] , n11_adj_13, \Kp[3] , \PID_CONTROLLER.err[3] , \PID_CONTROLLER.err[13] , 
            n415, n414, n13_adj_14, \PID_CONTROLLER.err[14] , \deadband[0] , 
            n15_adj_15, \PID_CONTROLLER.err[0] , PIN_7_c_1, n413, \Kp[4] , 
            n421, \Ki[4] , \Kp[5] , \Kp[6] , \Ki[5] , \Kp[7] , \Kd[1] , 
            \Kd[0] , VCC_net, \Ki[6] , \Kd[2] , \Kd[3] , \Kd[4] , 
            \deadband[1] , \Kd[5] , \Kd[6] , \Kd[7] , \Ki[0] , \deadband[2] , 
            \deadband[3] , \deadband[4] , \Ki[1] , \PID_CONTROLLER.err[9] , 
            \PID_CONTROLLER.err[6] , \PID_CONTROLLER.err[5] , \PID_CONTROLLER.err[4] , 
            \PID_CONTROLLER.err[2] , \PID_CONTROLLER.err[1] , pwm_count, 
            \Ki[2] , \deadband[5] , \deadband[6] , \deadband[7] , \deadband[8] , 
            \PID_CONTROLLER.err[19] , \PID_CONTROLLER.err[20] , \PID_CONTROLLER.err[18] , 
            \PID_CONTROLLER.err[17] , IntegralLimit, \motor_state[23] , 
            \motor_state[22] , \motor_state[21] , \motor_state[20] , \motor_state[19] , 
            \motor_state[18] , \motor_state[17] , \motor_state[16] , \motor_state[15] , 
            \motor_state[14] , \PID_CONTROLLER.err[22] , \PID_CONTROLLER.err[23] , 
            \motor_state[13] , \motor_state[12] , \motor_state[11] , \motor_state[10] , 
            \motor_state[9] , \motor_state[8] , \motor_state[7] , \motor_state[6] , 
            \motor_state[5] , \motor_state[4] , \motor_state[3] , \motor_state[2] , 
            \motor_state[1] , \PID_CONTROLLER.err[12] , \motor_state[0] , 
            \PID_CONTROLLER.err_prev[31] , \PID_CONTROLLER.err_prev[23] , 
            \PID_CONTROLLER.err_prev[22] , \PID_CONTROLLER.err_prev[21] , 
            \PID_CONTROLLER.err_prev[20] , \PID_CONTROLLER.err_prev[19] , 
            \PID_CONTROLLER.err_prev[18] , \PID_CONTROLLER.err_prev[17] , 
            \PID_CONTROLLER.err_prev[16] , \PID_CONTROLLER.err_prev[15] , 
            \PID_CONTROLLER.err_prev[14] , \PID_CONTROLLER.err_prev[13] , 
            \PID_CONTROLLER.err_prev[12] , \PID_CONTROLLER.err_prev[11] , 
            \PID_CONTROLLER.err_prev[10] , \PID_CONTROLLER.err_prev[9] , 
            \PID_CONTROLLER.err_prev[8] , \PID_CONTROLLER.err_prev[7] , 
            \PID_CONTROLLER.err_prev[6] , \PID_CONTROLLER.err_prev[5] , 
            \PID_CONTROLLER.err_prev[4] , \PID_CONTROLLER.err_prev[3] , 
            \PID_CONTROLLER.err_prev[2] , \PID_CONTROLLER.err_prev[1] , 
            \PID_CONTROLLER.err_prev[0] , n22, n21, n23900, n23899, 
            n23898, n23897, n23896, n23895, n23894, n23893, n23892, 
            n23891, n23890, n23889, n24, n23888, n23887, n23886, 
            n23885, n23884, n23883, n23882, n23881, n23880, n23879, 
            n23878, n20, n23877, n23, n19, n17, n48782, n18, 
            PIN_8_c_2, PIN_9_c_3, PIN_10_c_4, PIN_11_c_5, n868, \PID_CONTROLLER.err[10] , 
            \PID_CONTROLLER.err[11] , \PID_CONTROLLER.err[15] , \PID_CONTROLLER.err[16] , 
            \PID_CONTROLLER.err[21] , n869, n870, n871, PIN_6_c_0, 
            n872, n873, n874, n875, n47156, n23743, \PWMLimit[2] , 
            \PWMLimit[3] , hall3, \PWMLimit[5] , hall1, \PWMLimit[6] , 
            hall2, \PWMLimit[7] , n29, n30, n48778, n471, n470, 
            n469, n468, n467, n1, n28052, n1_adj_16, n463, n44626, 
            n462, n461, n460, n459, n458, n457, n456, n455, 
            n15_adj_17, n13_adj_18, n11_adj_19, setpoint, n47225, 
            n47180, n47182, n47188, n47186, n47184) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input \PWMLimit[4] ;
    input \PWMLimit[0] ;
    input \PWMLimit[1] ;
    output \PID_CONTROLLER.result[5] ;
    input n11;
    output \PID_CONTROLLER.result[6] ;
    input n13;
    output \PID_CONTROLLER.result[7] ;
    input n15;
    input \PWMLimit[8] ;
    input \PWMLimit[9] ;
    output \PID_CONTROLLER.err[31] ;
    output n387;
    input n11_adj_10;
    input n24384;
    output [23:0]pwm;
    input clk32MHz;
    input n24383;
    input n24382;
    input n24381;
    input n24380;
    input n42011;
    input n24377;
    input n24376;
    input n24375;
    input n24374;
    input n24373;
    input n24372;
    input n24371;
    input n24370;
    input n24369;
    input n24365;
    input n24364;
    input n24363;
    input n24362;
    input n24358;
    input \deadband[9] ;
    output \pwm_23__N_2951[5] ;
    output \pwm_23__N_2951[6] ;
    input n13_adj_11;
    input n15_adj_12;
    output \pwm_23__N_2951[7] ;
    output pwm_23__N_2948;
    input \Ki[7] ;
    input \Ki[3] ;
    input \Kp[1] ;
    output \PID_CONTROLLER.err[7] ;
    input \Kp[0] ;
    output \PID_CONTROLLER.err[8] ;
    input \Kp[2] ;
    input n11_adj_13;
    input \Kp[3] ;
    output \PID_CONTROLLER.err[3] ;
    output \PID_CONTROLLER.err[13] ;
    output n415;
    output n414;
    input n13_adj_14;
    output \PID_CONTROLLER.err[14] ;
    input \deadband[0] ;
    input n15_adj_15;
    output \PID_CONTROLLER.err[0] ;
    output PIN_7_c_1;
    output n413;
    input \Kp[4] ;
    output n421;
    input \Ki[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Ki[5] ;
    input \Kp[7] ;
    input \Kd[1] ;
    input \Kd[0] ;
    input VCC_net;
    input \Ki[6] ;
    input \Kd[2] ;
    input \Kd[3] ;
    input \Kd[4] ;
    input \deadband[1] ;
    input \Kd[5] ;
    input \Kd[6] ;
    input \Kd[7] ;
    input \Ki[0] ;
    input \deadband[2] ;
    input \deadband[3] ;
    input \deadband[4] ;
    input \Ki[1] ;
    output \PID_CONTROLLER.err[9] ;
    output \PID_CONTROLLER.err[6] ;
    output \PID_CONTROLLER.err[5] ;
    output \PID_CONTROLLER.err[4] ;
    output \PID_CONTROLLER.err[2] ;
    output \PID_CONTROLLER.err[1] ;
    output [8:0]pwm_count;
    input \Ki[2] ;
    input \deadband[5] ;
    input \deadband[6] ;
    input \deadband[7] ;
    input \deadband[8] ;
    output \PID_CONTROLLER.err[19] ;
    output \PID_CONTROLLER.err[20] ;
    output \PID_CONTROLLER.err[18] ;
    output \PID_CONTROLLER.err[17] ;
    input [23:0]IntegralLimit;
    input \motor_state[23] ;
    input \motor_state[22] ;
    input \motor_state[21] ;
    input \motor_state[20] ;
    input \motor_state[19] ;
    input \motor_state[18] ;
    input \motor_state[17] ;
    input \motor_state[16] ;
    input \motor_state[15] ;
    input \motor_state[14] ;
    output \PID_CONTROLLER.err[22] ;
    output \PID_CONTROLLER.err[23] ;
    input \motor_state[13] ;
    input \motor_state[12] ;
    input \motor_state[11] ;
    input \motor_state[10] ;
    input \motor_state[9] ;
    input \motor_state[8] ;
    input \motor_state[7] ;
    input \motor_state[6] ;
    input \motor_state[5] ;
    input \motor_state[4] ;
    input \motor_state[3] ;
    input \motor_state[2] ;
    input \motor_state[1] ;
    output \PID_CONTROLLER.err[12] ;
    input \motor_state[0] ;
    output \PID_CONTROLLER.err_prev[31] ;
    output \PID_CONTROLLER.err_prev[23] ;
    output \PID_CONTROLLER.err_prev[22] ;
    output \PID_CONTROLLER.err_prev[21] ;
    output \PID_CONTROLLER.err_prev[20] ;
    output \PID_CONTROLLER.err_prev[19] ;
    output \PID_CONTROLLER.err_prev[18] ;
    output \PID_CONTROLLER.err_prev[17] ;
    output \PID_CONTROLLER.err_prev[16] ;
    output \PID_CONTROLLER.err_prev[15] ;
    output \PID_CONTROLLER.err_prev[14] ;
    output \PID_CONTROLLER.err_prev[13] ;
    output \PID_CONTROLLER.err_prev[12] ;
    output \PID_CONTROLLER.err_prev[11] ;
    output \PID_CONTROLLER.err_prev[10] ;
    output \PID_CONTROLLER.err_prev[9] ;
    output \PID_CONTROLLER.err_prev[8] ;
    output \PID_CONTROLLER.err_prev[7] ;
    output \PID_CONTROLLER.err_prev[6] ;
    output \PID_CONTROLLER.err_prev[5] ;
    output \PID_CONTROLLER.err_prev[4] ;
    output \PID_CONTROLLER.err_prev[3] ;
    output \PID_CONTROLLER.err_prev[2] ;
    output \PID_CONTROLLER.err_prev[1] ;
    output \PID_CONTROLLER.err_prev[0] ;
    output n22;
    output n21;
    input n23900;
    input n23899;
    input n23898;
    input n23897;
    input n23896;
    input n23895;
    input n23894;
    input n23893;
    input n23892;
    input n23891;
    input n23890;
    input n23889;
    output n24;
    input n23888;
    input n23887;
    input n23886;
    input n23885;
    input n23884;
    input n23883;
    input n23882;
    input n23881;
    input n23880;
    input n23879;
    input n23878;
    output n20;
    input n23877;
    output n23;
    output n19;
    output n17;
    input n48782;
    output n18;
    output PIN_8_c_2;
    output PIN_9_c_3;
    output PIN_10_c_4;
    output PIN_11_c_5;
    output n868;
    output \PID_CONTROLLER.err[10] ;
    output \PID_CONTROLLER.err[11] ;
    output \PID_CONTROLLER.err[15] ;
    output \PID_CONTROLLER.err[16] ;
    output \PID_CONTROLLER.err[21] ;
    output n869;
    output n870;
    output n871;
    output PIN_6_c_0;
    output n872;
    output n873;
    output n874;
    output n875;
    output n47156;
    input n23743;
    input \PWMLimit[2] ;
    input \PWMLimit[3] ;
    input hall3;
    input \PWMLimit[5] ;
    input hall1;
    input \PWMLimit[6] ;
    input hall2;
    input \PWMLimit[7] ;
    input n29;
    input n30;
    input n48778;
    output n471;
    output n470;
    output n469;
    output n468;
    output n467;
    input n1;
    input n28052;
    input n1_adj_16;
    output n463;
    output n44626;
    output n462;
    output n461;
    output n460;
    output n459;
    output n458;
    output n457;
    output n456;
    output n455;
    input n15_adj_17;
    input n13_adj_18;
    input n11_adj_19;
    input [23:0]setpoint;
    output n47225;
    output n47180;
    output n47182;
    output n47188;
    output n47186;
    output n47184;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n38854;
    wire [21:0]n8451;
    
    wire n38855;
    wire [25:0]n8081;
    wire [24:0]n8109;
    
    wire n501, n38233, n38614;
    wire [13:0]n15853;
    
    wire n38615, n38234;
    wire [25:0]n10674;
    wire [24:0]n11361;
    
    wire n37450;
    wire [22:0]n1804;
    
    wire n38853, n404, n38232, n37451, n37234;
    wire [17:0]n14796;
    
    wire n619, n37235;
    wire [18:0]n14437;
    
    wire n522, n37233, n37033;
    wire [23:0]n57;
    
    wire n37034;
    wire [14:0]n15643;
    
    wire n38613, n33, n37032;
    wire [9:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(26[22:30])
    
    wire n37449, n425, n37232, n38852, n307, n38231, n210, n38230, 
        n38612, n37448, n31, n37031, n38611, n38610, n38851, n38609, 
        n728, n38608, n38850, n20_c, n113, n536, n38849, n631, 
        n38607;
    wire [26:0]n8052;
    
    wire n38229, n534, n38606, n38228, n463_c, n38848, n437, n38605, 
        n38227, n38226, n340, n38604, n38225, n243, n38603, n390, 
        n38847, n53, n146, n317, n38846, n38224, n244, n38845;
    wire [6:0]n16623;
    wire [5:0]n16632;
    
    wire n752, n38602, n38223, n658, n38601, n38222, n558, n38600, 
        n171, n38844, n464_adj_3377, n38599, n38221, n370, n38598, 
        n35, n98, n37447, n276, n38597, n38220, n37446, n86, 
        n182, n38219, n328, n37231, n37445, n38218, n231, n37230, 
        n29_c, n37030;
    wire [12:0]n16034;
    
    wire n38596, n38217, n41, n134, n37444;
    wire [22:0]n1803;
    
    wire n38842, n1711, n27, n37029, n38216, n38841, n38595, n37443, 
        n38215, n38594, n38214;
    wire [8:0]n16508;
    wire [7:0]n16574;
    
    wire n37229, n37442, n37228, n25, n37028, n37441, n38213, 
        n38593, n746, n37227, n23_c, n37027, n38840, n38212, n38592, 
        n649, n37226, n37440, n37439, n552, n37225, n455_c, n37224, 
        n38211, n358, n37223, n37438, n21_c, n37026, n261, n37222, 
        n38591, n37437, n71, n164, n38210;
    wire [31:0]\PID_CONTROLLER.result ;   // verilog/motorControl.v(25[23:29])
    wire [31:0]pwm_23__N_2951;
    
    wire n19_c, n17_c, n7, n9_adj_3378, n38590, n692, n38209, 
        n595, n38208, n38839, n731, n38589, n498, n38207, n401, 
        n38206, n634, n38588, n304, n38205, n207, n38204, n38838, 
        n537_adj_3379, n38587, n17_adj_3380, n110;
    wire [27:0]n8022;
    
    wire n38203, n440, n38586, n38202, n38201, n38837, n343, n38585, 
        n38200, n38199, n246, n38584, n38198, n38197, n19_adj_3381, 
        n37025, n38836, n56, n149, n38196, n38195, n9_adj_3382;
    wire [11:0]n16188;
    
    wire n38583, n37436, n38194, n38582, n38193, n38835, n38192, 
        n38581, n38191, n38190, n38580, n38189, n38834, n4, n38188, 
        n38579, n48723, n38187, n38186, n48724, n38578, n38185, 
        n38833, n38184, n734, n38577, n38183, n47692, n48303, 
        n689, n38182, n637, n38576, n592, n38181, n38832, n495, 
        n38180, n540, n38575, n398, n38179, n6, n8_adj_3385, n48155, 
        n301, n38178, n443, n38574, n204, n38177, n48773, n38831, 
        n14_adj_3387, n107, n346, n38573;
    wire [28:0]n7991;
    
    wire n38176, n18_c, n38175, n38174, n249, n38572, n38173, 
        n38830, n38172, n59, n152, n38171, n38170;
    wire [10:0]n16317;
    
    wire n38571, n44807, n38169, n38829, n38570, n38168, n38167, 
        n38569, n44584, n38166, n26, n38165, n38828, n38568, n38164, 
        n38163, n38567, n38162, n38161, n38827, n737, n38566, 
        n38160, n38159, n640, n38565, n38158, n38157, n533, n38826, 
        n44823, n44578, n34, n543, n38564, n38156, n38155, n460_c, 
        n38825, n446, n38563, n686, n38154, n589, n38153, n349, 
        n38562, n492, n38152, n395, n38151, n387_c, n38824, n252, 
        n38561;
    wire [0:0]n5789;
    wire [29:0]n6545;
    
    wire n37636, n298, n38150;
    wire [55:0]n58;
    
    wire n37635, n201, n38149, n62, n155, n37634, n11_adj_3389, 
        n104, n37633;
    wire [0:0]n7064;
    wire [29:0]n7959;
    
    wire n38148;
    wire [31:0]n61;
    
    wire n49, n62_adj_3390, n44899, n314, n38823;
    wire [20:0]n8475;
    
    wire n38560;
    wire [55:0]n191;
    
    wire n38147, n37632, n38559, n38146, n37631, n38145, n37630, 
        n38558, n38144, n37629, n241, n38822, n38143, n37628, 
        n38557, n43221, n44883, n38142, n37627, n38141, n37626, 
        n38556, n38140, n37625, n168, n38821, n38139, n37624, 
        n38555, n56_adj_3392, n26_adj_3393, n95, n38138, n37623, 
        n38137, n37622, n38136, n37621, n38135, n38554, n37620, 
        n38134;
    wire [22:0]n1802;
    
    wire n38819, n44853, n37619, n38133, n38553, n37618, n38132, 
        n1707, n37617, n38131, n38552, n37616, n38130, n43147, 
        n38818, n37615, n38129, n38551, n37614, n38128, n37613, 
        n38127, n38550, n680_adj_3398, n37612, n38126, n38817, n583, 
        n37611, n38125, n38549, n486, n37610, n680_adj_3400, n38124, 
        n389, n37609, n583_adj_3402, n38123, n38548, n292, n37608, 
        n486_adj_3404, n38122, n38816, n195, n37607, n389_adj_3407, 
        n38121, n38547, n5, n98_adj_3408, n292_adj_3410, n38120, 
        n195_adj_3412, n38119, n38546, n5_adj_3414, n98_adj_3415, 
        n38815;
    wire [19:0]n9330;
    wire [18:0]n10121;
    
    wire n38118, n545, n38545, n38117, n4_adj_3416, n38116, n472, 
        n38544, n38115, n38814, n25_adj_3417, n38114, n399, n38543, 
        n38113;
    wire [28:0]n7763;
    
    wire n37599, n22_c, n38112, n37598, n326, n38542, n38111, 
        n37597, n30_c, n38813, n38110, n37596, n253, n38541, n38109, 
        n37595, n38108, n37594, n180, n38540, n38107, n37593, 
        n38812, n38106, n37592, n107_adj_3418, n28, n38105, n37591, 
        n29_adj_3419, n38104, n37590;
    wire [6:0]n8442;
    wire [5:0]n9322;
    
    wire n752_adj_3420, n38539, n38103, n37589, n27_adj_3421, n38811, 
        n655, n38538, n38102, n37588, n5_adj_3422, n47720, n8_adj_3424, 
        n42013, n6_adj_3425, n24368, n24367, n24366, n16_adj_3426, 
        n50, n47123, n47126, n4_adj_3427, n48727, n48728, n24_c, 
        n32, n36, n23_adj_3429, n47711, n38101, n47708, n49079, 
        n48153, n45055, n49221, n48337, n56_adj_3431, n60, n37587, 
        pwm_23__N_2950, n48769;
    wire [31:0]n63;
    
    wire n17_adj_3432, n43145, n14_adj_3433, n15_adj_3434, n6_adj_3435, 
        n583_adj_3436, n229_adj_3437, n119, n7_adj_3438, n9_adj_3439, 
        n26_adj_3440, n19_adj_3441, n216, n18_adj_3442, n24_adj_3443, 
        n5_adj_3444, n47660, n301_adj_3446, n137_adj_3447, n4_adj_3448, 
        n48721, n38100, n48722, n10_adj_3450, n22_adj_3451, n44, 
        n313, n12_adj_3452, n16_adj_3453, n26_adj_3454, n28729, n47241, 
        n37586, n25_adj_3455, n558_adj_3456, n38537, n6_adj_3457, 
        n48913;
    wire [31:0]n64;
    
    wire n48914, n37585, n37584, n37583, n44998, n658_adj_3459, 
        n38099, n37582, n234_adj_3460, n38810;
    wire [4:0]n10114;
    
    wire n564, n38098, n461_adj_3461, n38536, n464_adj_3462, n38097, 
        n37581;
    wire [2:0]n11529;
    
    wire n370_adj_3463, n38096, n37580, n364, n38535, n276_adj_3464, 
        n38095, n37579, n38809, n86_adj_3465, n182_adj_3466;
    wire [31:0]\PID_CONTROLLER.result_31__N_2994 ;
    
    wire n47635;
    wire [17:0]n10855;
    
    wire n38094;
    wire [24:0]\PID_CONTROLLER.err_31__N_2816 ;
    
    wire n38093;
    wire [5:0]PHASES_5__N_2779;
    
    wire n23569, n48163, n37578, n267, n38534, n38092, n37577, 
        n38808, n48591, n38091, n683_adj_3468, n37576, n410_adj_3469, 
        n170, n20_adj_3470, n38090, n586, n37575, n38807, n48775, 
        n331;
    wire [7:0]n8432;
    
    wire n38533, n38089, n489, n37574, n392, n37573, n749, n38532, 
        n38088, n302, n507, n295, n37572, n38806, n38087, n198, 
        n37571, n652, n38531, n38086, n8_adj_3471, n101, n38085;
    wire [27:0]n9128;
    
    wire n37570, n37569, n555, n38530, n38084, n37568, n38805, 
        n38083, n37567, n458_c, n38529, n38082, n17_adj_3472, n37024, 
        n37566, n604, n38081, n38804, n398_adj_3475, n38080, n38079, 
        n530, n38803, n38078, n38077, n457_c, n38802;
    wire [16:0]n11534;
    
    wire n38076, n38075, n384, n38801, n38074, n37565, n361, n38528, 
        n37435, n38073, n695, n37434, n311, n38800, n264, n38527, 
        n598, n37433, n38072, n74, n167, n38071, n501_adj_3477, 
        n37432, n238_adj_3479, n38799;
    wire [8:0]n8421;
    
    wire n38526, n38070, n38525, n404_adj_3480, n37431, n38069, 
        n307_adj_3481, n37430, n746_adj_3482, n38524, n38068, n210_adj_3483, 
        n37429;
    wire [31:0]n66;
    
    wire n37216, n38067, n20_adj_3484, n113_adj_3485, n37215, n165_adj_3486, 
        n38798, n649_adj_3487, n38523;
    wire [10:0]n14563;
    wire [9:0]n14915;
    
    wire n37428, n37214, n37427, n38066, n37213, n15_adj_3488, n37023, 
        n37426, n23_adj_3490, n92, n552_adj_3491, n38522, n37212, 
        n13_adj_3492, n37022, n38065, n37425, n37211, n455_adj_3494, 
        n38521, n37210, n11_adj_3495, n37021, n37424, n37209, n9_adj_3497, 
        n37020, n38064, n37208, n37423, n358_adj_3499, n38520, n37207, 
        n7_adj_3500, n37019;
    wire [22:0]n1801;
    
    wire n38796, n38063, n37422, n37206, n5_adj_3502, n37018, n37205, 
        n261_adj_3504, n38519, n37421, n3, n37017, n37204, n38062, 
        n37564, n375, n1703, n38061, n71_adj_3506, n164_adj_3507, 
        n38060, n38795, n37420;
    wire [9:0]n8409;
    
    wire n38518, n37563;
    wire [15:0]n12160;
    
    wire n38059, n37562, n37419, n38058, n38517, n38057, n428, 
        n38056, n38794, n38516, n38055, n701, n38054, n525, n37561, 
        n743, n38515, n38053, n38793, n646, n38514, n38052, n37203, 
        n37560, n622, n37559, n38051, n38792, n38050;
    wire [23:0]n11995;
    
    wire n37418, n549, n38513, n38049, n37558, n38048, n37417, 
        n452, n38512, n719, n38047, n355, n38511, n38046, n37557, 
        n37202, n38791, n38045, n37416, n38044, n38790, n258, 
        n38510, n37201, n140_adj_3508, n47;
    wire [23:0]n67;
    
    wire n37556, n37555, n448;
    wire [14:0]n12735;
    
    wire n38043, n37415, n68, n161, n38042, n38789, n38041;
    wire [10:0]n8396;
    
    wire n38509, n38040, n38508, n38039, n37554, n37414, n38038, 
        n38788, n38507, n38037, n38036, n38506, n38035, n37553, 
        n37413, n38034, n38787, n740, n38505, n38033, n38032, 
        n643, n38504, n38031, n37552, n37412, n38030, n38786, 
        n546, n38503, n38029, n449, n38502, n37551, n37411, n495_adj_3511, 
        n38785, n352, n38501, n255, n38500, n37550, n37410, n38784, 
        n65, n158;
    wire [11:0]n8382;
    
    wire n38499, n37549, n37409, n38498, n38783, n38497, n237_adj_3512, 
        n38496, n334, n38782, n37200, n686_adj_3513, n37548, n37408, 
        n589_adj_3514, n37547, n38781, n492_adj_3515, n37546, n38495, 
        n395_adj_3516, n37545, n527, n38780, n737_adj_3517, n38494, 
        n431, n640_adj_3518, n38493, n298_adj_3519, n37544, n37407, 
        n521, n543_adj_3520, n38492, n454, n38779, n446_adj_3522, 
        n38491, n349_adj_3523, n38490, n37199, n201_adj_3524, n37543, 
        n11_adj_3525, n104_adj_3526, n37406;
    wire [13:0]n13259;
    wire [12:0]n13737;
    
    wire n37542, n252_adj_3527, n38489, n37405, n62_adj_3529, n155_adj_3530, 
        n381, n38778, n37016, n592_adj_3531, n528_adj_3532, n625, 
        n689_adj_3533, n722;
    wire [33:0]n282;
    
    wire n308, n38777, n143_adj_3536, n235_adj_3538, n38776, n50_adj_3539, 
        n162, n38775, n240_adj_3540, n337, n20_adj_3541, n89;
    wire [22:0]n1800;
    
    wire n38773, n434, n531_adj_3542, n1699, n38772;
    wire [12:0]n8367;
    
    wire n38488, n37541, n38487, n37198, n37540, n38486, n37539, 
        n628, n38771, n725, n38485;
    wire [6:0]n69;
    wire [6:0]Kd_delay_counter;   // verilog/motorControl.v(20[13:29])
    
    wire n38484, n37538, n38483, n734_adj_3543, n38482, n38770, 
        n37404, n38769, n637_adj_3544, n38481, n540_adj_3545, n38480, 
        n37403, n37197, n37015, n443_adj_3547, n38479, n38768, n346_adj_3548, 
        n38478, n37402, n37537, n249_adj_3549, n38477, n38767, n59_adj_3550, 
        n152_adj_3551, n37536, n37401, n37535, n38766;
    wire [13:0]n8351;
    
    wire n38476, n38475, n698, n37400, n38474, n37534, n601_adj_3552, 
        n37399, n86_adj_3553, n38765;
    wire [9:0]n70;
    
    wire n37982, n38473, n37981, n37980, n37533, n38764, n38472, 
        n504, n37398, n37979, n37978, n38471, n37977, n38763, 
        n17_adj_3557, n37976, n37975, n37532, n37196, n407, n37397, 
        n38470, n37974, n38762, n731_adj_3559, n38469;
    wire [8:0]n73;
    
    wire n37973, n37531, n37972, n310, n37396, n37971, n38761, 
        n634_adj_3561, n38468, n37970, n37195, n537_adj_3562, n38467, 
        n37530, n37969, n213, n37395, n37194, n440_adj_3564, n38466, 
        n37968, n37014, n38760, n37967, n343_adj_3568, n38465, n146_adj_3569, 
        n37966, n246_adj_3571, n38464;
    wire [26:0]n9932;
    
    wire n37529, n23_adj_3573, n116, n37965, n38759, n37964, n56_adj_3574, 
        n149_adj_3575, n53_adj_3576, n37963, n37962, n37961;
    wire [14:0]n8334;
    
    wire n38463, n38462, n37960, n37528, n37959, n37958;
    wire [8:0]n15229;
    
    wire n37394, n38758, n37013, n37393, n38461, n101_adj_3579, 
        n37957, n37956, n38460, n37527, n37955, n524, n38757, 
        n8_adj_3581, n38459, n37954, n37392, n37526, n37953, n451, 
        n38756, n38458, n37952, n37012, n38457, n37951, n198_adj_3584, 
        n37950, n37391, n37525, n37193, n37011, n38456, n37949, 
        n37390, n378, n38755, n37948, n728_adj_3586, n38455, n37947, 
        n37946, n37524, n295_adj_3587, n631_adj_3588, n38454, n305, 
        n38754, n37945, n243_adj_3589, n37944, n159, n534_adj_3590, 
        n38453, n37389, n37943, n392_adj_3591, n37523, n683_adj_3592, 
        n37942, n340_adj_3593, n232_adj_3595, n38753, n437_adj_3596, 
        n38452, n586_adj_3597, n37941, n489_adj_3598, n37940, n38451, 
        n37939, n37522, n38752, n38450, n37938, n37521, n37937, 
        n37388, n37387, n37192, n37936, n37935, n37520, n37934;
    wire [15:0]n8316;
    
    wire n38449, n37933, n38448, n37932, n37519, n37931, n38447, 
        n37010, n37386;
    wire [22:0]n1799;
    
    wire n38750, n38446, n37518, n37930, n37191, n1695, n38445, 
        n37929, n38444, n37928, n37517, n37927, n38749, n37926, 
        n38443, n37516, n37925, n37924, n38442, n37923, n38748, 
        n38747, n38441;
    wire [8:0]n7068;
    
    wire n37922, n37921, n37515, n38440, n37920, n38439, n37919, 
        n37918, n38746, n37917, n38438, n37514, n37916, n38745, 
        n37915, n38437, n37914, n38744, n38436, n37913, n37190;
    wire [22:0]n12578;
    
    wire n37379, n38435, n37912, n37513, n37378, n37911, n37910, 
        n38743, n37909, n37189;
    wire [16:0]n8297;
    
    wire n38434, n37908, n37512, n37377, n38742, n38433, n37907, 
        n37906, n38432, n37905, n37904, n37376, n38741, n37903, 
        n37511, n38431, n38430, n37902, n37901, n38740, n38429, 
        n37900, n37375, n37899, n37188, n37374, n37510, n37898, 
        n37187, n37186, n38428, n37897, n38739, n37896, n37373, 
        n38738, n38427, n37895, n37009, n37894, n37509, n37372, 
        n38737;
    wire [16:0]n15117;
    
    wire n37185, n37184, n37008, n38736, n38426, n37893, n37892, 
        n38425, n37183, n37371, n37891, n37182, n38424, n37890, 
        n37508, n38735, n37889, n38423, n37888, n37887, n37370, 
        n37181, n38422, n37180, n37886, n37507, n37179, n37007, 
        n37369, n37368, n38734, n38421, n37367, n38420, n37178, 
        n37177, n38419, n37366, n37506, n37176, n37175, n37365, 
        n38733, n37364, n37174, n37173, n37363;
    wire [17:0]n8277;
    
    wire n38418, n37172, n37362, n38417, n37171, n38732, n38416, 
        n37505, n37361, n38415, n37360, n38731, n37170, n37359, 
        n38414, n37169, n37358, n37504, n38413, n37357, n38730, 
        n38412, n37356, n37355, n38411, n510, n37354, n156_adj_3626, 
        n38729, n38410, n38409, n204_adj_3627, n37503, n437_adj_3628, 
        n37353, n14_adj_3629, n83, n38408, n364_adj_3630, n37352, 
        n291, n37351, n719_adj_3632, n38407, n14_adj_3633, n107_adj_3634, 
        n622_adj_3635, n38406, n218_adj_3636, n37350;
    wire [22:0]n1798;
    
    wire n38727, n1691, n525_adj_3637, n38405, n145_adj_3638, n37349, 
        n38726, n428_adj_3639, n38404;
    wire [11:0]n14171;
    
    wire n37502, n72, n37501, n38725, n331_adj_3640, n38403;
    wire [21:0]n13112;
    
    wire n37348, n234_adj_3641, n38402, n37500, n37347, n37346, 
        n44_adj_3642, n137_adj_3643, n38724, n37499, n37345, n38723;
    wire [18:0]n8256;
    
    wire n38401, n37344, n38400, n37343, n37342, n38722, n38399, 
        n37498, n38398, n37341, n38721, n38397, n38720, n38396, 
        n37497, n37340, n38395, n37339;
    wire [24:0]n75;
    
    wire n37145, n37144, n37143, n55_adj_3646, n38394, n38719, n37496, 
        n37338, n37142, n37141, n37337, n37140, n38393, n37139, 
        n38718, n38392, n37336, n37138, n38717, n38391, n37137, 
        n37335, n37136, n38390, n37495, n37334, n37135, n716, 
        n38389, n38716, n619_adj_3655, n38388, n37134, n37333, n37133, 
        n38715, n522_adj_3658, n38387, n37494, n704, n37332, n37132, 
        n607_adj_3660, n37331, n37131, n37130, n38714, n510_adj_3663, 
        n37330, n425_adj_3664, n38386, n37129, n413_adj_3666, n37329, 
        n37128, n38713, n38712, n328_adj_3669, n38385, n37127, n316_adj_3671, 
        n37328, n37126, n219_adj_3673, n37327, n231_adj_3674, n38384, 
        n37125, n518, n38711, n37124, n29_adj_3677, n122, n37123, 
        n37122;
    wire [9:0]n16423;
    
    wire n37326, n41_adj_3681, n134_adj_3682, n37325, n445, n38710, 
        n37324, n37323;
    wire [19:0]n8234;
    
    wire n38383, n38382, n38381, n740_adj_3684, n37322, n643_adj_3685, 
        n37321, n372, n38709, n38380, n546_adj_3686, n37320, n299_adj_3688, 
        n38708, n449_adj_3689, n37319, n38379, n37493, n226_adj_3691, 
        n38707, n352_adj_3692, n37318, n153_adj_3694, n38706, n255_adj_3695, 
        n37317, n38378, n38377, n65_adj_3696, n158_adj_3697, n11_adj_3698, 
        n80;
    wire [20:0]n13597;
    
    wire n37316, n37315, n38376, n37314, n37313, n38375, n37312;
    wire [22:0]n1797;
    
    wire n38704, n37311, n38374, n37310, n1687, n37309, n38373, 
        n37308, n37307, n38703, n37306, n38372, n37492, n37305, 
        n37304, n38702, n38371, n713, n38370, n37303, n37491, 
        n37302, n616, n38369, n38701, n519_adj_3699, n38368, n422, 
        n38367, n38700, n325, n38366, n707, n37301, n228_adj_3700, 
        n38365, n38_adj_3701, n131_adj_3702, n38699;
    wire [20:0]n8211;
    
    wire n38364, n38363, n38698, n38362, n610_adj_3703, n37300, 
        n513, n37299, n38697, n38361, n416_adj_3704, n37298, n38360, 
        n319, n37297;
    wire [31:0]n76;
    
    wire n37097, n37096, n38696, n222_adj_3706, n37296, n37095, 
        n37094, n32_adj_3711, n125, n38695, n38359;
    wire [19:0]n14038;
    
    wire n37295, n37093, n37294, n37092, n38358, n37091, n37293, 
        n37090, n38357, n37089, n37490, n37292, n37088, n38694, 
        n38356, n38355, n37489, n37291, n37087, n37086, n37085, 
        n38354, n37290, n38693, n38353, n37084, n38352, n38692, 
        n38351, n710, n38350, n38691, n38893, n37488, n613, n38349, 
        n38892, n37289, n516, n38348, n38891, n37083, n37288, 
        n38690, n37082, n37287, n37081, n37286, n37487, n37285, 
        n38689, n37080, n419_adj_3731, n38347, n37284, n37079, n322, 
        n38346, n225_adj_3733, n38345, n37078, n37283, n37077, n37076, 
        n37075, n38890, n515, n38688, n37282, n37074, n37073, 
        n35_adj_3741, n128_adj_3742, n710_adj_3743, n37281, n613_adj_3745, 
        n37280, PHASES_5__N_3046, n37072;
    wire [23:0]n852;
    wire [23:0]n79;
    
    wire n37071, n516_adj_3749, n37279, n419_adj_3750, n37278;
    wire [21:0]n8187;
    
    wire n38344, n442, n38687, n322_adj_3752, n37277, n38889, n38343, 
        n37070, n38342, n225_adj_3755, n37276, n35_adj_3756, n128_adj_3757, 
        n369, n38686, n37069, n37068, n296_adj_3764, n38685, n38341, 
        n38888, n37275, n37067, n37274, n38340, n37273, n37066, 
        n38339, n37065, n743_adj_3769, n37272, n37064, n223_adj_3772, 
        n38684, n38338, n37063, n646_adj_3774, n37271, n37062, n38337, 
        n37486, n549_adj_3777, n37270, n150_adj_3779, n38683, n37061, 
        n10_adj_3782, n10_adj_3783, n43196, n43194, n452_adj_3784, 
        n37269, n37060, n38336, n37059, n8_adj_3787, n77, n38335, 
        n38887, n37485, n355_adj_3788, n37268, n37058, n38334, n37057;
    wire [22:0]n1796;
    
    wire n38681, n258_adj_3791, n37267, n38333, n1683, n68_adj_3792, 
        n161_adj_3793, n38332, n38680, n37266, n37265, n37056, n38331, 
        n38679, n37264, n37055, n38886, n37484, n38678, n38330, 
        n37263, n37262, n37054, n707_adj_3797, n38329, n37261, n12_adj_3798, 
        n38677, n610_adj_3799, n38328, n37260, n37259, n37053, n513_adj_3801, 
        n38327, n37258, n37052, n416_adj_3803, n38326, n37051, n38676, 
        n319_adj_3805, n38325, n37257, n222_adj_3806, n38324, n37256, 
        n37483, n38675, n32_adj_3807, n125_adj_3808, n37255, n37050, 
        n37482, n28495, n37254;
    wire [22:0]n8162;
    
    wire n38323, n713_adj_3811, n37253, n616_adj_3812, n37252, n38885, 
        n38322, n38674, n38321, n519_adj_3813, n37251, n6_adj_3814, 
        n37049, n38320, n422_adj_3815, n37250, n37048, n38673;
    wire [31:0]n82;
    
    wire n37047, n325_adj_3817, n37249, n38884, n38672, n38319, 
        n38671, n38318, n38883, n38317, n38670, n38316, n38315, 
        n38669, n38314, n38882, n38313, n38668, n38312, n38311, 
        n38667, n38310, n38881, n38309, n38666, n38308, n704_adj_3818, 
        n38307, n512, n38665, n607_adj_3819, n38306, n38880, n510_adj_3820, 
        n38305, n439, n38664, n413_adj_3821, n38304, n316_adj_3822, 
        n38303, n366, n38663, n219_adj_3823, n38302, n38879, n29_adj_3824, 
        n122_adj_3825, n293, n38662;
    wire [23:0]n8136;
    
    wire n38301, n38300, n38299, n220_adj_3826, n38661, n38298, 
        n38878, n38297, n147_adj_3827, n38660, n38296, n37046, n228_adj_3829, 
        n37248, n37045, n38_adj_3831, n131_adj_3832, n38295, n5_adj_3833, 
        n74_adj_3834, n37247, n37246, n38294, n38877, n37044, n37043, 
        n37245, n37042, n37244, n38293;
    wire [15:0]n15402;
    
    wire n38659, n37041, n37243, n37242, n38292, n38658, n37481, 
        n38657, n38876, n38656, n37040, n37241, n37039, n45_adj_3843, 
        n37038, n37240, n38291, n43_adj_3845, n37037, n37239, n37238, 
        n38290, n38655, n38875, n41_adj_3847, n37036, n39_adj_3849, 
        n37035, n37237, n37_adj_3851, n37236, n38289, n35_adj_3853, 
        n716_adj_3854, n38288, n38654, n38653, n38874, n38652, n37480, 
        n37479, n38287, n37478, n37477, n38286, n38651, n38873, 
        n37476, n37475, n38285, n37474, n37473, n701_adj_3855, n38284, 
        n38650, n37472, n37471, n692_adj_3856, n37470, n595_adj_3857, 
        n37469, n722_adj_3858, n38649, n38872, n498_adj_3859, n37468, 
        n401_adj_3860, n37467, n304_adj_3861, n37466, n207_adj_3862, 
        n37465, n625_adj_3863, n38648, n17_adj_3864, n110_adj_3865, 
        n37464, n604_adj_3866, n38283, n37463, n37462, n507_adj_3867, 
        n38282, n528_adj_3868, n38647, n38871, n37461, n37460, n410_adj_3869, 
        n38281, n37459, n37458, n313_adj_3870, n38280, n431_adj_3871, 
        n38646, n37457, n37456, n37455, n37454, n334_adj_3872, n38645, 
        n38870, n37453, n37452, n237_adj_3873, n38644, n216_adj_3874, 
        n38279, n26_adj_3875, n119_adj_3876, n47_adj_3877, n140_adj_3878, 
        n38869, n38278, n38277, n38643, n749_adj_3879, n38642, n38868, 
        n652_adj_3880, n38641, n38276, n555_adj_3881, n38640, n38275, 
        n38867, n38274, n458_adj_3882, n38639, n38273, n361_adj_3883, 
        n38638, n38866, n264_adj_3884, n38637, n38272, n167_adj_3885, 
        n38271, n38270, n38636, n38269, n38635, n38268, n38267, 
        n38634, n38865, n38266, n38265, n38633, n38864, n38264, 
        n38263, n38632, n38262, n38261, n38631, n38863, n698_adj_3886, 
        n38260, n601_adj_3887, n38259, n38630, n504_adj_3888, n38258, 
        n407_adj_3889, n38257, n38629, n38862, n38628, n725_adj_3890, 
        n38627, n38861, n628_adj_3891, n38626, n531_adj_3892, n38625, 
        n38860, n310_adj_3893, n38256, n213_adj_3894, n38255, n434_adj_3895, 
        n38624, n23_adj_3896, n116_adj_3897, n38254, n337_adj_3898, 
        n38623, n38859, n38253, n38252, n240_adj_3899, n38622, n38251, 
        n38250, n50_adj_3900, n143_adj_3901, n38858, n38249, n38248, 
        n44573, n38621, n38247;
    wire [4:0]n16640;
    
    wire n38620, n38246, n38857, n38245;
    wire [3:0]n16647;
    
    wire n38619, n38244, n38243;
    wire [2:0]n16653;
    
    wire n38618, n38242, n38856, n38241, n38617, n38240, n38239, 
        n38238, n38237, n38616, n38236, n695_adj_3902, n38235, n598_adj_3903, 
        n36452, n6_adj_3904, n9_adj_3905, n7_adj_3906, n43578, n880, 
        n892, n911, n19566, n19600, n934, n22310, n19608, n878, 
        n36747, n19292, n902_adj_3909, n4_adj_3910, n7_adj_3911, n24_adj_3912, 
        n26_adj_3913, n25_adj_3914, n27_adj_3915, n17_adj_3916, n20352, 
        n44847, n6_adj_3917;
    wire [5:0]PHASES_5__N_3039;
    
    wire n47234, n44840, n47079, n16801, n36732, n8_adj_3918, n8_adj_3919, 
        n47229, n44015, n44039, n47230, n44079, n44081, n47192, 
        n19615, n44011, n12_adj_3922, n47227, n7_adj_3928, n9_adj_3929, 
        n17_adj_3930, n48413, n48409, n48423, n48391, n48375, n30_adj_3934, 
        n48431, n48665, n48417, n48903, n47808, n48651, n49063, 
        n49207, n6_adj_3935, n48735, n48347, n24_adj_3936, n47757, 
        n50294, n8_adj_3937, n48997, n48143, n4_adj_3938, n48731, 
        n47787, n50272, n10_adj_3939, n49105, n48145, n49227, n49228, 
        n47761, n49180, n48151, n49223, n38898, n8_adj_3940, n18_adj_3941, 
        n24_adj_3942, n22_adj_3943, n26_adj_3944, n45037, n11_adj_3945, 
        n9_adj_3946, n17_adj_3947, n48465, n48463, n47856, n50467, 
        n48469, n48457, n47870, n50455, n10_adj_3948, n30_adj_3949, 
        n5_adj_3950, n48473, n48471, n47886, n48685, n49077, n48459, 
        n48909, n49146, n49245, n6_adj_3951, n47955, n24_adj_3952, 
        n48743, n47862, n50420, n48761, n48131, n4_adj_3953, n48737, 
        n48738, n8_adj_3954, n47850, n6_adj_3955, n16_adj_3956, n47852, 
        n48871, n48141, n49127, n4_adj_3957, n48741, n47872, n49103, 
        n48133, n49225, n49226, n48445, n49011, n48139, n49128, 
        n49125, n6_adj_3958, n4_adj_3959;
    
    SB_CARRY mult_14_add_1219_13 (.CI(n38854), .I0(n8451[10]), .I1(GND_net), 
            .CO(n38855));
    SB_LUT4 add_3088_6_lut (.I0(GND_net), .I1(n8109[3]), .I2(n501), .I3(n38233), 
            .O(n8081[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_14 (.CI(n38614), .I0(n15853[11]), .I1(GND_net), 
            .CO(n38615));
    SB_CARRY add_3088_6 (.CI(n38233), .I0(n8109[3]), .I1(n501), .CO(n38234));
    SB_LUT4 add_3198_24_lut (.I0(GND_net), .I1(n11361[21]), .I2(GND_net), 
            .I3(n37450), .O(n10674[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_12_lut (.I0(GND_net), .I1(n8451[9]), .I2(GND_net), 
            .I3(n38853), .O(n1804[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_5_lut (.I0(GND_net), .I1(n8109[2]), .I2(n404), .I3(n38232), 
            .O(n8081[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_5 (.CI(n38232), .I0(n8109[2]), .I1(n404), .CO(n38233));
    SB_CARRY add_3198_24 (.CI(n37450), .I0(n11361[21]), .I1(GND_net), 
            .CO(n37451));
    SB_CARRY add_3363_7 (.CI(n37234), .I0(n14796[4]), .I1(n619), .CO(n37235));
    SB_LUT4 add_3363_6_lut (.I0(GND_net), .I1(n14796[3]), .I2(n522), .I3(n37233), 
            .O(n14437[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n37033), .I0(GND_net), .I1(n57[17]), 
            .CO(n37034));
    SB_LUT4 add_3432_13_lut (.I0(GND_net), .I1(n15853[10]), .I2(GND_net), 
            .I3(n38613), .O(n15643[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_12 (.CI(n38853), .I0(n8451[9]), .I1(GND_net), 
            .CO(n38854));
    SB_CARRY add_3432_13 (.CI(n38613), .I0(n15853[10]), .I1(GND_net), 
            .CO(n38614));
    SB_CARRY add_3363_6 (.CI(n37233), .I0(n14796[3]), .I1(n522), .CO(n37234));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[16]), .I3(n37032), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3198_23_lut (.I0(GND_net), .I1(n11361[20]), .I2(GND_net), 
            .I3(n37449), .O(n10674[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_5_lut (.I0(GND_net), .I1(n14796[2]), .I2(n425), .I3(n37232), 
            .O(n14437[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n37032), .I0(GND_net), .I1(n57[16]), 
            .CO(n37033));
    SB_LUT4 mult_14_add_1219_11_lut (.I0(GND_net), .I1(n8451[8]), .I2(GND_net), 
            .I3(n38852), .O(n1804[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_4_lut (.I0(GND_net), .I1(n8109[1]), .I2(n307), .I3(n38231), 
            .O(n8081[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_4 (.CI(n38231), .I0(n8109[1]), .I1(n307), .CO(n38232));
    SB_LUT4 add_3088_3_lut (.I0(GND_net), .I1(n8109[0]), .I2(n210), .I3(n38230), 
            .O(n8081[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_23 (.CI(n37449), .I0(n11361[20]), .I1(GND_net), 
            .CO(n37450));
    SB_LUT4 add_3432_12_lut (.I0(GND_net), .I1(n15853[9]), .I2(GND_net), 
            .I3(n38612), .O(n15643[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_12 (.CI(n38612), .I0(n15853[9]), .I1(GND_net), .CO(n38613));
    SB_LUT4 add_3198_22_lut (.I0(GND_net), .I1(n11361[19]), .I2(GND_net), 
            .I3(n37448), .O(n10674[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[15]), .I3(n37031), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3432_11_lut (.I0(GND_net), .I1(n15853[8]), .I2(GND_net), 
            .I3(n38611), .O(n15643[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_11 (.CI(n38852), .I0(n8451[8]), .I1(GND_net), 
            .CO(n38853));
    SB_CARRY add_3432_11 (.CI(n38611), .I0(n15853[8]), .I1(GND_net), .CO(n38612));
    SB_LUT4 add_3432_10_lut (.I0(GND_net), .I1(n15853[7]), .I2(GND_net), 
            .I3(n38610), .O(n15643[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_10 (.CI(n38610), .I0(n15853[7]), .I1(GND_net), .CO(n38611));
    SB_LUT4 mult_14_add_1219_10_lut (.I0(GND_net), .I1(n8451[7]), .I2(GND_net), 
            .I3(n38851), .O(n1804[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_10 (.CI(n38851), .I0(n8451[7]), .I1(GND_net), 
            .CO(n38852));
    SB_LUT4 add_3432_9_lut (.I0(GND_net), .I1(n15853[6]), .I2(GND_net), 
            .I3(n38609), .O(n15643[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_3 (.CI(n38230), .I0(n8109[0]), .I1(n210), .CO(n38231));
    SB_CARRY add_3432_9 (.CI(n38609), .I0(n15853[6]), .I1(GND_net), .CO(n38610));
    SB_LUT4 add_3432_8_lut (.I0(GND_net), .I1(n15853[5]), .I2(n728), .I3(n38608), 
            .O(n15643[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_9_lut (.I0(GND_net), .I1(n8451[6]), .I2(GND_net), 
            .I3(n38850), .O(n1804[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_2_lut (.I0(GND_net), .I1(n20_c), .I2(n113), .I3(GND_net), 
            .O(n8081[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_9 (.CI(n38850), .I0(n8451[6]), .I1(GND_net), 
            .CO(n38851));
    SB_CARRY add_3088_2 (.CI(GND_net), .I0(n20_c), .I1(n113), .CO(n38230));
    SB_CARRY add_3198_22 (.CI(n37448), .I0(n11361[19]), .I1(GND_net), 
            .CO(n37449));
    SB_CARRY add_3363_5 (.CI(n37232), .I0(n14796[2]), .I1(n425), .CO(n37233));
    SB_LUT4 mult_14_add_1219_8_lut (.I0(GND_net), .I1(n8451[5]), .I2(n536), 
            .I3(n38849), .O(n1804[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_8 (.CI(n38608), .I0(n15853[5]), .I1(n728), .CO(n38609));
    SB_LUT4 add_3432_7_lut (.I0(GND_net), .I1(n15853[4]), .I2(n631), .I3(n38607), 
            .O(n15643[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_7 (.CI(n38607), .I0(n15853[4]), .I1(n631), .CO(n38608));
    SB_LUT4 add_3087_28_lut (.I0(GND_net), .I1(n8081[25]), .I2(GND_net), 
            .I3(n38229), .O(n8052[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_8 (.CI(n38849), .I0(n8451[5]), .I1(n536), 
            .CO(n38850));
    SB_LUT4 add_3432_6_lut (.I0(GND_net), .I1(n15853[3]), .I2(n534), .I3(n38606), 
            .O(n15643[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_27_lut (.I0(GND_net), .I1(n8081[24]), .I2(GND_net), 
            .I3(n38228), .O(n8052[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_6 (.CI(n38606), .I0(n15853[3]), .I1(n534), .CO(n38607));
    SB_CARRY add_3087_27 (.CI(n38228), .I0(n8081[24]), .I1(GND_net), .CO(n38229));
    SB_LUT4 mult_14_add_1219_7_lut (.I0(GND_net), .I1(n8451[4]), .I2(n463_c), 
            .I3(n38848), .O(n1804[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3432_5_lut (.I0(GND_net), .I1(n15853[2]), .I2(n437), .I3(n38605), 
            .O(n15643[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_26_lut (.I0(GND_net), .I1(n8081[23]), .I2(GND_net), 
            .I3(n38227), .O(n8052[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_5 (.CI(n38605), .I0(n15853[2]), .I1(n437), .CO(n38606));
    SB_CARRY add_3087_26 (.CI(n38227), .I0(n8081[23]), .I1(GND_net), .CO(n38228));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n37031), .I0(GND_net), .I1(n57[15]), 
            .CO(n37032));
    SB_LUT4 add_3087_25_lut (.I0(GND_net), .I1(n8081[22]), .I2(GND_net), 
            .I3(n38226), .O(n8052[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_7 (.CI(n38848), .I0(n8451[4]), .I1(n463_c), 
            .CO(n38849));
    SB_LUT4 add_3432_4_lut (.I0(GND_net), .I1(n15853[1]), .I2(n340), .I3(n38604), 
            .O(n15643[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_25 (.CI(n38226), .I0(n8081[22]), .I1(GND_net), .CO(n38227));
    SB_CARRY add_3432_4 (.CI(n38604), .I0(n15853[1]), .I1(n340), .CO(n38605));
    SB_LUT4 add_3087_24_lut (.I0(GND_net), .I1(n8081[21]), .I2(GND_net), 
            .I3(n38225), .O(n8052[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3432_3_lut (.I0(GND_net), .I1(n15853[0]), .I2(n243), .I3(n38603), 
            .O(n15643[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_6_lut (.I0(GND_net), .I1(n8451[3]), .I2(n390), 
            .I3(n38847), .O(n1804[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3432_3 (.CI(n38603), .I0(n15853[0]), .I1(n243), .CO(n38604));
    SB_CARRY mult_14_add_1219_6 (.CI(n38847), .I0(n8451[3]), .I1(n390), 
            .CO(n38848));
    SB_LUT4 add_3432_2_lut (.I0(GND_net), .I1(n53), .I2(n146), .I3(GND_net), 
            .O(n15643[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_5_lut (.I0(GND_net), .I1(n8451[2]), .I2(n317), 
            .I3(n38846), .O(n1804[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_24 (.CI(n38225), .I0(n8081[21]), .I1(GND_net), .CO(n38226));
    SB_CARRY add_3432_2 (.CI(GND_net), .I0(n53), .I1(n146), .CO(n38603));
    SB_LUT4 add_3087_23_lut (.I0(GND_net), .I1(n8081[20]), .I2(GND_net), 
            .I3(n38224), .O(n8052[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_5 (.CI(n38846), .I0(n8451[2]), .I1(n317), 
            .CO(n38847));
    SB_LUT4 mult_14_add_1219_4_lut (.I0(GND_net), .I1(n8451[1]), .I2(n244), 
            .I3(n38845), .O(n1804[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3516_8_lut (.I0(GND_net), .I1(n16632[5]), .I2(n752), .I3(n38602), 
            .O(n16623[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_23 (.CI(n38224), .I0(n8081[20]), .I1(GND_net), .CO(n38225));
    SB_LUT4 add_3087_22_lut (.I0(GND_net), .I1(n8081[19]), .I2(GND_net), 
            .I3(n38223), .O(n8052[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3516_7_lut (.I0(GND_net), .I1(n16632[4]), .I2(n658), .I3(n38601), 
            .O(n16623[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_22 (.CI(n38223), .I0(n8081[19]), .I1(GND_net), .CO(n38224));
    SB_CARRY mult_14_add_1219_4 (.CI(n38845), .I0(n8451[1]), .I1(n244), 
            .CO(n38846));
    SB_CARRY add_3516_7 (.CI(n38601), .I0(n16632[4]), .I1(n658), .CO(n38602));
    SB_LUT4 add_3087_21_lut (.I0(GND_net), .I1(n8081[18]), .I2(GND_net), 
            .I3(n38222), .O(n8052[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3516_6_lut (.I0(GND_net), .I1(n16632[3]), .I2(n558), .I3(n38600), 
            .O(n16623[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_3_lut (.I0(GND_net), .I1(n8451[0]), .I2(n171), 
            .I3(n38844), .O(n1804[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_6 (.CI(n38600), .I0(n16632[3]), .I1(n558), .CO(n38601));
    SB_CARRY add_3087_21 (.CI(n38222), .I0(n8081[18]), .I1(GND_net), .CO(n38223));
    SB_LUT4 add_3516_5_lut (.I0(GND_net), .I1(n16632[2]), .I2(n464_adj_3377), 
            .I3(n38599), .O(n16623[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_3 (.CI(n38844), .I0(n8451[0]), .I1(n171), 
            .CO(n38845));
    SB_LUT4 add_3087_20_lut (.I0(GND_net), .I1(n8081[17]), .I2(GND_net), 
            .I3(n38221), .O(n8052[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_5 (.CI(n38599), .I0(n16632[2]), .I1(n464_adj_3377), 
            .CO(n38600));
    SB_LUT4 add_3516_4_lut (.I0(GND_net), .I1(n16632[1]), .I2(n370), .I3(n38598), 
            .O(n16623[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_2_lut (.I0(GND_net), .I1(n35), .I2(n98), 
            .I3(GND_net), .O(n1804[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_21_lut (.I0(GND_net), .I1(n11361[18]), .I2(GND_net), 
            .I3(n37447), .O(n10674[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_20 (.CI(n38221), .I0(n8081[17]), .I1(GND_net), .CO(n38222));
    SB_CARRY add_3516_4 (.CI(n38598), .I0(n16632[1]), .I1(n370), .CO(n38599));
    SB_LUT4 add_3516_3_lut (.I0(GND_net), .I1(n16632[0]), .I2(n276), .I3(n38597), 
            .O(n16623[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_19_lut (.I0(GND_net), .I1(n8081[16]), .I2(GND_net), 
            .I3(n38220), .O(n8052[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3516_3 (.CI(n38597), .I0(n16632[0]), .I1(n276), .CO(n38598));
    SB_CARRY add_3198_21 (.CI(n37447), .I0(n11361[18]), .I1(GND_net), 
            .CO(n37448));
    SB_CARRY add_3087_19 (.CI(n38220), .I0(n8081[16]), .I1(GND_net), .CO(n38221));
    SB_LUT4 add_3198_20_lut (.I0(GND_net), .I1(n11361[17]), .I2(GND_net), 
            .I3(n37446), .O(n10674[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3516_2_lut (.I0(GND_net), .I1(n86), .I2(n182), .I3(GND_net), 
            .O(n16623[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3516_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_2 (.CI(GND_net), .I0(n35), .I1(n98), .CO(n38844));
    SB_CARRY add_3516_2 (.CI(GND_net), .I0(n86), .I1(n182), .CO(n38597));
    SB_LUT4 add_3087_18_lut (.I0(GND_net), .I1(n8081[15]), .I2(GND_net), 
            .I3(n38219), .O(n8052[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_4_lut (.I0(GND_net), .I1(n14796[1]), .I2(n328), .I3(n37231), 
            .O(n14437[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_20 (.CI(n37446), .I0(n11361[17]), .I1(GND_net), 
            .CO(n37447));
    SB_CARRY add_3087_18 (.CI(n38219), .I0(n8081[15]), .I1(GND_net), .CO(n38220));
    SB_LUT4 add_3198_19_lut (.I0(GND_net), .I1(n11361[16]), .I2(GND_net), 
            .I3(n37445), .O(n10674[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_4 (.CI(n37231), .I0(n14796[1]), .I1(n328), .CO(n37232));
    SB_LUT4 add_3087_17_lut (.I0(GND_net), .I1(n8081[14]), .I2(GND_net), 
            .I3(n38218), .O(n8052[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_3_lut (.I0(GND_net), .I1(n14796[0]), .I2(n231), .I3(n37230), 
            .O(n14437[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[14]), .I3(n37030), .O(n29_c)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3446_15_lut (.I0(GND_net), .I1(n16034[12]), .I2(GND_net), 
            .I3(n38596), .O(n15853[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_17 (.CI(n38218), .I0(n8081[14]), .I1(GND_net), .CO(n38219));
    SB_CARRY add_3198_19 (.CI(n37445), .I0(n11361[16]), .I1(GND_net), 
            .CO(n37446));
    SB_CARRY add_3363_3 (.CI(n37230), .I0(n14796[0]), .I1(n231), .CO(n37231));
    SB_LUT4 add_3087_16_lut (.I0(GND_net), .I1(n8081[13]), .I2(GND_net), 
            .I3(n38217), .O(n8052[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_2_lut (.I0(GND_net), .I1(n41), .I2(n134), .I3(GND_net), 
            .O(n14437[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n37030), .I0(GND_net), .I1(n57[14]), 
            .CO(n37031));
    SB_CARRY add_3087_16 (.CI(n38217), .I0(n8081[13]), .I1(GND_net), .CO(n38218));
    SB_LUT4 add_3198_18_lut (.I0(GND_net), .I1(n11361[15]), .I2(GND_net), 
            .I3(n37444), .O(n10674[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_24_lut (.I0(GND_net), .I1(n1804[21]), .I2(GND_net), 
            .I3(n38842), .O(n1803[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_24 (.CI(n38842), .I0(n1804[21]), .I1(GND_net), 
            .CO(n1711));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[13]), .I3(n37029), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n37029), .I0(GND_net), .I1(n57[13]), 
            .CO(n37030));
    SB_LUT4 add_3087_15_lut (.I0(GND_net), .I1(n8081[12]), .I2(GND_net), 
            .I3(n38216), .O(n8052[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_23_lut (.I0(GND_net), .I1(n1804[20]), .I2(GND_net), 
            .I3(n38841), .O(n1803[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_18 (.CI(n37444), .I0(n11361[15]), .I1(GND_net), 
            .CO(n37445));
    SB_CARRY add_3363_2 (.CI(GND_net), .I0(n41), .I1(n134), .CO(n37230));
    SB_LUT4 add_3446_14_lut (.I0(GND_net), .I1(n16034[11]), .I2(GND_net), 
            .I3(n38595), .O(n15853[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_14 (.CI(n38595), .I0(n16034[11]), .I1(GND_net), 
            .CO(n38596));
    SB_CARRY add_3087_15 (.CI(n38216), .I0(n8081[12]), .I1(GND_net), .CO(n38217));
    SB_LUT4 add_3198_17_lut (.I0(GND_net), .I1(n11361[14]), .I2(GND_net), 
            .I3(n37443), .O(n10674[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_14_lut (.I0(GND_net), .I1(n8081[11]), .I2(GND_net), 
            .I3(n38215), .O(n8052[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_14 (.CI(n38215), .I0(n8081[11]), .I1(GND_net), .CO(n38216));
    SB_LUT4 add_3446_13_lut (.I0(GND_net), .I1(n16034[10]), .I2(GND_net), 
            .I3(n38594), .O(n15853[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_13_lut (.I0(GND_net), .I1(n8081[10]), .I2(GND_net), 
            .I3(n38214), .O(n8052[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_17 (.CI(n37443), .I0(n11361[14]), .I1(GND_net), 
            .CO(n37444));
    SB_LUT4 add_3501_10_lut (.I0(GND_net), .I1(n16574[7]), .I2(GND_net), 
            .I3(n37229), .O(n16508[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_16_lut (.I0(GND_net), .I1(n11361[13]), .I2(GND_net), 
            .I3(n37442), .O(n10674[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3501_9_lut (.I0(GND_net), .I1(n16574[6]), .I2(GND_net), 
            .I3(n37228), .O(n16508[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[12]), .I3(n37028), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3446_13 (.CI(n38594), .I0(n16034[10]), .I1(GND_net), 
            .CO(n38595));
    SB_CARRY add_3087_13 (.CI(n38214), .I0(n8081[10]), .I1(GND_net), .CO(n38215));
    SB_CARRY add_3198_16 (.CI(n37442), .I0(n11361[13]), .I1(GND_net), 
            .CO(n37443));
    SB_LUT4 add_3198_15_lut (.I0(GND_net), .I1(n11361[12]), .I2(GND_net), 
            .I3(n37441), .O(n10674[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3087_12_lut (.I0(GND_net), .I1(n8081[9]), .I2(GND_net), 
            .I3(n38213), .O(n8052[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n37028), .I0(GND_net), .I1(n57[12]), 
            .CO(n37029));
    SB_CARRY mult_14_add_1218_23 (.CI(n38841), .I0(n1804[20]), .I1(GND_net), 
            .CO(n38842));
    SB_LUT4 add_3446_12_lut (.I0(GND_net), .I1(n16034[9]), .I2(GND_net), 
            .I3(n38593), .O(n15853[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_9 (.CI(n37228), .I0(n16574[6]), .I1(GND_net), .CO(n37229));
    SB_CARRY add_3087_12 (.CI(n38213), .I0(n8081[9]), .I1(GND_net), .CO(n38214));
    SB_CARRY add_3198_15 (.CI(n37441), .I0(n11361[12]), .I1(GND_net), 
            .CO(n37442));
    SB_LUT4 add_3501_8_lut (.I0(GND_net), .I1(n16574[5]), .I2(n746), .I3(n37227), 
            .O(n16508[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[11]), .I3(n37027), .O(n23_c)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1218_22_lut (.I0(GND_net), .I1(n1804[19]), .I2(GND_net), 
            .I3(n38840), .O(n1803[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n37027), .I0(GND_net), .I1(n57[11]), 
            .CO(n37028));
    SB_CARRY add_3446_12 (.CI(n38593), .I0(n16034[9]), .I1(GND_net), .CO(n38594));
    SB_LUT4 add_3087_11_lut (.I0(GND_net), .I1(n8081[8]), .I2(GND_net), 
            .I3(n38212), .O(n8052[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_11_lut (.I0(GND_net), .I1(n16034[8]), .I2(GND_net), 
            .I3(n38592), .O(n15853[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_11 (.CI(n38212), .I0(n8081[8]), .I1(GND_net), .CO(n38213));
    SB_CARRY add_3501_8 (.CI(n37227), .I0(n16574[5]), .I1(n746), .CO(n37228));
    SB_LUT4 add_3501_7_lut (.I0(GND_net), .I1(n16574[4]), .I2(n649), .I3(n37226), 
            .O(n16508[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_14_lut (.I0(GND_net), .I1(n11361[11]), .I2(GND_net), 
            .I3(n37440), .O(n10674[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_7 (.CI(n37226), .I0(n16574[4]), .I1(n649), .CO(n37227));
    SB_CARRY add_3198_14 (.CI(n37440), .I0(n11361[11]), .I1(GND_net), 
            .CO(n37441));
    SB_LUT4 add_3198_13_lut (.I0(GND_net), .I1(n11361[10]), .I2(GND_net), 
            .I3(n37439), .O(n10674[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3501_6_lut (.I0(GND_net), .I1(n16574[3]), .I2(n552), .I3(n37225), 
            .O(n16508[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_6 (.CI(n37225), .I0(n16574[3]), .I1(n552), .CO(n37226));
    SB_LUT4 add_3501_5_lut (.I0(GND_net), .I1(n16574[2]), .I2(n455_c), 
            .I3(n37224), .O(n16508[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_11 (.CI(n38592), .I0(n16034[8]), .I1(GND_net), .CO(n38593));
    SB_LUT4 add_3087_10_lut (.I0(GND_net), .I1(n8081[7]), .I2(GND_net), 
            .I3(n38211), .O(n8052[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_13 (.CI(n37439), .I0(n11361[10]), .I1(GND_net), 
            .CO(n37440));
    SB_CARRY add_3501_5 (.CI(n37224), .I0(n16574[2]), .I1(n455_c), .CO(n37225));
    SB_LUT4 add_3501_4_lut (.I0(GND_net), .I1(n16574[1]), .I2(n358), .I3(n37223), 
            .O(n16508[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_12_lut (.I0(GND_net), .I1(n11361[9]), .I2(GND_net), 
            .I3(n37438), .O(n10674[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[10]), .I3(n37026), .O(n21_c)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3501_4 (.CI(n37223), .I0(n16574[1]), .I1(n358), .CO(n37224));
    SB_LUT4 add_3501_3_lut (.I0(GND_net), .I1(n16574[0]), .I2(n261), .I3(n37222), 
            .O(n16508[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_10_lut (.I0(GND_net), .I1(n16034[7]), .I2(GND_net), 
            .I3(n38591), .O(n15853[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_3 (.CI(n37222), .I0(n16574[0]), .I1(n261), .CO(n37223));
    SB_CARRY add_3087_10 (.CI(n38211), .I0(n8081[7]), .I1(GND_net), .CO(n38212));
    SB_CARRY add_3198_12 (.CI(n37438), .I0(n11361[9]), .I1(GND_net), .CO(n37439));
    SB_LUT4 add_3198_11_lut (.I0(GND_net), .I1(n11361[8]), .I2(GND_net), 
            .I3(n37437), .O(n10674[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_10 (.CI(n38591), .I0(n16034[7]), .I1(GND_net), .CO(n38592));
    SB_LUT4 add_3501_2_lut (.I0(GND_net), .I1(n71), .I2(n164), .I3(GND_net), 
            .O(n16508[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3501_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3501_2 (.CI(GND_net), .I0(n71), .I1(n164), .CO(n37222));
    SB_LUT4 add_3087_9_lut (.I0(GND_net), .I1(n8081[6]), .I2(GND_net), 
            .I3(n38210), .O(n8052[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_23__I_816_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(pwm_23__N_2951[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_c));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_816_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(pwm_23__N_2951[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_c));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_816_i7_2_lut (.I0(\PID_CONTROLLER.result [3]), .I1(pwm_23__N_2951[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 pwm_23__I_816_i9_2_lut (.I0(\PID_CONTROLLER.result [4]), .I1(pwm_23__N_2951[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3378));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n37026), .I0(GND_net), .I1(n57[10]), 
            .CO(n37027));
    SB_CARRY mult_14_add_1218_22 (.CI(n38840), .I0(n1804[19]), .I1(GND_net), 
            .CO(n38841));
    SB_LUT4 add_3446_9_lut (.I0(GND_net), .I1(n16034[6]), .I2(GND_net), 
            .I3(n38590), .O(n15853[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_9 (.CI(n38210), .I0(n8081[6]), .I1(GND_net), .CO(n38211));
    SB_LUT4 add_3087_8_lut (.I0(GND_net), .I1(n8081[5]), .I2(n692), .I3(n38209), 
            .O(n8052[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_9 (.CI(n38590), .I0(n16034[6]), .I1(GND_net), .CO(n38591));
    SB_CARRY add_3087_8 (.CI(n38209), .I0(n8081[5]), .I1(n692), .CO(n38210));
    SB_LUT4 add_3087_7_lut (.I0(GND_net), .I1(n8081[4]), .I2(n595), .I3(n38208), 
            .O(n8052[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_21_lut (.I0(GND_net), .I1(n1804[18]), .I2(GND_net), 
            .I3(n38839), .O(n1803[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_8_lut (.I0(GND_net), .I1(n16034[5]), .I2(n731), .I3(n38589), 
            .O(n15853[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_7 (.CI(n38208), .I0(n8081[4]), .I1(n595), .CO(n38209));
    SB_LUT4 add_3087_6_lut (.I0(GND_net), .I1(n8081[3]), .I2(n498), .I3(n38207), 
            .O(n8052[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_8 (.CI(n38589), .I0(n16034[5]), .I1(n731), .CO(n38590));
    SB_CARRY add_3087_6 (.CI(n38207), .I0(n8081[3]), .I1(n498), .CO(n38208));
    SB_LUT4 add_3087_5_lut (.I0(GND_net), .I1(n8081[2]), .I2(n401), .I3(n38206), 
            .O(n8052[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_21 (.CI(n38839), .I0(n1804[18]), .I1(GND_net), 
            .CO(n38840));
    SB_LUT4 add_3446_7_lut (.I0(GND_net), .I1(n16034[4]), .I2(n634), .I3(n38588), 
            .O(n15853[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_5 (.CI(n38206), .I0(n8081[2]), .I1(n401), .CO(n38207));
    SB_LUT4 add_3087_4_lut (.I0(GND_net), .I1(n8081[1]), .I2(n304), .I3(n38205), 
            .O(n8052[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_7 (.CI(n38588), .I0(n16034[4]), .I1(n634), .CO(n38589));
    SB_CARRY add_3087_4 (.CI(n38205), .I0(n8081[1]), .I1(n304), .CO(n38206));
    SB_LUT4 add_3087_3_lut (.I0(GND_net), .I1(n8081[0]), .I2(n207), .I3(n38204), 
            .O(n8052[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_20_lut (.I0(GND_net), .I1(n1804[17]), .I2(GND_net), 
            .I3(n38838), .O(n1803[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_6_lut (.I0(GND_net), .I1(n16034[3]), .I2(n537_adj_3379), 
            .I3(n38587), .O(n15853[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3087_3 (.CI(n38204), .I0(n8081[0]), .I1(n207), .CO(n38205));
    SB_LUT4 add_3087_2_lut (.I0(GND_net), .I1(n17_adj_3380), .I2(n110), 
            .I3(GND_net), .O(n8052[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3087_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3446_6 (.CI(n38587), .I0(n16034[3]), .I1(n537_adj_3379), 
            .CO(n38588));
    SB_CARRY add_3087_2 (.CI(GND_net), .I0(n17_adj_3380), .I1(n110), .CO(n38204));
    SB_LUT4 add_3086_29_lut (.I0(GND_net), .I1(n8052[26]), .I2(GND_net), 
            .I3(n38203), .O(n8022[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_20 (.CI(n38838), .I0(n1804[17]), .I1(GND_net), 
            .CO(n38839));
    SB_LUT4 add_3446_5_lut (.I0(GND_net), .I1(n16034[2]), .I2(n440), .I3(n38586), 
            .O(n15853[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_28_lut (.I0(GND_net), .I1(n8052[25]), .I2(GND_net), 
            .I3(n38202), .O(n8022[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_28 (.CI(n38202), .I0(n8052[25]), .I1(GND_net), .CO(n38203));
    SB_CARRY add_3446_5 (.CI(n38586), .I0(n16034[2]), .I1(n440), .CO(n38587));
    SB_LUT4 add_3086_27_lut (.I0(GND_net), .I1(n8052[24]), .I2(GND_net), 
            .I3(n38201), .O(n8022[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_27 (.CI(n38201), .I0(n8052[24]), .I1(GND_net), .CO(n38202));
    SB_LUT4 mult_14_add_1218_19_lut (.I0(GND_net), .I1(n1804[16]), .I2(GND_net), 
            .I3(n38837), .O(n1803[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_4_lut (.I0(GND_net), .I1(n16034[1]), .I2(n343), .I3(n38585), 
            .O(n15853[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_26_lut (.I0(GND_net), .I1(n8052[23]), .I2(GND_net), 
            .I3(n38200), .O(n8022[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_26 (.CI(n38200), .I0(n8052[23]), .I1(GND_net), .CO(n38201));
    SB_CARRY add_3446_4 (.CI(n38585), .I0(n16034[1]), .I1(n343), .CO(n38586));
    SB_LUT4 add_3086_25_lut (.I0(GND_net), .I1(n8052[22]), .I2(GND_net), 
            .I3(n38199), .O(n8022[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_25 (.CI(n38199), .I0(n8052[22]), .I1(GND_net), .CO(n38200));
    SB_CARRY mult_14_add_1218_19 (.CI(n38837), .I0(n1804[16]), .I1(GND_net), 
            .CO(n38838));
    SB_LUT4 add_3446_3_lut (.I0(GND_net), .I1(n16034[0]), .I2(n246), .I3(n38584), 
            .O(n15853[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_24_lut (.I0(GND_net), .I1(n8052[21]), .I2(GND_net), 
            .I3(n38198), .O(n8022[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_24 (.CI(n38198), .I0(n8052[21]), .I1(GND_net), .CO(n38199));
    SB_CARRY add_3446_3 (.CI(n38584), .I0(n16034[0]), .I1(n246), .CO(n38585));
    SB_LUT4 add_3086_23_lut (.I0(GND_net), .I1(n8052[20]), .I2(GND_net), 
            .I3(n38197), .O(n8022[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[9]), .I3(n37025), .O(n19_adj_3381)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3198_11 (.CI(n37437), .I0(n11361[8]), .I1(GND_net), .CO(n37438));
    SB_CARRY add_3086_23 (.CI(n38197), .I0(n8052[20]), .I1(GND_net), .CO(n38198));
    SB_LUT4 mult_14_add_1218_18_lut (.I0(GND_net), .I1(n1804[15]), .I2(GND_net), 
            .I3(n38836), .O(n1803[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3446_2_lut (.I0(GND_net), .I1(n56), .I2(n149), .I3(GND_net), 
            .O(n15853[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3446_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_22_lut (.I0(GND_net), .I1(n8052[19]), .I2(GND_net), 
            .I3(n38196), .O(n8022[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_22 (.CI(n38196), .I0(n8052[19]), .I1(GND_net), .CO(n38197));
    SB_CARRY add_3446_2 (.CI(GND_net), .I0(n56), .I1(n149), .CO(n38584));
    SB_LUT4 add_3086_21_lut (.I0(GND_net), .I1(n8052[18]), .I2(GND_net), 
            .I3(n38195), .O(n8022[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_21 (.CI(n38195), .I0(n8052[18]), .I1(GND_net), .CO(n38196));
    SB_LUT4 LessThan_20_i9_2_lut (.I0(\PWMLimit[4] ), .I1(\PID_CONTROLLER.result [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3382));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_14_add_1218_18 (.CI(n38836), .I0(n1804[15]), .I1(GND_net), 
            .CO(n38837));
    SB_LUT4 add_3459_14_lut (.I0(GND_net), .I1(n16188[11]), .I2(GND_net), 
            .I3(n38583), .O(n16034[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_10_lut (.I0(GND_net), .I1(n11361[7]), .I2(GND_net), 
            .I3(n37436), .O(n10674[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_20_lut (.I0(GND_net), .I1(n8052[17]), .I2(GND_net), 
            .I3(n38194), .O(n8022[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_20 (.CI(n38194), .I0(n8052[17]), .I1(GND_net), .CO(n38195));
    SB_LUT4 add_3459_13_lut (.I0(GND_net), .I1(n16188[10]), .I2(GND_net), 
            .I3(n38582), .O(n16034[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_19_lut (.I0(GND_net), .I1(n8052[16]), .I2(GND_net), 
            .I3(n38193), .O(n8022[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_19 (.CI(n38193), .I0(n8052[16]), .I1(GND_net), .CO(n38194));
    SB_LUT4 mult_14_add_1218_17_lut (.I0(GND_net), .I1(n1804[14]), .I2(GND_net), 
            .I3(n38835), .O(n1803[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_13 (.CI(n38582), .I0(n16188[10]), .I1(GND_net), 
            .CO(n38583));
    SB_LUT4 add_3086_18_lut (.I0(GND_net), .I1(n8052[15]), .I2(GND_net), 
            .I3(n38192), .O(n8022[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_18 (.CI(n38192), .I0(n8052[15]), .I1(GND_net), .CO(n38193));
    SB_LUT4 add_3459_12_lut (.I0(GND_net), .I1(n16188[9]), .I2(GND_net), 
            .I3(n38581), .O(n16034[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_17_lut (.I0(GND_net), .I1(n8052[14]), .I2(GND_net), 
            .I3(n38191), .O(n8022[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_17 (.CI(n38191), .I0(n8052[14]), .I1(GND_net), .CO(n38192));
    SB_CARRY mult_14_add_1218_17 (.CI(n38835), .I0(n1804[14]), .I1(GND_net), 
            .CO(n38836));
    SB_CARRY add_3459_12 (.CI(n38581), .I0(n16188[9]), .I1(GND_net), .CO(n38582));
    SB_LUT4 add_3086_16_lut (.I0(GND_net), .I1(n8052[13]), .I2(GND_net), 
            .I3(n38190), .O(n8022[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_16 (.CI(n38190), .I0(n8052[13]), .I1(GND_net), .CO(n38191));
    SB_LUT4 add_3459_11_lut (.I0(GND_net), .I1(n16188[8]), .I2(GND_net), 
            .I3(n38580), .O(n16034[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_15_lut (.I0(GND_net), .I1(n8052[12]), .I2(GND_net), 
            .I3(n38189), .O(n8022[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_15 (.CI(n38189), .I0(n8052[12]), .I1(GND_net), .CO(n38190));
    SB_LUT4 mult_14_add_1218_16_lut (.I0(GND_net), .I1(n1804[13]), .I2(GND_net), 
            .I3(n38834), .O(n1803[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i4_4_lut (.I0(\PWMLimit[0] ), .I1(\PID_CONTROLLER.result [1]), 
            .I2(\PWMLimit[1] ), .I3(\PID_CONTROLLER.result [0]), .O(n4));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_3459_11 (.CI(n38580), .I0(n16188[8]), .I1(GND_net), .CO(n38581));
    SB_LUT4 add_3086_14_lut (.I0(GND_net), .I1(n8052[11]), .I2(GND_net), 
            .I3(n38188), .O(n8022[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_14 (.CI(n38188), .I0(n8052[11]), .I1(GND_net), .CO(n38189));
    SB_LUT4 add_3459_10_lut (.I0(GND_net), .I1(n16188[7]), .I2(GND_net), 
            .I3(n38579), .O(n16034[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33221_3_lut (.I0(n4), .I1(\PID_CONTROLLER.result[5] ), .I2(n11), 
            .I3(GND_net), .O(n48723));   // verilog/motorControl.v(38[12:27])
    defparam i33221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3086_13_lut (.I0(GND_net), .I1(n8052[10]), .I2(GND_net), 
            .I3(n38187), .O(n8022[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_13 (.CI(n38187), .I0(n8052[10]), .I1(GND_net), .CO(n38188));
    SB_CARRY mult_14_add_1218_16 (.CI(n38834), .I0(n1804[13]), .I1(GND_net), 
            .CO(n38835));
    SB_CARRY add_3459_10 (.CI(n38579), .I0(n16188[7]), .I1(GND_net), .CO(n38580));
    SB_LUT4 add_3086_12_lut (.I0(GND_net), .I1(n8052[9]), .I2(GND_net), 
            .I3(n38186), .O(n8022[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33222_3_lut (.I0(n48723), .I1(\PID_CONTROLLER.result[6] ), 
            .I2(n13), .I3(GND_net), .O(n48724));   // verilog/motorControl.v(38[12:27])
    defparam i33222_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3086_12 (.CI(n38186), .I0(n8052[9]), .I1(GND_net), .CO(n38187));
    SB_LUT4 add_3459_9_lut (.I0(GND_net), .I1(n16188[6]), .I2(GND_net), 
            .I3(n38578), .O(n16034[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_11_lut (.I0(GND_net), .I1(n8052[8]), .I2(GND_net), 
            .I3(n38185), .O(n8022[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_11 (.CI(n38185), .I0(n8052[8]), .I1(GND_net), .CO(n38186));
    SB_LUT4 mult_14_add_1218_15_lut (.I0(GND_net), .I1(n1804[12]), .I2(GND_net), 
            .I3(n38833), .O(n1803[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_9 (.CI(n38578), .I0(n16188[6]), .I1(GND_net), .CO(n38579));
    SB_LUT4 add_3086_10_lut (.I0(GND_net), .I1(n8052[7]), .I2(GND_net), 
            .I3(n38184), .O(n8022[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_10 (.CI(n38184), .I0(n8052[7]), .I1(GND_net), .CO(n38185));
    SB_LUT4 add_3459_8_lut (.I0(GND_net), .I1(n16188[5]), .I2(n734), .I3(n38577), 
            .O(n16034[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_9_lut (.I0(GND_net), .I1(n8052[6]), .I2(GND_net), 
            .I3(n38183), .O(n8022[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_9 (.CI(n38183), .I0(n8052[6]), .I1(GND_net), .CO(n38184));
    SB_CARRY mult_14_add_1218_15 (.CI(n38833), .I0(n1804[12]), .I1(GND_net), 
            .CO(n38834));
    SB_LUT4 i32801_4_lut (.I0(n13), .I1(n11), .I2(n9_adj_3382), .I3(n47692), 
            .O(n48303));
    defparam i32801_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_3459_8 (.CI(n38577), .I0(n16188[5]), .I1(n734), .CO(n38578));
    SB_LUT4 add_3086_8_lut (.I0(GND_net), .I1(n8052[5]), .I2(n689), .I3(n38182), 
            .O(n8022[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_8 (.CI(n38182), .I0(n8052[5]), .I1(n689), .CO(n38183));
    SB_LUT4 add_3459_7_lut (.I0(GND_net), .I1(n16188[4]), .I2(n637), .I3(n38576), 
            .O(n16034[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_7_lut (.I0(GND_net), .I1(n8052[4]), .I2(n592), .I3(n38181), 
            .O(n8022[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_7 (.CI(n38181), .I0(n8052[4]), .I1(n592), .CO(n38182));
    SB_LUT4 mult_14_add_1218_14_lut (.I0(GND_net), .I1(n1804[11]), .I2(GND_net), 
            .I3(n38832), .O(n1803[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_7 (.CI(n38576), .I0(n16188[4]), .I1(n637), .CO(n38577));
    SB_LUT4 add_3086_6_lut (.I0(GND_net), .I1(n8052[3]), .I2(n495), .I3(n38180), 
            .O(n8022[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_6 (.CI(n38180), .I0(n8052[3]), .I1(n495), .CO(n38181));
    SB_LUT4 add_3459_6_lut (.I0(GND_net), .I1(n16188[3]), .I2(n540), .I3(n38575), 
            .O(n16034[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_5_lut (.I0(GND_net), .I1(n8052[2]), .I2(n398), .I3(n38179), 
            .O(n8022[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_20_i8_3_lut (.I0(n6), .I1(\PID_CONTROLLER.result [4]), 
            .I2(n9_adj_3382), .I3(GND_net), .O(n8_adj_3385));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32653_3_lut (.I0(n48724), .I1(\PID_CONTROLLER.result[7] ), 
            .I2(n15), .I3(GND_net), .O(n48155));   // verilog/motorControl.v(38[12:27])
    defparam i32653_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3086_5 (.CI(n38179), .I0(n8052[2]), .I1(n398), .CO(n38180));
    SB_CARRY mult_14_add_1218_14 (.CI(n38832), .I0(n1804[11]), .I1(GND_net), 
            .CO(n38833));
    SB_CARRY add_3459_6 (.CI(n38575), .I0(n16188[3]), .I1(n540), .CO(n38576));
    SB_LUT4 add_3086_4_lut (.I0(GND_net), .I1(n8052[1]), .I2(n301), .I3(n38178), 
            .O(n8022[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_4 (.CI(n38178), .I0(n8052[1]), .I1(n301), .CO(n38179));
    SB_LUT4 add_3459_5_lut (.I0(GND_net), .I1(n16188[2]), .I2(n443), .I3(n38574), 
            .O(n16034[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3086_3_lut (.I0(GND_net), .I1(n8052[0]), .I2(n204), .I3(n38177), 
            .O(n8022[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33271_4_lut (.I0(n48155), .I1(n8_adj_3385), .I2(n15), .I3(n48303), 
            .O(n48773));   // verilog/motorControl.v(38[12:27])
    defparam i33271_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_3086_3 (.CI(n38177), .I0(n8052[0]), .I1(n204), .CO(n38178));
    SB_LUT4 mult_14_add_1218_13_lut (.I0(GND_net), .I1(n1804[10]), .I2(GND_net), 
            .I3(n38831), .O(n1803[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_5 (.CI(n38574), .I0(n16188[2]), .I1(n443), .CO(n38575));
    SB_LUT4 add_3086_2_lut (.I0(GND_net), .I1(n14_adj_3387), .I2(n107), 
            .I3(GND_net), .O(n8022[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3086_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3086_2 (.CI(GND_net), .I0(n14_adj_3387), .I1(n107), .CO(n38177));
    SB_LUT4 add_3459_4_lut (.I0(GND_net), .I1(n16188[1]), .I2(n346), .I3(n38573), 
            .O(n16034[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3085_30_lut (.I0(GND_net), .I1(n8022[27]), .I2(GND_net), 
            .I3(n38176), .O(n7991[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33272_3_lut (.I0(n48773), .I1(\PID_CONTROLLER.result [8]), 
            .I2(\PWMLimit[8] ), .I3(GND_net), .O(n18_c));   // verilog/motorControl.v(38[12:27])
    defparam i33272_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3085_29_lut (.I0(GND_net), .I1(n8022[26]), .I2(GND_net), 
            .I3(n38175), .O(n7991[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_13 (.CI(n38831), .I0(n1804[10]), .I1(GND_net), 
            .CO(n38832));
    SB_CARRY add_3459_4 (.CI(n38573), .I0(n16188[1]), .I1(n346), .CO(n38574));
    SB_CARRY add_3085_29 (.CI(n38175), .I0(n8022[26]), .I1(GND_net), .CO(n38176));
    SB_LUT4 add_3085_28_lut (.I0(GND_net), .I1(n8022[25]), .I2(GND_net), 
            .I3(n38174), .O(n7991[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3459_3_lut (.I0(GND_net), .I1(n16188[0]), .I2(n249), .I3(n38572), 
            .O(n16034[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_28 (.CI(n38174), .I0(n8022[25]), .I1(GND_net), .CO(n38175));
    SB_LUT4 add_3085_27_lut (.I0(GND_net), .I1(n8022[24]), .I2(GND_net), 
            .I3(n38173), .O(n7991[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_12_lut (.I0(GND_net), .I1(n1804[9]), .I2(GND_net), 
            .I3(n38830), .O(n1803[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3459_3 (.CI(n38572), .I0(n16188[0]), .I1(n249), .CO(n38573));
    SB_CARRY add_3085_27 (.CI(n38173), .I0(n8022[24]), .I1(GND_net), .CO(n38174));
    SB_LUT4 add_3085_26_lut (.I0(GND_net), .I1(n8022[23]), .I2(GND_net), 
            .I3(n38172), .O(n7991[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3459_2_lut (.I0(GND_net), .I1(n59), .I2(n152), .I3(GND_net), 
            .O(n16034[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3459_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_26 (.CI(n38172), .I0(n8022[23]), .I1(GND_net), .CO(n38173));
    SB_LUT4 add_3085_25_lut (.I0(GND_net), .I1(n8022[22]), .I2(GND_net), 
            .I3(n38171), .O(n7991[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_12 (.CI(n38830), .I0(n1804[9]), .I1(GND_net), 
            .CO(n38831));
    SB_CARRY add_3459_2 (.CI(GND_net), .I0(n59), .I1(n152), .CO(n38572));
    SB_CARRY add_3085_25 (.CI(n38171), .I0(n8022[22]), .I1(GND_net), .CO(n38172));
    SB_LUT4 add_3085_24_lut (.I0(GND_net), .I1(n8022[21]), .I2(GND_net), 
            .I3(n38170), .O(n7991[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_13_lut (.I0(GND_net), .I1(n16317[10]), .I2(GND_net), 
            .I3(n38571), .O(n16188[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n18_c), .I2(\PID_CONTROLLER.result [9]), 
            .I3(\PID_CONTROLLER.result [10]), .O(n44807));   // verilog/motorControl.v(38[12:27])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3085_24 (.CI(n38170), .I0(n8022[21]), .I1(GND_net), .CO(n38171));
    SB_LUT4 add_3085_23_lut (.I0(GND_net), .I1(n8022[20]), .I2(GND_net), 
            .I3(n38169), .O(n7991[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_11_lut (.I0(GND_net), .I1(n1804[8]), .I2(GND_net), 
            .I3(n38829), .O(n1803[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_12_lut (.I0(GND_net), .I1(n16317[9]), .I2(GND_net), 
            .I3(n38570), .O(n16188[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_23 (.CI(n38169), .I0(n8022[20]), .I1(GND_net), .CO(n38170));
    SB_LUT4 add_3085_22_lut (.I0(GND_net), .I1(n8022[19]), .I2(GND_net), 
            .I3(n38168), .O(n7991[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_12 (.CI(n38570), .I0(n16317[9]), .I1(GND_net), .CO(n38571));
    SB_CARRY add_3085_22 (.CI(n38168), .I0(n8022[19]), .I1(GND_net), .CO(n38169));
    SB_LUT4 add_3085_21_lut (.I0(GND_net), .I1(n8022[18]), .I2(GND_net), 
            .I3(n38167), .O(n7991[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_11 (.CI(n38829), .I0(n1804[8]), .I1(GND_net), 
            .CO(n38830));
    SB_LUT4 add_3471_11_lut (.I0(GND_net), .I1(n16317[8]), .I2(GND_net), 
            .I3(n38569), .O(n16188[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_21 (.CI(n38167), .I0(n8022[18]), .I1(GND_net), .CO(n38168));
    SB_LUT4 i2_4_lut (.I0(n18_c), .I1(\PID_CONTROLLER.result [10]), .I2(\PID_CONTROLLER.result [9]), 
            .I3(\PID_CONTROLLER.result [11]), .O(n44584));   // verilog/motorControl.v(38[12:27])
    defparam i2_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3085_20_lut (.I0(GND_net), .I1(n8022[17]), .I2(GND_net), 
            .I3(n38166), .O(n7991[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_11 (.CI(n38569), .I0(n16317[8]), .I1(GND_net), .CO(n38570));
    SB_CARRY add_3085_20 (.CI(n38166), .I0(n8022[17]), .I1(GND_net), .CO(n38167));
    SB_LUT4 i1_4_lut (.I0(\PID_CONTROLLER.result [12]), .I1(\PWMLimit[9] ), 
            .I2(n44584), .I3(n44807), .O(n26));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut.LUT_INIT = 16'hb3a2;
    SB_LUT4 add_3085_19_lut (.I0(GND_net), .I1(n8022[16]), .I2(GND_net), 
            .I3(n38165), .O(n7991[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_10_lut (.I0(GND_net), .I1(n1804[7]), .I2(GND_net), 
            .I3(n38828), .O(n1803[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_10_lut (.I0(GND_net), .I1(n16317[7]), .I2(GND_net), 
            .I3(n38568), .O(n16188[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_19 (.CI(n38165), .I0(n8022[16]), .I1(GND_net), .CO(n38166));
    SB_LUT4 add_3085_18_lut (.I0(GND_net), .I1(n8022[15]), .I2(GND_net), 
            .I3(n38164), .O(n7991[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_10 (.CI(n38568), .I0(n16317[7]), .I1(GND_net), .CO(n38569));
    SB_CARRY add_3085_18 (.CI(n38164), .I0(n8022[15]), .I1(GND_net), .CO(n38165));
    SB_LUT4 add_3085_17_lut (.I0(GND_net), .I1(n8022[14]), .I2(GND_net), 
            .I3(n38163), .O(n7991[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_10 (.CI(n38828), .I0(n1804[7]), .I1(GND_net), 
            .CO(n38829));
    SB_LUT4 add_3471_9_lut (.I0(GND_net), .I1(n16317[6]), .I2(GND_net), 
            .I3(n38567), .O(n16188[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_17 (.CI(n38163), .I0(n8022[14]), .I1(GND_net), .CO(n38164));
    SB_LUT4 add_3085_16_lut (.I0(GND_net), .I1(n8022[13]), .I2(GND_net), 
            .I3(n38162), .O(n7991[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_9 (.CI(n38567), .I0(n16317[6]), .I1(GND_net), .CO(n38568));
    SB_CARRY add_3085_16 (.CI(n38162), .I0(n8022[13]), .I1(GND_net), .CO(n38163));
    SB_LUT4 add_3085_15_lut (.I0(GND_net), .I1(n8022[12]), .I2(GND_net), 
            .I3(n38161), .O(n7991[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_9_lut (.I0(GND_net), .I1(n1804[6]), .I2(GND_net), 
            .I3(n38827), .O(n1803[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_8_lut (.I0(GND_net), .I1(n16317[5]), .I2(n737), .I3(n38566), 
            .O(n16188[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_15 (.CI(n38161), .I0(n8022[12]), .I1(GND_net), .CO(n38162));
    SB_LUT4 add_3085_14_lut (.I0(GND_net), .I1(n8022[11]), .I2(GND_net), 
            .I3(n38160), .O(n7991[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_8 (.CI(n38566), .I0(n16317[5]), .I1(n737), .CO(n38567));
    SB_CARRY add_3085_14 (.CI(n38160), .I0(n8022[11]), .I1(GND_net), .CO(n38161));
    SB_LUT4 add_3085_13_lut (.I0(GND_net), .I1(n8022[10]), .I2(GND_net), 
            .I3(n38159), .O(n7991[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_9 (.CI(n38827), .I0(n1804[6]), .I1(GND_net), 
            .CO(n38828));
    SB_LUT4 add_3471_7_lut (.I0(GND_net), .I1(n16317[4]), .I2(n640), .I3(n38565), 
            .O(n16188[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_13 (.CI(n38159), .I0(n8022[10]), .I1(GND_net), .CO(n38160));
    SB_LUT4 add_3085_12_lut (.I0(GND_net), .I1(n8022[9]), .I2(GND_net), 
            .I3(n38158), .O(n7991[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_7 (.CI(n38565), .I0(n16317[4]), .I1(n640), .CO(n38566));
    SB_CARRY add_3085_12 (.CI(n38158), .I0(n8022[9]), .I1(GND_net), .CO(n38159));
    SB_LUT4 add_3085_11_lut (.I0(GND_net), .I1(n8022[8]), .I2(GND_net), 
            .I3(n38157), .O(n7991[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_8_lut (.I0(GND_net), .I1(n1804[5]), .I2(n533), 
            .I3(n38826), .O(n1803[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_8 (.CI(n38826), .I0(n1804[5]), .I1(n533), 
            .CO(n38827));
    SB_LUT4 i3_4_lut_adj_1403 (.I0(\PID_CONTROLLER.result [15]), .I1(n26), 
            .I2(\PID_CONTROLLER.result [13]), .I3(\PID_CONTROLLER.result [14]), 
            .O(n44823));   // verilog/motorControl.v(38[12:27])
    defparam i3_4_lut_adj_1403.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1404 (.I0(n26), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [13]), .I3(\PID_CONTROLLER.result [15]), 
            .O(n44578));   // verilog/motorControl.v(38[12:27])
    defparam i2_4_lut_adj_1404.LUT_INIT = 16'h8000;
    SB_LUT4 i1_4_lut_adj_1405 (.I0(\PID_CONTROLLER.result [16]), .I1(\PWMLimit[9] ), 
            .I2(n44578), .I3(n44823), .O(n34));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1405.LUT_INIT = 16'hb3a2;
    SB_LUT4 add_3471_6_lut (.I0(GND_net), .I1(n16317[3]), .I2(n543), .I3(n38564), 
            .O(n16188[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_11 (.CI(n38157), .I0(n8022[8]), .I1(GND_net), .CO(n38158));
    SB_LUT4 add_3085_10_lut (.I0(GND_net), .I1(n8022[7]), .I2(GND_net), 
            .I3(n38156), .O(n7991[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_6 (.CI(n38564), .I0(n16317[3]), .I1(n543), .CO(n38565));
    SB_CARRY add_3085_10 (.CI(n38156), .I0(n8022[7]), .I1(GND_net), .CO(n38157));
    SB_LUT4 add_3085_9_lut (.I0(GND_net), .I1(n8022[6]), .I2(GND_net), 
            .I3(n38155), .O(n7991[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_7_lut (.I0(GND_net), .I1(n1804[4]), .I2(n460_c), 
            .I3(n38825), .O(n1803[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_5_lut (.I0(GND_net), .I1(n16317[2]), .I2(n446), .I3(n38563), 
            .O(n16188[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_9 (.CI(n38155), .I0(n8022[6]), .I1(GND_net), .CO(n38156));
    SB_LUT4 add_3085_8_lut (.I0(GND_net), .I1(n8022[5]), .I2(n686), .I3(n38154), 
            .O(n7991[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_5 (.CI(n38563), .I0(n16317[2]), .I1(n446), .CO(n38564));
    SB_CARRY add_3085_8 (.CI(n38154), .I0(n8022[5]), .I1(n686), .CO(n38155));
    SB_LUT4 add_3085_7_lut (.I0(GND_net), .I1(n8022[4]), .I2(n589), .I3(n38153), 
            .O(n7991[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_7 (.CI(n38825), .I0(n1804[4]), .I1(n460_c), 
            .CO(n38826));
    SB_LUT4 add_3471_4_lut (.I0(GND_net), .I1(n16317[1]), .I2(n349), .I3(n38562), 
            .O(n16188[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_7 (.CI(n38153), .I0(n8022[4]), .I1(n589), .CO(n38154));
    SB_LUT4 add_3085_6_lut (.I0(GND_net), .I1(n8022[3]), .I2(n492), .I3(n38152), 
            .O(n7991[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_4 (.CI(n38562), .I0(n16317[1]), .I1(n349), .CO(n38563));
    SB_CARRY add_3085_6 (.CI(n38152), .I0(n8022[3]), .I1(n492), .CO(n38153));
    SB_LUT4 add_3085_5_lut (.I0(GND_net), .I1(n8022[2]), .I2(n395), .I3(n38151), 
            .O(n7991[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1218_6_lut (.I0(GND_net), .I1(n1804[3]), .I2(n387_c), 
            .I3(n38824), .O(n1803[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3471_3_lut (.I0(GND_net), .I1(n16317[0]), .I2(n252), .I3(n38561), 
            .O(n16188[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_5 (.CI(n38151), .I0(n8022[2]), .I1(n395), .CO(n38152));
    SB_LUT4 mult_10_add_2137_32_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(n6545[29]), 
            .I2(GND_net), .I3(n37636), .O(n5789[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3085_4_lut (.I0(GND_net), .I1(n8022[1]), .I2(n298), .I3(n38150), 
            .O(n7991[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_3 (.CI(n38561), .I0(n16317[0]), .I1(n252), .CO(n38562));
    SB_CARRY add_3085_4 (.CI(n38150), .I0(n8022[1]), .I1(n298), .CO(n38151));
    SB_LUT4 mult_10_add_2137_31_lut (.I0(GND_net), .I1(n6545[28]), .I2(GND_net), 
            .I3(n37635), .O(n58[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_31 (.CI(n37635), .I0(n6545[28]), .I1(GND_net), 
            .CO(n37636));
    SB_LUT4 add_3085_3_lut (.I0(GND_net), .I1(n8022[0]), .I2(n201), .I3(n38149), 
            .O(n7991[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_6 (.CI(n38824), .I0(n1804[3]), .I1(n387_c), 
            .CO(n38825));
    SB_LUT4 add_3471_2_lut (.I0(GND_net), .I1(n62), .I2(n155), .I3(GND_net), 
            .O(n16188[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3471_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3085_3 (.CI(n38149), .I0(n8022[0]), .I1(n201), .CO(n38150));
    SB_LUT4 mult_10_add_2137_30_lut (.I0(GND_net), .I1(n6545[27]), .I2(GND_net), 
            .I3(n37634), .O(n58[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_30 (.CI(n37634), .I0(n6545[27]), .I1(GND_net), 
            .CO(n37635));
    SB_LUT4 add_3085_2_lut (.I0(GND_net), .I1(n11_adj_3389), .I2(n104), 
            .I3(GND_net), .O(n7991[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3085_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3471_2 (.CI(GND_net), .I0(n62), .I1(n155), .CO(n38561));
    SB_CARRY add_3085_2 (.CI(GND_net), .I0(n11_adj_3389), .I1(n104), .CO(n38149));
    SB_LUT4 mult_10_add_2137_29_lut (.I0(GND_net), .I1(n6545[26]), .I2(GND_net), 
            .I3(n37633), .O(n58[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_29 (.CI(n37633), .I0(n6545[26]), .I1(GND_net), 
            .CO(n37634));
    SB_LUT4 mult_12_add_2137_32_lut (.I0(n61[25]), .I1(n7959[29]), .I2(GND_net), 
            .I3(n38148), .O(n7064[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_32_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1406 (.I0(\PID_CONTROLLER.result [26]), .I1(n34), 
            .I2(n49), .I3(n62_adj_3390), .O(n44899));   // verilog/motorControl.v(31[14] 52[8])
    defparam i3_4_lut_adj_1406.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_14_add_1218_5_lut (.I0(GND_net), .I1(n1804[2]), .I2(n314), 
            .I3(n38823), .O(n1803[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_23_lut (.I0(GND_net), .I1(n8475[20]), .I2(GND_net), 
            .I3(n38560), .O(n8451[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_31_lut (.I0(GND_net), .I1(n7959[28]), .I2(GND_net), 
            .I3(n38147), .O(n191[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_28_lut (.I0(GND_net), .I1(n6545[25]), .I2(GND_net), 
            .I3(n37632), .O(n58[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_28 (.CI(n37632), .I0(n6545[25]), .I1(GND_net), 
            .CO(n37633));
    SB_CARRY mult_12_add_2137_31 (.CI(n38147), .I0(n7959[28]), .I1(GND_net), 
            .CO(n38148));
    SB_LUT4 add_3108_22_lut (.I0(GND_net), .I1(n8475[19]), .I2(GND_net), 
            .I3(n38559), .O(n8451[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_30_lut (.I0(GND_net), .I1(n7959[27]), .I2(GND_net), 
            .I3(n38146), .O(n191[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_27_lut (.I0(GND_net), .I1(n6545[24]), .I2(GND_net), 
            .I3(n37631), .O(n58[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_27 (.CI(n37631), .I0(n6545[24]), .I1(GND_net), 
            .CO(n37632));
    SB_CARRY mult_12_add_2137_30 (.CI(n38146), .I0(n7959[27]), .I1(GND_net), 
            .CO(n38147));
    SB_CARRY mult_14_add_1218_5 (.CI(n38823), .I0(n1804[2]), .I1(n314), 
            .CO(n38824));
    SB_CARRY add_3108_22 (.CI(n38559), .I0(n8475[19]), .I1(GND_net), .CO(n38560));
    SB_LUT4 mult_12_add_2137_29_lut (.I0(GND_net), .I1(n7959[26]), .I2(GND_net), 
            .I3(n38145), .O(n191[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_26_lut (.I0(GND_net), .I1(n6545[23]), .I2(GND_net), 
            .I3(n37630), .O(n58[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_26 (.CI(n37630), .I0(n6545[23]), .I1(GND_net), 
            .CO(n37631));
    SB_CARRY mult_12_add_2137_29 (.CI(n38145), .I0(n7959[26]), .I1(GND_net), 
            .CO(n38146));
    SB_LUT4 add_3108_21_lut (.I0(GND_net), .I1(n8475[18]), .I2(GND_net), 
            .I3(n38558), .O(n8451[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_28_lut (.I0(GND_net), .I1(n7959[25]), .I2(GND_net), 
            .I3(n38144), .O(n191[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_25_lut (.I0(GND_net), .I1(n6545[22]), .I2(GND_net), 
            .I3(n37629), .O(n58[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_25 (.CI(n37629), .I0(n6545[22]), .I1(GND_net), 
            .CO(n37630));
    SB_CARRY mult_12_add_2137_28 (.CI(n38144), .I0(n7959[25]), .I1(GND_net), 
            .CO(n38145));
    SB_LUT4 mult_14_add_1218_4_lut (.I0(GND_net), .I1(n1804[1]), .I2(n241), 
            .I3(n38822), .O(n1803[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_21 (.CI(n38558), .I0(n8475[18]), .I1(GND_net), .CO(n38559));
    SB_LUT4 mult_12_add_2137_27_lut (.I0(GND_net), .I1(n7959[24]), .I2(GND_net), 
            .I3(n38143), .O(n191[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_24_lut (.I0(GND_net), .I1(n6545[21]), .I2(GND_net), 
            .I3(n37628), .O(n58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_24 (.CI(n37628), .I0(n6545[21]), .I1(GND_net), 
            .CO(n37629));
    SB_CARRY mult_12_add_2137_27 (.CI(n38143), .I0(n7959[24]), .I1(GND_net), 
            .CO(n38144));
    SB_LUT4 add_3108_20_lut (.I0(GND_net), .I1(n8475[17]), .I2(GND_net), 
            .I3(n38557), .O(n8451[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut (.I0(n43221), .I1(\PID_CONTROLLER.result [26]), .I2(n34), 
            .I3(GND_net), .O(n44883));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mult_12_add_2137_26_lut (.I0(GND_net), .I1(n7959[23]), .I2(GND_net), 
            .I3(n38142), .O(n191[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_23_lut (.I0(GND_net), .I1(n6545[20]), .I2(GND_net), 
            .I3(n37627), .O(n58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_23 (.CI(n37627), .I0(n6545[20]), .I1(GND_net), 
            .CO(n37628));
    SB_CARRY mult_12_add_2137_26 (.CI(n38142), .I0(n7959[23]), .I1(GND_net), 
            .CO(n38143));
    SB_CARRY mult_14_add_1218_4 (.CI(n38822), .I0(n1804[1]), .I1(n241), 
            .CO(n38823));
    SB_CARRY add_3108_20 (.CI(n38557), .I0(n8475[17]), .I1(GND_net), .CO(n38558));
    SB_LUT4 mult_12_add_2137_25_lut (.I0(GND_net), .I1(n7959[22]), .I2(GND_net), 
            .I3(n38141), .O(n191[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_22_lut (.I0(GND_net), .I1(n6545[19]), .I2(GND_net), 
            .I3(n37626), .O(n58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_22 (.CI(n37626), .I0(n6545[19]), .I1(GND_net), 
            .CO(n37627));
    SB_CARRY mult_12_add_2137_25 (.CI(n38141), .I0(n7959[22]), .I1(GND_net), 
            .CO(n38142));
    SB_LUT4 add_3108_19_lut (.I0(GND_net), .I1(n8475[16]), .I2(GND_net), 
            .I3(n38556), .O(n8451[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_24_lut (.I0(GND_net), .I1(n7959[21]), .I2(GND_net), 
            .I3(n38140), .O(n191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_21_lut (.I0(GND_net), .I1(n6545[18]), .I2(GND_net), 
            .I3(n37625), .O(n58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_21 (.CI(n37625), .I0(n6545[18]), .I1(GND_net), 
            .CO(n37626));
    SB_CARRY mult_12_add_2137_24 (.CI(n38140), .I0(n7959[21]), .I1(GND_net), 
            .CO(n38141));
    SB_LUT4 mult_14_add_1218_3_lut (.I0(GND_net), .I1(n1804[0]), .I2(n168), 
            .I3(n38821), .O(n1803[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_19 (.CI(n38556), .I0(n8475[16]), .I1(GND_net), .CO(n38557));
    SB_LUT4 mult_12_add_2137_23_lut (.I0(GND_net), .I1(n7959[20]), .I2(GND_net), 
            .I3(n38139), .O(n191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_2137_20_lut (.I0(GND_net), .I1(n6545[17]), .I2(GND_net), 
            .I3(n37624), .O(n58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_20 (.CI(n37624), .I0(n6545[17]), .I1(GND_net), 
            .CO(n37625));
    SB_CARRY mult_12_add_2137_23 (.CI(n38139), .I0(n7959[20]), .I1(GND_net), 
            .CO(n38140));
    SB_LUT4 add_3108_18_lut (.I0(GND_net), .I1(n8475[15]), .I2(GND_net), 
            .I3(n38555), .O(n8451[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1407 (.I0(\PID_CONTROLLER.result [27]), .I1(\PWMLimit[9] ), 
            .I2(n44883), .I3(n44899), .O(n56_adj_3392));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1407.LUT_INIT = 16'hb3a2;
    SB_CARRY mult_14_add_1218_3 (.CI(n38821), .I0(n1804[0]), .I1(n168), 
            .CO(n38822));
    SB_LUT4 mult_14_add_1218_2_lut (.I0(GND_net), .I1(n26_adj_3393), .I2(n95), 
            .I3(GND_net), .O(n1803[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1218_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_add_2137_22_lut (.I0(GND_net), .I1(n7959[19]), .I2(GND_net), 
            .I3(n38138), .O(n191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_22 (.CI(n38138), .I0(n7959[19]), .I1(GND_net), 
            .CO(n38139));
    SB_LUT4 mult_10_add_2137_19_lut (.I0(GND_net), .I1(n6545[16]), .I2(GND_net), 
            .I3(n37623), .O(n58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_19 (.CI(n37623), .I0(n6545[16]), .I1(GND_net), 
            .CO(n37624));
    SB_LUT4 mult_12_add_2137_21_lut (.I0(GND_net), .I1(n7959[18]), .I2(GND_net), 
            .I3(n38137), .O(n191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_21 (.CI(n38137), .I0(n7959[18]), .I1(GND_net), 
            .CO(n38138));
    SB_LUT4 mult_10_add_2137_18_lut (.I0(GND_net), .I1(n6545[15]), .I2(GND_net), 
            .I3(n37622), .O(n58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_18 (.CI(n37622), .I0(n6545[15]), .I1(GND_net), 
            .CO(n37623));
    SB_LUT4 mult_12_add_2137_20_lut (.I0(GND_net), .I1(n7959[17]), .I2(GND_net), 
            .I3(n38136), .O(n191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1218_2 (.CI(GND_net), .I0(n26_adj_3393), .I1(n95), 
            .CO(n38821));
    SB_CARRY add_3108_18 (.CI(n38555), .I0(n8475[15]), .I1(GND_net), .CO(n38556));
    SB_CARRY mult_12_add_2137_20 (.CI(n38136), .I0(n7959[17]), .I1(GND_net), 
            .CO(n38137));
    SB_LUT4 mult_10_add_2137_17_lut (.I0(GND_net), .I1(n6545[14]), .I2(GND_net), 
            .I3(n37621), .O(n58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_17 (.CI(n37621), .I0(n6545[14]), .I1(GND_net), 
            .CO(n37622));
    SB_LUT4 mult_12_add_2137_19_lut (.I0(GND_net), .I1(n7959[16]), .I2(GND_net), 
            .I3(n38135), .O(n191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_17_lut (.I0(GND_net), .I1(n8475[14]), .I2(GND_net), 
            .I3(n38554), .O(n8451[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_19 (.CI(n38135), .I0(n7959[16]), .I1(GND_net), 
            .CO(n38136));
    SB_LUT4 mult_10_add_2137_16_lut (.I0(GND_net), .I1(n6545[13]), .I2(GND_net), 
            .I3(n37620), .O(n58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_16 (.CI(n37620), .I0(n6545[13]), .I1(GND_net), 
            .CO(n37621));
    SB_LUT4 mult_12_add_2137_18_lut (.I0(GND_net), .I1(n7959[15]), .I2(GND_net), 
            .I3(n38134), .O(n191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_24_lut (.I0(GND_net), .I1(n1803[21]), .I2(GND_net), 
            .I3(n38819), .O(n1802[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1408 (.I0(\PID_CONTROLLER.result [30]), .I1(n56_adj_3392), 
            .I2(\PID_CONTROLLER.result [28]), .I3(\PID_CONTROLLER.result [29]), 
            .O(n44853));   // verilog/motorControl.v(38[12:27])
    defparam i3_4_lut_adj_1408.LUT_INIT = 16'hfffe;
    SB_CARRY add_3108_17 (.CI(n38554), .I0(n8475[14]), .I1(GND_net), .CO(n38555));
    SB_CARRY mult_12_add_2137_18 (.CI(n38134), .I0(n7959[15]), .I1(GND_net), 
            .CO(n38135));
    SB_LUT4 mult_10_add_2137_15_lut (.I0(GND_net), .I1(n6545[12]), .I2(GND_net), 
            .I3(n37619), .O(n58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_15 (.CI(n37619), .I0(n6545[12]), .I1(GND_net), 
            .CO(n37620));
    SB_LUT4 mult_12_add_2137_17_lut (.I0(GND_net), .I1(n7959[14]), .I2(GND_net), 
            .I3(n38133), .O(n191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_16_lut (.I0(GND_net), .I1(n8475[13]), .I2(GND_net), 
            .I3(n38553), .O(n8451[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_17 (.CI(n38133), .I0(n7959[14]), .I1(GND_net), 
            .CO(n38134));
    SB_LUT4 mult_10_add_2137_14_lut (.I0(GND_net), .I1(n6545[11]), .I2(GND_net), 
            .I3(n37618), .O(n58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_14 (.CI(n37618), .I0(n6545[11]), .I1(GND_net), 
            .CO(n37619));
    SB_LUT4 mult_12_add_2137_16_lut (.I0(GND_net), .I1(n7959[13]), .I2(GND_net), 
            .I3(n38132), .O(n191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_24 (.CI(n38819), .I0(n1803[21]), .I1(GND_net), 
            .CO(n1707));
    SB_CARRY add_3108_16 (.CI(n38553), .I0(n8475[13]), .I1(GND_net), .CO(n38554));
    SB_CARRY mult_12_add_2137_16 (.CI(n38132), .I0(n7959[13]), .I1(GND_net), 
            .CO(n38133));
    SB_LUT4 mult_10_add_2137_13_lut (.I0(GND_net), .I1(n6545[10]), .I2(GND_net), 
            .I3(n37617), .O(n58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_13 (.CI(n37617), .I0(n6545[10]), .I1(GND_net), 
            .CO(n37618));
    SB_LUT4 mult_12_add_2137_15_lut (.I0(GND_net), .I1(n7959[12]), .I2(GND_net), 
            .I3(n38131), .O(n191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_15_lut (.I0(GND_net), .I1(n8475[12]), .I2(GND_net), 
            .I3(n38552), .O(n8451[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_15 (.CI(n38131), .I0(n7959[12]), .I1(GND_net), 
            .CO(n38132));
    SB_LUT4 mult_10_add_2137_12_lut (.I0(GND_net), .I1(n6545[9]), .I2(GND_net), 
            .I3(n37616), .O(n58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_12 (.CI(n37616), .I0(n6545[9]), .I1(GND_net), 
            .CO(n37617));
    SB_LUT4 mult_12_add_2137_14_lut (.I0(GND_net), .I1(n7959[11]), .I2(GND_net), 
            .I3(n38130), .O(n191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1409 (.I0(\PWMLimit[9] ), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n43147), .I3(n44853), .O(n387));   // verilog/motorControl.v(38[12:27])
    defparam i1_4_lut_adj_1409.LUT_INIT = 16'hb3a2;
    SB_LUT4 mult_14_add_1217_23_lut (.I0(GND_net), .I1(n1803[20]), .I2(GND_net), 
            .I3(n38818), .O(n1802[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_15 (.CI(n38552), .I0(n8475[12]), .I1(GND_net), .CO(n38553));
    SB_CARRY mult_12_add_2137_14 (.CI(n38130), .I0(n7959[11]), .I1(GND_net), 
            .CO(n38131));
    SB_LUT4 mult_10_add_2137_11_lut (.I0(GND_net), .I1(n6545[8]), .I2(GND_net), 
            .I3(n37615), .O(n58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_11 (.CI(n37615), .I0(n6545[8]), .I1(GND_net), 
            .CO(n37616));
    SB_LUT4 mult_12_add_2137_13_lut (.I0(GND_net), .I1(n7959[10]), .I2(GND_net), 
            .I3(n38129), .O(n191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_14_lut (.I0(GND_net), .I1(n8475[11]), .I2(GND_net), 
            .I3(n38551), .O(n8451[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_13 (.CI(n38129), .I0(n7959[10]), .I1(GND_net), 
            .CO(n38130));
    SB_LUT4 mult_10_add_2137_10_lut (.I0(GND_net), .I1(n6545[7]), .I2(GND_net), 
            .I3(n37614), .O(n58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_10 (.CI(n37614), .I0(n6545[7]), .I1(GND_net), 
            .CO(n37615));
    SB_LUT4 mult_12_add_2137_12_lut (.I0(GND_net), .I1(n7959[9]), .I2(GND_net), 
            .I3(n38128), .O(n191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_23 (.CI(n38818), .I0(n1803[20]), .I1(GND_net), 
            .CO(n38819));
    SB_CARRY add_3108_14 (.CI(n38551), .I0(n8475[11]), .I1(GND_net), .CO(n38552));
    SB_CARRY mult_12_add_2137_12 (.CI(n38128), .I0(n7959[9]), .I1(GND_net), 
            .CO(n38129));
    SB_LUT4 mult_10_add_2137_9_lut (.I0(GND_net), .I1(n6545[6]), .I2(GND_net), 
            .I3(n37613), .O(n58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_9 (.CI(n37613), .I0(n6545[6]), .I1(GND_net), 
            .CO(n37614));
    SB_LUT4 mult_12_add_2137_11_lut (.I0(GND_net), .I1(n7959[8]), .I2(GND_net), 
            .I3(n38127), .O(n191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_13_lut (.I0(GND_net), .I1(n8475[10]), .I2(GND_net), 
            .I3(n38550), .O(n8451[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_11 (.CI(n38127), .I0(n7959[8]), .I1(GND_net), 
            .CO(n38128));
    SB_LUT4 mult_10_add_2137_8_lut (.I0(GND_net), .I1(n6545[5]), .I2(n680_adj_3398), 
            .I3(n37612), .O(n58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_8 (.CI(n37612), .I0(n6545[5]), .I1(n680_adj_3398), 
            .CO(n37613));
    SB_LUT4 mult_12_add_2137_10_lut (.I0(GND_net), .I1(n7959[7]), .I2(GND_net), 
            .I3(n38126), .O(n191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_22_lut (.I0(GND_net), .I1(n1803[19]), .I2(GND_net), 
            .I3(n38817), .O(n1802[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_13 (.CI(n38550), .I0(n8475[10]), .I1(GND_net), .CO(n38551));
    SB_CARRY mult_12_add_2137_10 (.CI(n38126), .I0(n7959[7]), .I1(GND_net), 
            .CO(n38127));
    SB_LUT4 mult_10_add_2137_7_lut (.I0(GND_net), .I1(n6545[4]), .I2(n583), 
            .I3(n37611), .O(n58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_7 (.CI(n37611), .I0(n6545[4]), .I1(n583), 
            .CO(n37612));
    SB_LUT4 mult_12_add_2137_9_lut (.I0(GND_net), .I1(n7959[6]), .I2(GND_net), 
            .I3(n38125), .O(n191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_12_lut (.I0(GND_net), .I1(n8475[9]), .I2(GND_net), 
            .I3(n38549), .O(n8451[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_9 (.CI(n38125), .I0(n7959[6]), .I1(GND_net), 
            .CO(n38126));
    SB_LUT4 mult_10_add_2137_6_lut (.I0(GND_net), .I1(n6545[3]), .I2(n486), 
            .I3(n37610), .O(n58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_6 (.CI(n37610), .I0(n6545[3]), .I1(n486), 
            .CO(n37611));
    SB_LUT4 mult_12_add_2137_8_lut (.I0(GND_net), .I1(n7959[5]), .I2(n680_adj_3400), 
            .I3(n38124), .O(n191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_22 (.CI(n38817), .I0(n1803[19]), .I1(GND_net), 
            .CO(n38818));
    SB_CARRY add_3108_12 (.CI(n38549), .I0(n8475[9]), .I1(GND_net), .CO(n38550));
    SB_CARRY mult_12_add_2137_8 (.CI(n38124), .I0(n7959[5]), .I1(n680_adj_3400), 
            .CO(n38125));
    SB_LUT4 mult_10_add_2137_5_lut (.I0(GND_net), .I1(n6545[2]), .I2(n389), 
            .I3(n37609), .O(n58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_5 (.CI(n37609), .I0(n6545[2]), .I1(n389), 
            .CO(n37610));
    SB_LUT4 mult_12_add_2137_7_lut (.I0(GND_net), .I1(n7959[4]), .I2(n583_adj_3402), 
            .I3(n38123), .O(n191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_11_lut (.I0(GND_net), .I1(n8475[8]), .I2(GND_net), 
            .I3(n38548), .O(n8451[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_7 (.CI(n38123), .I0(n7959[4]), .I1(n583_adj_3402), 
            .CO(n38124));
    SB_LUT4 mult_10_add_2137_4_lut (.I0(GND_net), .I1(n6545[1]), .I2(n292), 
            .I3(n37608), .O(n58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_4 (.CI(n37608), .I0(n6545[1]), .I1(n292), 
            .CO(n37609));
    SB_LUT4 mult_12_add_2137_6_lut (.I0(GND_net), .I1(n7959[3]), .I2(n486_adj_3404), 
            .I3(n38122), .O(n191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_21_lut (.I0(GND_net), .I1(n1803[18]), .I2(GND_net), 
            .I3(n38816), .O(n1802[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_11 (.CI(n38548), .I0(n8475[8]), .I1(GND_net), .CO(n38549));
    SB_CARRY mult_12_add_2137_6 (.CI(n38122), .I0(n7959[3]), .I1(n486_adj_3404), 
            .CO(n38123));
    SB_LUT4 mult_10_add_2137_3_lut (.I0(GND_net), .I1(n6545[0]), .I2(n195), 
            .I3(n37607), .O(n58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_3 (.CI(n37607), .I0(n6545[0]), .I1(n195), 
            .CO(n37608));
    SB_LUT4 mult_12_add_2137_5_lut (.I0(GND_net), .I1(n7959[2]), .I2(n389_adj_3407), 
            .I3(n38121), .O(n191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_10_lut (.I0(GND_net), .I1(n8475[7]), .I2(GND_net), 
            .I3(n38547), .O(n8451[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_5 (.CI(n38121), .I0(n7959[2]), .I1(n389_adj_3407), 
            .CO(n38122));
    SB_LUT4 mult_10_add_2137_2_lut (.I0(GND_net), .I1(n5), .I2(n98_adj_3408), 
            .I3(GND_net), .O(n58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_2137_2 (.CI(GND_net), .I0(n5), .I1(n98_adj_3408), 
            .CO(n37607));
    SB_LUT4 mult_12_add_2137_4_lut (.I0(GND_net), .I1(n7959[1]), .I2(n292_adj_3410), 
            .I3(n38120), .O(n191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_21 (.CI(n38816), .I0(n1803[18]), .I1(GND_net), 
            .CO(n38817));
    SB_CARRY add_3108_10 (.CI(n38547), .I0(n8475[7]), .I1(GND_net), .CO(n38548));
    SB_CARRY mult_12_add_2137_4 (.CI(n38120), .I0(n7959[1]), .I1(n292_adj_3410), 
            .CO(n38121));
    SB_LUT4 mult_12_add_2137_3_lut (.I0(GND_net), .I1(n7959[0]), .I2(n195_adj_3412), 
            .I3(n38119), .O(n191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_9_lut (.I0(GND_net), .I1(n8475[6]), .I2(GND_net), 
            .I3(n38546), .O(n8451[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_12_add_2137_3 (.CI(n38119), .I0(n7959[0]), .I1(n195_adj_3412), 
            .CO(n38120));
    SB_LUT4 mult_12_add_2137_2_lut (.I0(GND_net), .I1(n5_adj_3414), .I2(n98_adj_3415), 
            .I3(GND_net), .O(n191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_12_add_2137_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_20_lut (.I0(GND_net), .I1(n1803[17]), .I2(GND_net), 
            .I3(n38815), .O(n1802[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_9 (.CI(n38546), .I0(n8475[6]), .I1(GND_net), .CO(n38547));
    SB_CARRY mult_12_add_2137_2 (.CI(GND_net), .I0(n5_adj_3414), .I1(n98_adj_3415), 
            .CO(n38119));
    SB_LUT4 add_3149_21_lut (.I0(GND_net), .I1(n10121[18]), .I2(GND_net), 
            .I3(n38118), .O(n9330[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3108_8_lut (.I0(GND_net), .I1(n8475[5]), .I2(n545), .I3(n38545), 
            .O(n8451[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_20_lut (.I0(GND_net), .I1(n10121[17]), .I2(GND_net), 
            .I3(n38117), .O(n9330[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_20 (.CI(n38117), .I0(n10121[17]), .I1(GND_net), 
            .CO(n38118));
    SB_LUT4 i1_3_lut (.I0(\PID_CONTROLLER.result [22]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n4_adj_3416));   // verilog/motorControl.v(37[31:51])
    defparam i1_3_lut.LUT_INIT = 16'h7e7e;
    SB_CARRY mult_14_add_1217_20 (.CI(n38815), .I0(n1803[17]), .I1(GND_net), 
            .CO(n38816));
    SB_CARRY add_3108_8 (.CI(n38545), .I0(n8475[5]), .I1(n545), .CO(n38546));
    SB_LUT4 add_3149_19_lut (.I0(GND_net), .I1(n10121[16]), .I2(GND_net), 
            .I3(n38116), .O(n9330[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_19 (.CI(n38116), .I0(n10121[16]), .I1(GND_net), 
            .CO(n38117));
    SB_LUT4 add_3108_7_lut (.I0(GND_net), .I1(n8475[4]), .I2(n472), .I3(n38544), 
            .O(n8451[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_18_lut (.I0(GND_net), .I1(n10121[15]), .I2(GND_net), 
            .I3(n38115), .O(n9330[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_18 (.CI(n38115), .I0(n10121[15]), .I1(GND_net), 
            .CO(n38116));
    SB_LUT4 mult_14_add_1217_19_lut (.I0(GND_net), .I1(n1803[16]), .I2(GND_net), 
            .I3(n38814), .O(n1802[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_7 (.CI(n38544), .I0(n8475[4]), .I1(n472), .CO(n38545));
    SB_LUT4 i6_4_lut (.I0(\PID_CONTROLLER.result [13]), .I1(\PID_CONTROLLER.result [23]), 
            .I2(n4_adj_3416), .I3(pwm_23__N_2951[10]), .O(n25_adj_3417));   // verilog/motorControl.v(37[31:51])
    defparam i6_4_lut.LUT_INIT = 16'hf7fe;
    SB_LUT4 add_3149_17_lut (.I0(GND_net), .I1(n10121[14]), .I2(GND_net), 
            .I3(n38114), .O(n9330[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_17 (.CI(n38114), .I0(n10121[14]), .I1(GND_net), 
            .CO(n38115));
    SB_LUT4 add_3108_6_lut (.I0(GND_net), .I1(n8475[3]), .I2(n399), .I3(n38543), 
            .O(n8451[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_16_lut (.I0(GND_net), .I1(n10121[13]), .I2(GND_net), 
            .I3(n38113), .O(n9330[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_31_lut (.I0(GND_net), .I1(n7763[28]), .I2(GND_net), 
            .I3(n37599), .O(n6545[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_16 (.CI(n38113), .I0(n10121[13]), .I1(GND_net), 
            .CO(n38114));
    SB_LUT4 i3_3_lut (.I0(\PID_CONTROLLER.result [15]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n22_c));   // verilog/motorControl.v(37[31:51])
    defparam i3_3_lut.LUT_INIT = 16'h7e7e;
    SB_CARRY mult_14_add_1217_19 (.CI(n38814), .I0(n1803[16]), .I1(GND_net), 
            .CO(n38815));
    SB_CARRY add_3108_6 (.CI(n38543), .I0(n8475[3]), .I1(n399), .CO(n38544));
    SB_LUT4 add_3149_15_lut (.I0(GND_net), .I1(n10121[12]), .I2(GND_net), 
            .I3(n38112), .O(n9330[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_30_lut (.I0(GND_net), .I1(n7763[27]), .I2(GND_net), 
            .I3(n37598), .O(n6545[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_30 (.CI(n37598), .I0(n7763[27]), .I1(GND_net), .CO(n37599));
    SB_CARRY add_3149_15 (.CI(n38112), .I0(n10121[12]), .I1(GND_net), 
            .CO(n38113));
    SB_LUT4 add_3108_5_lut (.I0(GND_net), .I1(n8475[2]), .I2(n326), .I3(n38542), 
            .O(n8451[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_14_lut (.I0(GND_net), .I1(n10121[11]), .I2(GND_net), 
            .I3(n38111), .O(n9330[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_29_lut (.I0(GND_net), .I1(n7763[26]), .I2(GND_net), 
            .I3(n37597), .O(n6545[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_29 (.CI(n37597), .I0(n7763[26]), .I1(GND_net), .CO(n37598));
    SB_CARRY add_3149_14 (.CI(n38111), .I0(n10121[11]), .I1(GND_net), 
            .CO(n38112));
    SB_LUT4 i11_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(n22_c), .I2(\PID_CONTROLLER.result [11]), 
            .I3(pwm_23__N_2951[10]), .O(n30_c));   // verilog/motorControl.v(37[31:51])
    defparam i11_4_lut.LUT_INIT = 16'hdffe;
    SB_LUT4 mult_14_add_1217_18_lut (.I0(GND_net), .I1(n1803[15]), .I2(GND_net), 
            .I3(n38813), .O(n1802[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_5 (.CI(n38542), .I0(n8475[2]), .I1(n326), .CO(n38543));
    SB_LUT4 add_3149_13_lut (.I0(GND_net), .I1(n10121[10]), .I2(GND_net), 
            .I3(n38110), .O(n9330[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_28_lut (.I0(GND_net), .I1(n7763[25]), .I2(GND_net), 
            .I3(n37596), .O(n6545[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_28 (.CI(n37596), .I0(n7763[25]), .I1(GND_net), .CO(n37597));
    SB_CARRY add_3149_13 (.CI(n38110), .I0(n10121[10]), .I1(GND_net), 
            .CO(n38111));
    SB_LUT4 add_3108_4_lut (.I0(GND_net), .I1(n8475[1]), .I2(n253), .I3(n38541), 
            .O(n8451[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_12_lut (.I0(GND_net), .I1(n10121[9]), .I2(GND_net), 
            .I3(n38109), .O(n9330[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_27_lut (.I0(GND_net), .I1(n7763[24]), .I2(GND_net), 
            .I3(n37595), .O(n6545[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_27 (.CI(n37595), .I0(n7763[24]), .I1(GND_net), .CO(n37596));
    SB_CARRY add_3149_12 (.CI(n38109), .I0(n10121[9]), .I1(GND_net), .CO(n38110));
    SB_CARRY mult_14_add_1217_18 (.CI(n38813), .I0(n1803[15]), .I1(GND_net), 
            .CO(n38814));
    SB_CARRY add_3108_4 (.CI(n38541), .I0(n8475[1]), .I1(n253), .CO(n38542));
    SB_LUT4 add_3149_11_lut (.I0(GND_net), .I1(n10121[8]), .I2(GND_net), 
            .I3(n38108), .O(n9330[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_26_lut (.I0(GND_net), .I1(n7763[23]), .I2(GND_net), 
            .I3(n37594), .O(n6545[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_26 (.CI(n37594), .I0(n7763[23]), .I1(GND_net), .CO(n37595));
    SB_CARRY add_3149_11 (.CI(n38108), .I0(n10121[8]), .I1(GND_net), .CO(n38109));
    SB_LUT4 add_3108_3_lut (.I0(GND_net), .I1(n8475[0]), .I2(n180), .I3(n38540), 
            .O(n8451[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_10_lut (.I0(GND_net), .I1(n10121[7]), .I2(GND_net), 
            .I3(n38107), .O(n9330[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_25_lut (.I0(GND_net), .I1(n7763[22]), .I2(GND_net), 
            .I3(n37593), .O(n6545[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_25 (.CI(n37593), .I0(n7763[22]), .I1(GND_net), .CO(n37594));
    SB_CARRY add_3149_10 (.CI(n38107), .I0(n10121[7]), .I1(GND_net), .CO(n38108));
    SB_LUT4 mult_14_add_1217_17_lut (.I0(GND_net), .I1(n1803[14]), .I2(GND_net), 
            .I3(n38812), .O(n1802[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3108_3 (.CI(n38540), .I0(n8475[0]), .I1(n180), .CO(n38541));
    SB_LUT4 add_3149_9_lut (.I0(GND_net), .I1(n10121[6]), .I2(GND_net), 
            .I3(n38106), .O(n9330[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_24_lut (.I0(GND_net), .I1(n7763[21]), .I2(GND_net), 
            .I3(n37592), .O(n6545[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_24 (.CI(n37592), .I0(n7763[21]), .I1(GND_net), .CO(n37593));
    SB_CARRY add_3149_9 (.CI(n38106), .I0(n10121[6]), .I1(GND_net), .CO(n38107));
    SB_LUT4 add_3108_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n8451[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3108_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_3_lut (.I0(\PID_CONTROLLER.result [30]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n28));   // verilog/motorControl.v(37[31:51])
    defparam i9_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 add_3149_8_lut (.I0(GND_net), .I1(n10121[5]), .I2(n545), .I3(n38105), 
            .O(n9330[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_23_lut (.I0(GND_net), .I1(n7763[20]), .I2(GND_net), 
            .I3(n37591), .O(n6545[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut (.I0(\PID_CONTROLLER.result [25]), .I1(\PID_CONTROLLER.result [18]), 
            .I2(pwm_23__N_2951[10]), .I3(\PID_CONTROLLER.result [26]), .O(n29_adj_3419));   // verilog/motorControl.v(37[31:51])
    defparam i10_4_lut.LUT_INIT = 16'h7ffe;
    SB_CARRY add_3010_23 (.CI(n37591), .I0(n7763[20]), .I1(GND_net), .CO(n37592));
    SB_CARRY add_3149_8 (.CI(n38105), .I0(n10121[5]), .I1(n545), .CO(n38106));
    SB_CARRY mult_14_add_1217_17 (.CI(n38812), .I0(n1803[14]), .I1(GND_net), 
            .CO(n38813));
    SB_CARRY add_3108_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n38540));
    SB_LUT4 add_3149_7_lut (.I0(GND_net), .I1(n10121[4]), .I2(n472), .I3(n38104), 
            .O(n9330[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_22_lut (.I0(GND_net), .I1(n7763[19]), .I2(GND_net), 
            .I3(n37590), .O(n6545[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_22 (.CI(n37590), .I0(n7763[19]), .I1(GND_net), .CO(n37591));
    SB_CARRY add_3149_7 (.CI(n38104), .I0(n10121[4]), .I1(n472), .CO(n38105));
    SB_LUT4 add_3107_8_lut (.I0(GND_net), .I1(n9322[5]), .I2(n752_adj_3420), 
            .I3(n38539), .O(n8442[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_6_lut (.I0(GND_net), .I1(n10121[3]), .I2(n399), .I3(n38103), 
            .O(n9330[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_21_lut (.I0(GND_net), .I1(n7763[18]), .I2(GND_net), 
            .I3(n37589), .O(n6545[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_21 (.CI(n37589), .I0(n7763[18]), .I1(GND_net), .CO(n37590));
    SB_CARRY add_3149_6 (.CI(n38103), .I0(n10121[3]), .I1(n399), .CO(n38104));
    SB_LUT4 i8_3_lut (.I0(\PID_CONTROLLER.result [27]), .I1(\PID_CONTROLLER.result [28]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n27_adj_3421));   // verilog/motorControl.v(37[31:51])
    defparam i8_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 mult_14_add_1217_16_lut (.I0(GND_net), .I1(n1803[13]), .I2(GND_net), 
            .I3(n38811), .O(n1802[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3107_7_lut (.I0(GND_net), .I1(n9322[4]), .I2(n655), .I3(n38538), 
            .O(n8442[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_5_lut (.I0(GND_net), .I1(n10121[2]), .I2(n326), .I3(n38102), 
            .O(n9330[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_20_lut (.I0(GND_net), .I1(n7763[17]), .I2(GND_net), 
            .I3(n37588), .O(n6545[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_20 (.CI(n37588), .I0(n7763[17]), .I1(GND_net), .CO(n37589));
    SB_CARRY add_3149_5 (.CI(n38102), .I0(n10121[2]), .I1(n326), .CO(n38103));
    SB_LUT4 pwm_23__I_816_i5_2_lut (.I0(\PID_CONTROLLER.result [2]), .I1(pwm_23__N_2951[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3422));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32218_4_lut (.I0(n11_adj_10), .I1(n9_adj_3378), .I2(n7), 
            .I3(n5_adj_3422), .O(n47720));
    defparam i32218_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 pwm_23__I_816_i8_3_lut (.I0(pwm_23__N_2951[4]), .I1(pwm_23__N_2951[8]), 
            .I2(n17_c), .I3(GND_net), .O(n8_adj_3424));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm__i23 (.Q(pwm[23]), .C(clk32MHz), .D(n24384));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i22 (.Q(pwm[22]), .C(clk32MHz), .D(n24383));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i21 (.Q(pwm[21]), .C(clk32MHz), .D(n24382));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i20 (.Q(pwm[20]), .C(clk32MHz), .D(n24381));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i19 (.Q(pwm[19]), .C(clk32MHz), .D(n24380));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i18 (.Q(pwm[18]), .C(clk32MHz), .D(n42013));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i17 (.Q(pwm[17]), .C(clk32MHz), .D(n42011));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i16 (.Q(pwm[16]), .C(clk32MHz), .D(n24377));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i15 (.Q(pwm[15]), .C(clk32MHz), .D(n24376));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 pwm_23__I_816_i6_3_lut (.I0(pwm_23__N_2951[2]), .I1(pwm_23__N_2951[3]), 
            .I2(n7), .I3(GND_net), .O(n6_adj_3425));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm__i14 (.Q(pwm[14]), .C(clk32MHz), .D(n24375));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i13 (.Q(pwm[13]), .C(clk32MHz), .D(n24374));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i12 (.Q(pwm[12]), .C(clk32MHz), .D(n24373));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i11 (.Q(pwm[11]), .C(clk32MHz), .D(n24372));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i10 (.Q(pwm[10]), .C(clk32MHz), .D(n24371));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i9 (.Q(pwm[9]), .C(clk32MHz), .D(n24370));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i8 (.Q(pwm[8]), .C(clk32MHz), .D(n24369));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i7 (.Q(pwm[7]), .C(clk32MHz), .D(n24368));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i6 (.Q(pwm[6]), .C(clk32MHz), .D(n24367));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i5 (.Q(pwm[5]), .C(clk32MHz), .D(n24366));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i4 (.Q(pwm[4]), .C(clk32MHz), .D(n24365));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i3 (.Q(pwm[3]), .C(clk32MHz), .D(n24364));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i2 (.Q(pwm[2]), .C(clk32MHz), .D(n24363));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i1 (.Q(pwm[1]), .C(clk32MHz), .D(n24362));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF pwm__i0 (.Q(pwm[0]), .C(clk32MHz), .D(n24358));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 pwm_23__I_816_i16_3_lut (.I0(n8_adj_3424), .I1(pwm_23__N_2951[9]), 
            .I2(n19_c), .I3(GND_net), .O(n16_adj_3426));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31974_4_lut (.I0(n50), .I1(\PID_CONTROLLER.result [26]), .I2(\deadband[9] ), 
            .I3(\PID_CONTROLLER.result [25]), .O(n47123));   // verilog/motorControl.v(37[10:27])
    defparam i31974_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 pwm_23__I_816_i4_3_lut (.I0(n47126), .I1(pwm_23__N_2951[1]), 
            .I2(\PID_CONTROLLER.result [1]), .I3(GND_net), .O(n4_adj_3427));   // verilog/motorControl.v(37[31:51])
    defparam pwm_23__I_816_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33225_3_lut (.I0(n4_adj_3427), .I1(\pwm_23__N_2951[5] ), .I2(n11_adj_10), 
            .I3(GND_net), .O(n48727));   // verilog/motorControl.v(37[31:51])
    defparam i33225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33226_3_lut (.I0(n48727), .I1(\pwm_23__N_2951[6] ), .I2(n13_adj_11), 
            .I3(GND_net), .O(n48728));   // verilog/motorControl.v(37[31:51])
    defparam i33226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut (.I0(\PID_CONTROLLER.result [19]), .I1(\PID_CONTROLLER.result [29]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n24_c));   // verilog/motorControl.v(37[31:51])
    defparam i5_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i13_4_lut (.I0(n25_adj_3417), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [16]), .I3(pwm_23__N_2951[10]), .O(n32));   // verilog/motorControl.v(37[31:51])
    defparam i13_4_lut.LUT_INIT = 16'hbffe;
    SB_LUT4 i17_4_lut (.I0(n27_adj_3421), .I1(n29_adj_3419), .I2(n28), 
            .I3(n30_c), .O(n36));   // verilog/motorControl.v(37[31:51])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut (.I0(\PID_CONTROLLER.result [12]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(pwm_23__N_2951[10]), .I3(GND_net), .O(n23_adj_3429));   // verilog/motorControl.v(37[31:51])
    defparam i4_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i32209_4_lut (.I0(n17_c), .I1(n15_adj_12), .I2(n13_adj_11), 
            .I3(n47720), .O(n47711));
    defparam i32209_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n37025), .I0(GND_net), .I1(n57[9]), 
            .CO(n37026));
    SB_LUT4 add_3149_4_lut (.I0(GND_net), .I1(n10121[1]), .I2(n253), .I3(n38101), 
            .O(n9330[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33577_4_lut (.I0(n16_adj_3426), .I1(n6_adj_3425), .I2(n19_c), 
            .I3(n47708), .O(n49079));   // verilog/motorControl.v(37[31:51])
    defparam i33577_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32651_3_lut (.I0(n48728), .I1(\pwm_23__N_2951[7] ), .I2(n15_adj_12), 
            .I3(GND_net), .O(n48153));   // verilog/motorControl.v(37[31:51])
    defparam i32651_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3107_7 (.CI(n38538), .I0(n9322[4]), .I1(n655), .CO(n38539));
    SB_LUT4 i18_4_lut (.I0(n23_adj_3429), .I1(n36), .I2(n32), .I3(n24_c), 
            .O(n45055));   // verilog/motorControl.v(37[31:51])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_3149_4 (.CI(n38101), .I0(n10121[1]), .I1(n253), .CO(n38102));
    SB_LUT4 i33719_4_lut (.I0(n48153), .I1(n49079), .I2(n19_c), .I3(n47711), 
            .O(n49221));   // verilog/motorControl.v(37[31:51])
    defparam i33719_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32835_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [29]), 
            .I2(\PID_CONTROLLER.result [30]), .I3(\PID_CONTROLLER.result [28]), 
            .O(n48337));
    defparam i32835_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i56_3_lut  (.I0(n47123), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n56_adj_3431));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i56_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i60_4_lut  (.I0(\PID_CONTROLLER.result [28]), 
            .I1(\PID_CONTROLLER.result [30]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [29]), 
            .O(n60));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i60_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 add_3010_19_lut (.I0(GND_net), .I1(n7763[16]), .I2(GND_net), 
            .I3(n37587), .O(n6545[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33685_4_lut (.I0(n49221), .I1(\PID_CONTROLLER.result [31]), 
            .I2(pwm_23__N_2951[10]), .I3(n45055), .O(pwm_23__N_2950));   // verilog/motorControl.v(37[31:51])
    defparam i33685_4_lut.LUT_INIT = 16'hcc8e;
    SB_LUT4 i33267_3_lut (.I0(n60), .I1(n56_adj_3431), .I2(n48337), .I3(GND_net), 
            .O(n48769));   // verilog/motorControl.v(37[10:27])
    defparam i33267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 pwm_23__I_815_4_lut (.I0(n48769), .I1(pwm_23__N_2950), .I2(\deadband[9] ), 
            .I3(\PID_CONTROLLER.result [31]), .O(pwm_23__N_2948));   // verilog/motorControl.v(37[10:51])
    defparam pwm_23__I_815_4_lut.LUT_INIT = 16'hecfe;
    SB_CARRY add_3010_19 (.CI(n37587), .I0(n7763[16]), .I1(GND_net), .CO(n37588));
    SB_LUT4 LessThan_22_i17_2_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n63[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3432));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1410 (.I0(\PID_CONTROLLER.result [28]), .I1(\PID_CONTROLLER.result [30]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(GND_net), .O(n43145));   // verilog/motorControl.v(38[12:27])
    defparam i2_3_lut_adj_1410.LUT_INIT = 16'h8080;
    SB_LUT4 i5_3_lut_adj_1411 (.I0(\PID_CONTROLLER.result [20]), .I1(\PID_CONTROLLER.result [22]), 
            .I2(\PID_CONTROLLER.result [18]), .I3(GND_net), .O(n14_adj_3433));
    defparam i5_3_lut_adj_1411.LUT_INIT = 16'h8080;
    SB_LUT4 i6_4_lut_adj_1412 (.I0(\PID_CONTROLLER.result [23]), .I1(\PID_CONTROLLER.result [25]), 
            .I2(\PID_CONTROLLER.result [24]), .I3(\PID_CONTROLLER.result [19]), 
            .O(n15_adj_3434));
    defparam i6_4_lut_adj_1412.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n15_adj_3434), .I1(\PID_CONTROLLER.result [21]), 
            .I2(n14_adj_3433), .I3(\PID_CONTROLLER.result [17]), .O(n43221));
    defparam i8_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i3_4_lut_adj_1413 (.I0(\PID_CONTROLLER.result [23]), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\PID_CONTROLLER.result [22]), .I3(\PID_CONTROLLER.result [25]), 
            .O(n62_adj_3390));   // verilog/motorControl.v(31[14] 52[8])
    defparam i3_4_lut_adj_1413.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [19]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3435));   // verilog/motorControl.v(31[14] 52[8])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(\PID_CONTROLLER.result [20]), .I1(\PID_CONTROLLER.result [17]), 
            .I2(\PID_CONTROLLER.result [18]), .I3(n6_adj_3435), .O(n49));   // verilog/motorControl.v(31[14] 52[8])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_14_i392_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n583_adj_3436));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i392_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_3437));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i7_2_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n63[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3438));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_22_i9_2_lut (.I0(\PID_CONTROLLER.result [4]), .I1(n63[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3439));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3440));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i19_2_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n63[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_3441));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i146_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n216));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_2_lut (.I0(\PID_CONTROLLER.result [14]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_3442));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1414 (.I0(\PID_CONTROLLER.result [11]), .I1(\PID_CONTROLLER.result [27]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(\PID_CONTROLLER.result [10]), 
            .O(n24_adj_3443));
    defparam i10_4_lut_adj_1414.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_22_i5_2_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n63[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3444));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32159_4_lut (.I0(n11_adj_13), .I1(n9_adj_3439), .I2(n7_adj_3438), 
            .I3(n5_adj_3444), .O(n47660));
    defparam i32159_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i203_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n301_adj_3446));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i93_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n137_adj_3447));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_22_i4_4_lut (.I0(n63[0]), .I1(n63[1]), .I2(\PID_CONTROLLER.result [1]), 
            .I3(\PID_CONTROLLER.result [0]), .O(n4_adj_3448));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i33219_3_lut (.I0(n4_adj_3448), .I1(n415), .I2(n11_adj_13), 
            .I3(GND_net), .O(n48721));   // verilog/motorControl.v(40[21:37])
    defparam i33219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3149_3_lut (.I0(GND_net), .I1(n10121[0]), .I2(n180), .I3(n38100), 
            .O(n9330[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33220_3_lut (.I0(n48721), .I1(n414), .I2(n13_adj_14), .I3(GND_net), 
            .O(n48722));   // verilog/motorControl.v(40[21:37])
    defparam i33220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1415 (.I0(\PID_CONTROLLER.result [27]), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(GND_net), .O(n10_adj_3450));   // verilog/motorControl.v(31[14] 52[8])
    defparam i1_3_lut_adj_1415.LUT_INIT = 16'h8080;
    SB_LUT4 i8_4_lut_adj_1416 (.I0(\PID_CONTROLLER.result [30]), .I1(n49), 
            .I2(\PID_CONTROLLER.result [12]), .I3(\PID_CONTROLLER.result [28]), 
            .O(n22_adj_3451));
    defparam i8_4_lut_adj_1416.LUT_INIT = 16'hfffe;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i211_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n313));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut_adj_1417 (.I0(\PID_CONTROLLER.result [16]), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(GND_net), .O(n12_adj_3452));   // verilog/motorControl.v(31[14] 52[8])
    defparam i3_3_lut_adj_1417.LUT_INIT = 16'h8080;
    SB_LUT4 i7_4_lut (.I0(n63[10]), .I1(\PID_CONTROLLER.result [12]), .I2(\PID_CONTROLLER.result [26]), 
            .I3(n10_adj_3450), .O(n16_adj_3453));   // verilog/motorControl.v(31[14] 52[8])
    defparam i7_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i12_4_lut (.I0(\PID_CONTROLLER.result [29]), .I1(n24_adj_3443), 
            .I2(n18_adj_3442), .I3(n62_adj_3390), .O(n26_adj_3454));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15326_1_lut (.I0(\PID_CONTROLLER.result [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n28729));   // verilog/motorControl.v(31[14] 52[8])
    defparam i15326_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31880_4_lut (.I0(n43221), .I1(n16_adj_3453), .I2(n12_adj_3452), 
            .I3(n43145), .O(n47241));   // verilog/motorControl.v(31[14] 52[8])
    defparam i31880_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3010_18_lut (.I0(GND_net), .I1(n7763[15]), .I2(GND_net), 
            .I3(n37586), .O(n6545[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_3 (.CI(n38100), .I0(n10121[0]), .I1(n180), .CO(n38101));
    SB_LUT4 i11_3_lut (.I0(\PID_CONTROLLER.result [26]), .I1(n22_adj_3451), 
            .I2(n63[10]), .I3(GND_net), .O(n25_adj_3455));
    defparam i11_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 add_3107_6_lut (.I0(GND_net), .I1(n9322[3]), .I2(n558_adj_3456), 
            .I3(n38537), .O(n8442[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_22_i6_3_lut (.I0(n63[2]), .I1(n63[3]), .I2(n7_adj_3438), 
            .I3(GND_net), .O(n6_adj_3457));   // verilog/motorControl.v(40[21:37])
    defparam LessThan_22_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33411_3_lut (.I0(n6_adj_3457), .I1(n63[4]), .I2(n9_adj_3439), 
            .I3(GND_net), .O(n48913));   // verilog/motorControl.v(40[21:37])
    defparam i33411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_17_inv_0_i1_1_lut (.I0(\deadband[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[0]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33412_3_lut (.I0(n48913), .I1(n63[8]), .I2(n17_adj_3432), 
            .I3(GND_net), .O(n48914));   // verilog/motorControl.v(40[21:37])
    defparam i33412_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3010_18 (.CI(n37586), .I0(n7763[15]), .I1(GND_net), .CO(n37587));
    SB_LUT4 add_3010_17_lut (.I0(GND_net), .I1(n7763[14]), .I2(GND_net), 
            .I3(n37585), .O(n6545[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n9330[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_17 (.CI(n37585), .I0(n7763[14]), .I1(GND_net), .CO(n37586));
    SB_LUT4 add_3010_16_lut (.I0(GND_net), .I1(n7763[13]), .I2(GND_net), 
            .I3(n37584), .O(n6545[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_16 (.CI(n38811), .I0(n1803[13]), .I1(GND_net), 
            .CO(n38812));
    SB_CARRY add_3149_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n38100));
    SB_CARRY add_3010_16 (.CI(n37584), .I0(n7763[13]), .I1(GND_net), .CO(n37585));
    SB_LUT4 add_3010_15_lut (.I0(GND_net), .I1(n7763[12]), .I2(GND_net), 
            .I3(n37583), .O(n6545[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_7_lut (.I0(GND_net), .I1(n44998), .I2(n658_adj_3459), 
            .I3(n38099), .O(n9322[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_15 (.CI(n37583), .I0(n7763[12]), .I1(GND_net), .CO(n37584));
    SB_LUT4 add_3010_14_lut (.I0(GND_net), .I1(n7763[11]), .I2(GND_net), 
            .I3(n37582), .O(n6545[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i158_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n234_adj_3460));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1217_15_lut (.I0(GND_net), .I1(n1803[12]), .I2(GND_net), 
            .I3(n38810), .O(n1802[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3107_6 (.CI(n38537), .I0(n9322[3]), .I1(n558_adj_3456), 
            .CO(n38538));
    SB_LUT4 add_3148_6_lut (.I0(GND_net), .I1(n10114[3]), .I2(n564), .I3(n38098), 
            .O(n9322[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_6 (.CI(n38098), .I0(n10114[3]), .I1(n564), .CO(n38099));
    SB_CARRY add_3010_14 (.CI(n37582), .I0(n7763[11]), .I1(GND_net), .CO(n37583));
    SB_LUT4 add_3107_5_lut (.I0(GND_net), .I1(n9322[2]), .I2(n461_adj_3461), 
            .I3(n38536), .O(n8442[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_5_lut (.I0(GND_net), .I1(n10114[2]), .I2(n464_adj_3462), 
            .I3(n38097), .O(n9322[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_5 (.CI(n38097), .I0(n10114[2]), .I1(n464_adj_3462), 
            .CO(n38098));
    SB_LUT4 add_3010_13_lut (.I0(GND_net), .I1(n7763[10]), .I2(GND_net), 
            .I3(n37581), .O(n6545[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_13 (.CI(n37581), .I0(n7763[10]), .I1(GND_net), .CO(n37582));
    SB_CARRY mult_14_add_1217_15 (.CI(n38810), .I0(n1803[12]), .I1(GND_net), 
            .CO(n38811));
    SB_CARRY add_3107_5 (.CI(n38536), .I0(n9322[2]), .I1(n461_adj_3461), 
            .CO(n38537));
    SB_LUT4 add_3148_4_lut (.I0(GND_net), .I1(n11529[1]), .I2(n370_adj_3463), 
            .I3(n38096), .O(n9322[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_4 (.CI(n38096), .I0(n11529[1]), .I1(n370_adj_3463), 
            .CO(n38097));
    SB_LUT4 add_3010_12_lut (.I0(GND_net), .I1(n7763[9]), .I2(GND_net), 
            .I3(n37580), .O(n6545[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_12 (.CI(n37580), .I0(n7763[9]), .I1(GND_net), .CO(n37581));
    SB_LUT4 add_3107_4_lut (.I0(GND_net), .I1(n9322[1]), .I2(n364), .I3(n38535), 
            .O(n8442[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_3_lut (.I0(GND_net), .I1(n10114[0]), .I2(n276_adj_3464), 
            .I3(n38095), .O(n9322[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_3 (.CI(n38095), .I0(n10114[0]), .I1(n276_adj_3464), 
            .CO(n38096));
    SB_LUT4 add_3010_11_lut (.I0(GND_net), .I1(n7763[8]), .I2(GND_net), 
            .I3(n37579), .O(n6545[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_11 (.CI(n37579), .I0(n7763[8]), .I1(GND_net), .CO(n37580));
    SB_LUT4 mult_14_add_1217_14_lut (.I0(GND_net), .I1(n1803[11]), .I2(GND_net), 
            .I3(n38809), .O(n1802[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_2_lut (.I0(GND_net), .I1(n86_adj_3465), .I2(n182_adj_3466), 
            .I3(GND_net), .O(n9322[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3107_4 (.CI(n38535), .I0(n9322[1]), .I1(n364), .CO(n38536));
    SB_CARRY add_3148_2 (.CI(GND_net), .I0(n86_adj_3465), .I1(n182_adj_3466), 
            .CO(n38095));
    SB_CARRY mult_14_add_1217_14 (.CI(n38809), .I0(n1803[11]), .I1(GND_net), 
            .CO(n38810));
    SB_DFF \PID_CONTROLLER.result_i0  (.Q(\PID_CONTROLLER.result [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [0]));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3198_10 (.CI(n37436), .I0(n11361[7]), .I1(GND_net), .CO(n37437));
    SB_LUT4 i32134_4_lut (.I0(n17_adj_3432), .I1(n15_adj_15), .I2(n13_adj_14), 
            .I3(n47660), .O(n47635));
    defparam i32134_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3178_20_lut (.I0(GND_net), .I1(n10855[17]), .I2(GND_net), 
            .I3(n38094), .O(n10121[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err[0] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [0]));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3178_19_lut (.I0(GND_net), .I1(n10855[16]), .I2(GND_net), 
            .I3(n38093), .O(n10121[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_19_lut.LUT_INIT = 16'hC33C;
    SB_DFFE PHASES_i2 (.Q(PIN_7_c_1), .C(clk32MHz), .E(n23569), .D(PHASES_5__N_2779[1]));   // verilog/motorControl.v(57[10] 100[6])
    SB_LUT4 i32661_3_lut (.I0(n48722), .I1(n413), .I2(n15_adj_15), .I3(GND_net), 
            .O(n48163));   // verilog/motorControl.v(40[21:37])
    defparam i32661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3010_10_lut (.I0(GND_net), .I1(n7763[7]), .I2(GND_net), 
            .I3(n37578), .O(n6545[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_10 (.CI(n37578), .I0(n7763[7]), .I1(GND_net), .CO(n37579));
    SB_LUT4 add_3107_3_lut (.I0(GND_net), .I1(n9322[0]), .I2(n267), .I3(n38534), 
            .O(n8442[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_19 (.CI(n38093), .I0(n10855[16]), .I1(GND_net), 
            .CO(n38094));
    SB_LUT4 add_3178_18_lut (.I0(GND_net), .I1(n10855[15]), .I2(GND_net), 
            .I3(n38092), .O(n10121[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_9_lut (.I0(GND_net), .I1(n7763[6]), .I2(GND_net), 
            .I3(n37577), .O(n6545[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_9 (.CI(n37577), .I0(n7763[6]), .I1(GND_net), .CO(n37578));
    SB_LUT4 mult_14_add_1217_13_lut (.I0(GND_net), .I1(n1803[10]), .I2(GND_net), 
            .I3(n38808), .O(n1802[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33368_3_lut (.I0(n48914), .I1(n63[9]), .I2(n19_adj_3441), 
            .I3(GND_net), .O(n48591));   // verilog/motorControl.v(40[21:37])
    defparam i33368_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3107_3 (.CI(n38534), .I0(n9322[0]), .I1(n267), .CO(n38535));
    SB_CARRY add_3178_18 (.CI(n38092), .I0(n10855[15]), .I1(GND_net), 
            .CO(n38093));
    SB_LUT4 add_3178_17_lut (.I0(GND_net), .I1(n10855[14]), .I2(GND_net), 
            .I3(n38091), .O(n10121[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_8_lut (.I0(GND_net), .I1(n7763[5]), .I2(n683_adj_3468), 
            .I3(n37576), .O(n6545[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_13 (.CI(n38808), .I0(n1803[10]), .I1(GND_net), 
            .CO(n38809));
    SB_LUT4 mult_10_i276_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n410_adj_3469));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i276_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3010_8 (.CI(n37576), .I0(n7763[5]), .I1(n683_adj_3468), 
            .CO(n37577));
    SB_LUT4 add_3107_2_lut (.I0(GND_net), .I1(n86_adj_3465), .I2(n170), 
            .I3(GND_net), .O(n8442[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3107_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_17 (.CI(n38091), .I0(n10855[14]), .I1(GND_net), 
            .CO(n38092));
    SB_LUT4 i28_4_lut (.I0(n25_adj_3455), .I1(n47241), .I2(\PID_CONTROLLER.result [13]), 
            .I3(n26_adj_3454), .O(n20_adj_3470));   // verilog/motorControl.v(31[14] 52[8])
    defparam i28_4_lut.LUT_INIT = 16'hc0c5;
    SB_LUT4 add_3178_16_lut (.I0(GND_net), .I1(n10855[13]), .I2(GND_net), 
            .I3(n38090), .O(n10121[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_7_lut (.I0(GND_net), .I1(n7763[4]), .I2(n586), .I3(n37575), 
            .O(n6545[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_12_lut (.I0(GND_net), .I1(n1803[9]), .I2(GND_net), 
            .I3(n38807), .O(n1802[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_7 (.CI(n37575), .I0(n7763[4]), .I1(n586), .CO(n37576));
    SB_LUT4 i33273_4_lut (.I0(n48591), .I1(n48163), .I2(n19_adj_3441), 
            .I3(n47635), .O(n48775));   // verilog/motorControl.v(40[21:37])
    defparam i33273_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i33057_4_lut (.I0(n48775), .I1(\PID_CONTROLLER.result [31]), 
            .I2(n63[10]), .I3(n20_adj_3470), .O(n421));   // verilog/motorControl.v(40[21:37])
    defparam i33057_4_lut.LUT_INIT = 16'h8ecc;
    SB_CARRY mult_14_add_1217_12 (.CI(n38807), .I0(n1803[9]), .I1(GND_net), 
            .CO(n38808));
    SB_CARRY add_3107_2 (.CI(GND_net), .I0(n86_adj_3465), .I1(n170), .CO(n38534));
    SB_LUT4 mult_10_i223_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n331));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3106_9_lut (.I0(GND_net), .I1(n8442[6]), .I2(GND_net), 
            .I3(n38533), .O(n8432[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_16 (.CI(n38090), .I0(n10855[13]), .I1(GND_net), 
            .CO(n38091));
    SB_LUT4 add_3178_15_lut (.I0(GND_net), .I1(n10855[12]), .I2(GND_net), 
            .I3(n38089), .O(n10121[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3010_6_lut (.I0(GND_net), .I1(n7763[3]), .I2(n489), .I3(n37574), 
            .O(n6545[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_6 (.CI(n37574), .I0(n7763[3]), .I1(n489), .CO(n37575));
    SB_LUT4 add_3010_5_lut (.I0(GND_net), .I1(n7763[2]), .I2(n392), .I3(n37573), 
            .O(n6545[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3106_8_lut (.I0(GND_net), .I1(n8442[5]), .I2(n749), .I3(n38532), 
            .O(n8432[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_15 (.CI(n38089), .I0(n10855[12]), .I1(GND_net), 
            .CO(n38090));
    SB_LUT4 add_3178_14_lut (.I0(GND_net), .I1(n10855[11]), .I2(GND_net), 
            .I3(n38088), .O(n10121[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_5 (.CI(n37573), .I0(n7763[2]), .I1(n392), .CO(n37574));
    SB_LUT4 mult_14_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i341_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n507));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i341_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3178_14 (.CI(n38088), .I0(n10855[11]), .I1(GND_net), 
            .CO(n38089));
    SB_LUT4 add_3010_4_lut (.I0(GND_net), .I1(n7763[1]), .I2(n295), .I3(n37572), 
            .O(n6545[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_4 (.CI(n37572), .I0(n7763[1]), .I1(n295), .CO(n37573));
    SB_LUT4 mult_14_add_1217_11_lut (.I0(GND_net), .I1(n1803[8]), .I2(GND_net), 
            .I3(n38806), .O(n1802[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_8 (.CI(n38532), .I0(n8442[5]), .I1(n749), .CO(n38533));
    SB_LUT4 add_3178_13_lut (.I0(GND_net), .I1(n10855[10]), .I2(GND_net), 
            .I3(n38087), .O(n10121[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_13 (.CI(n38087), .I0(n10855[10]), .I1(GND_net), 
            .CO(n38088));
    SB_LUT4 add_3010_3_lut (.I0(GND_net), .I1(n7763[0]), .I2(n198), .I3(n37571), 
            .O(n6545[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_3 (.CI(n37571), .I0(n7763[0]), .I1(n198), .CO(n37572));
    SB_LUT4 add_3106_7_lut (.I0(GND_net), .I1(n8442[4]), .I2(n652), .I3(n38531), 
            .O(n8432[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_12_lut (.I0(GND_net), .I1(n10855[9]), .I2(GND_net), 
            .I3(n38086), .O(n10121[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_12 (.CI(n38086), .I0(n10855[9]), .I1(GND_net), .CO(n38087));
    SB_LUT4 add_3010_2_lut (.I0(GND_net), .I1(n8_adj_3471), .I2(n101), 
            .I3(GND_net), .O(n6545[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3010_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3010_2 (.CI(GND_net), .I0(n8_adj_3471), .I1(n101), .CO(n37571));
    SB_CARRY mult_14_add_1217_11 (.CI(n38806), .I0(n1803[8]), .I1(GND_net), 
            .CO(n38807));
    SB_CARRY add_3106_7 (.CI(n38531), .I0(n8442[4]), .I1(n652), .CO(n38532));
    SB_LUT4 add_3178_11_lut (.I0(GND_net), .I1(n10855[8]), .I2(GND_net), 
            .I3(n38085), .O(n10121[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_11 (.CI(n38085), .I0(n10855[8]), .I1(GND_net), .CO(n38086));
    SB_LUT4 add_3077_30_lut (.I0(GND_net), .I1(n9128[27]), .I2(GND_net), 
            .I3(n37570), .O(n7763[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_29_lut (.I0(GND_net), .I1(n9128[26]), .I2(GND_net), 
            .I3(n37569), .O(n7763[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3106_6_lut (.I0(GND_net), .I1(n8442[3]), .I2(n555), .I3(n38530), 
            .O(n8432[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_10_lut (.I0(GND_net), .I1(n10855[7]), .I2(GND_net), 
            .I3(n38084), .O(n10121[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_10 (.CI(n38084), .I0(n10855[7]), .I1(GND_net), .CO(n38085));
    SB_CARRY add_3077_29 (.CI(n37569), .I0(n9128[26]), .I1(GND_net), .CO(n37570));
    SB_LUT4 add_3077_28_lut (.I0(GND_net), .I1(n9128[25]), .I2(GND_net), 
            .I3(n37568), .O(n7763[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_10_lut (.I0(GND_net), .I1(n1803[7]), .I2(GND_net), 
            .I3(n38805), .O(n1802[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_6 (.CI(n38530), .I0(n8442[3]), .I1(n555), .CO(n38531));
    SB_LUT4 add_3178_9_lut (.I0(GND_net), .I1(n10855[6]), .I2(GND_net), 
            .I3(n38083), .O(n10121[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_9 (.CI(n38083), .I0(n10855[6]), .I1(GND_net), .CO(n38084));
    SB_CARRY add_3077_28 (.CI(n37568), .I0(n9128[25]), .I1(GND_net), .CO(n37569));
    SB_LUT4 add_3077_27_lut (.I0(GND_net), .I1(n9128[24]), .I2(GND_net), 
            .I3(n37567), .O(n7763[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3106_5_lut (.I0(GND_net), .I1(n8442[2]), .I2(n458_c), 
            .I3(n38529), .O(n8432[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_8_lut (.I0(GND_net), .I1(n10855[5]), .I2(n545), .I3(n38082), 
            .O(n10121[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_8 (.CI(n38082), .I0(n10855[5]), .I1(n545), .CO(n38083));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n57[8]), .I3(n37024), .O(n17_adj_3472)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3077_27 (.CI(n37567), .I0(n9128[24]), .I1(GND_net), .CO(n37568));
    SB_LUT4 add_3077_26_lut (.I0(GND_net), .I1(n9128[23]), .I2(GND_net), 
            .I3(n37566), .O(n7763[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n604));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1217_10 (.CI(n38805), .I0(n1803[7]), .I1(GND_net), 
            .CO(n38806));
    SB_LUT4 add_3178_7_lut (.I0(GND_net), .I1(n10855[4]), .I2(n472), .I3(n38081), 
            .O(n10121[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_7 (.CI(n38081), .I0(n10855[4]), .I1(n472), .CO(n38082));
    SB_LUT4 mult_14_add_1217_9_lut (.I0(GND_net), .I1(n1803[6]), .I2(GND_net), 
            .I3(n38804), .O(n1802[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i268_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n398_adj_3475));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3178_6_lut (.I0(GND_net), .I1(n10855[3]), .I2(n399), .I3(n38080), 
            .O(n10121[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_6 (.CI(n38080), .I0(n10855[3]), .I1(n399), .CO(n38081));
    SB_CARRY add_3077_26 (.CI(n37566), .I0(n9128[23]), .I1(GND_net), .CO(n37567));
    SB_CARRY mult_14_add_1217_9 (.CI(n38804), .I0(n1803[6]), .I1(GND_net), 
            .CO(n38805));
    SB_CARRY add_3106_5 (.CI(n38529), .I0(n8442[2]), .I1(n458_c), .CO(n38530));
    SB_LUT4 add_3178_5_lut (.I0(GND_net), .I1(n10855[2]), .I2(n326), .I3(n38079), 
            .O(n10121[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_5 (.CI(n38079), .I0(n10855[2]), .I1(n326), .CO(n38080));
    SB_LUT4 mult_14_add_1217_8_lut (.I0(GND_net), .I1(n1803[5]), .I2(n530), 
            .I3(n38803), .O(n1802[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_4_lut (.I0(GND_net), .I1(n10855[1]), .I2(n253), .I3(n38078), 
            .O(n10121[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_4 (.CI(n38078), .I0(n10855[1]), .I1(n253), .CO(n38079));
    SB_CARRY mult_14_add_1217_8 (.CI(n38803), .I0(n1803[5]), .I1(n530), 
            .CO(n38804));
    SB_LUT4 add_3178_3_lut (.I0(GND_net), .I1(n10855[0]), .I2(n180), .I3(n38077), 
            .O(n10121[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_3 (.CI(n38077), .I0(n10855[0]), .I1(n180), .CO(n38078));
    SB_LUT4 mult_14_add_1217_7_lut (.I0(GND_net), .I1(n1803[4]), .I2(n457_c), 
            .I3(n38802), .O(n1802[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3178_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n10121[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3178_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3178_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n38077));
    SB_CARRY mult_14_add_1217_7 (.CI(n38802), .I0(n1803[4]), .I1(n457_c), 
            .CO(n38803));
    SB_LUT4 add_3206_19_lut (.I0(GND_net), .I1(n11534[16]), .I2(GND_net), 
            .I3(n38076), .O(n10855[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_18_lut (.I0(GND_net), .I1(n11534[15]), .I2(GND_net), 
            .I3(n38075), .O(n10855[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1217_6_lut (.I0(GND_net), .I1(n1803[3]), .I2(n384), 
            .I3(n38801), .O(n1802[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_18 (.CI(n38075), .I0(n11534[15]), .I1(GND_net), 
            .CO(n38076));
    SB_LUT4 add_3206_17_lut (.I0(GND_net), .I1(n11534[14]), .I2(GND_net), 
            .I3(n38074), .O(n10855[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_25_lut (.I0(GND_net), .I1(n9128[22]), .I2(GND_net), 
            .I3(n37565), .O(n7763[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_6 (.CI(n38801), .I0(n1803[3]), .I1(n384), 
            .CO(n38802));
    SB_LUT4 add_3106_4_lut (.I0(GND_net), .I1(n8442[1]), .I2(n361), .I3(n38528), 
            .O(n8432[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_17 (.CI(n38074), .I0(n11534[14]), .I1(GND_net), 
            .CO(n38075));
    SB_LUT4 add_3198_9_lut (.I0(GND_net), .I1(n11361[6]), .I2(GND_net), 
            .I3(n37435), .O(n10674[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_9 (.CI(n37435), .I0(n11361[6]), .I1(GND_net), .CO(n37436));
    SB_CARRY add_3106_4 (.CI(n38528), .I0(n8442[1]), .I1(n361), .CO(n38529));
    SB_LUT4 add_3206_16_lut (.I0(GND_net), .I1(n11534[13]), .I2(GND_net), 
            .I3(n38073), .O(n10855[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_8_lut (.I0(GND_net), .I1(n11361[5]), .I2(n695), .I3(n37434), 
            .O(n10674[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_8 (.CI(n37434), .I0(n11361[5]), .I1(n695), .CO(n37435));
    SB_LUT4 mult_14_add_1217_5_lut (.I0(GND_net), .I1(n1803[2]), .I2(n311), 
            .I3(n38800), .O(n1802[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_5 (.CI(n38800), .I0(n1803[2]), .I1(n311), 
            .CO(n38801));
    SB_LUT4 add_3106_3_lut (.I0(GND_net), .I1(n8442[0]), .I2(n264), .I3(n38527), 
            .O(n8432[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_16 (.CI(n38073), .I0(n11534[13]), .I1(GND_net), 
            .CO(n38074));
    SB_LUT4 add_3198_7_lut (.I0(GND_net), .I1(n11361[4]), .I2(n598), .I3(n37433), 
            .O(n10674[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_3 (.CI(n38527), .I0(n8442[0]), .I1(n264), .CO(n38528));
    SB_CARRY add_3198_7 (.CI(n37433), .I0(n11361[4]), .I1(n598), .CO(n37434));
    SB_LUT4 add_3206_15_lut (.I0(GND_net), .I1(n11534[12]), .I2(GND_net), 
            .I3(n38072), .O(n10855[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3106_2_lut (.I0(GND_net), .I1(n74), .I2(n167), .I3(GND_net), 
            .O(n8432[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_15 (.CI(n38072), .I0(n11534[12]), .I1(GND_net), 
            .CO(n38073));
    SB_LUT4 add_3206_14_lut (.I0(GND_net), .I1(n11534[11]), .I2(GND_net), 
            .I3(n38071), .O(n10855[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_6_lut (.I0(GND_net), .I1(n11361[3]), .I2(n501_adj_3477), 
            .I3(n37432), .O(n10674[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_6 (.CI(n37432), .I0(n11361[3]), .I1(n501_adj_3477), 
            .CO(n37433));
    SB_CARRY add_3206_14 (.CI(n38071), .I0(n11534[11]), .I1(GND_net), 
            .CO(n38072));
    SB_LUT4 mult_14_add_1217_4_lut (.I0(GND_net), .I1(n1803[1]), .I2(n238_adj_3479), 
            .I3(n38799), .O(n1802[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3106_2 (.CI(GND_net), .I0(n74), .I1(n167), .CO(n38527));
    SB_LUT4 add_3105_10_lut (.I0(GND_net), .I1(n8432[7]), .I2(GND_net), 
            .I3(n38526), .O(n8421[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_13_lut (.I0(GND_net), .I1(n11534[10]), .I2(GND_net), 
            .I3(n38070), .O(n10855[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_9_lut (.I0(GND_net), .I1(n8432[6]), .I2(GND_net), 
            .I3(n38525), .O(n8421[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_5_lut (.I0(GND_net), .I1(n11361[2]), .I2(n404_adj_3480), 
            .I3(n37431), .O(n10674[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_5 (.CI(n37431), .I0(n11361[2]), .I1(n404_adj_3480), 
            .CO(n37432));
    SB_CARRY add_3206_13 (.CI(n38070), .I0(n11534[10]), .I1(GND_net), 
            .CO(n38071));
    SB_CARRY add_3105_9 (.CI(n38525), .I0(n8432[6]), .I1(GND_net), .CO(n38526));
    SB_LUT4 add_3206_12_lut (.I0(GND_net), .I1(n11534[9]), .I2(GND_net), 
            .I3(n38069), .O(n10855[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_12 (.CI(n38069), .I0(n11534[9]), .I1(GND_net), .CO(n38070));
    SB_LUT4 add_3198_4_lut (.I0(GND_net), .I1(n11361[1]), .I2(n307_adj_3481), 
            .I3(n37430), .O(n10674[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_4 (.CI(n37430), .I0(n11361[1]), .I1(n307_adj_3481), 
            .CO(n37431));
    SB_CARRY mult_14_add_1217_4 (.CI(n38799), .I0(n1803[1]), .I1(n238_adj_3479), 
            .CO(n38800));
    SB_LUT4 add_3105_8_lut (.I0(GND_net), .I1(n8432[5]), .I2(n746_adj_3482), 
            .I3(n38524), .O(n8421[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_11_lut (.I0(GND_net), .I1(n11534[8]), .I2(GND_net), 
            .I3(n38068), .O(n10855[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_11 (.CI(n38068), .I0(n11534[8]), .I1(GND_net), .CO(n38069));
    SB_LUT4 add_3198_3_lut (.I0(GND_net), .I1(n11361[0]), .I2(n210_adj_3483), 
            .I3(n37429), .O(n10674[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_3 (.CI(n37429), .I0(n11361[0]), .I1(n210_adj_3483), 
            .CO(n37430));
    SB_CARRY unary_minus_5_add_3_10 (.CI(n37024), .I0(GND_net), .I1(n57[8]), 
            .CO(n37025));
    SB_LUT4 add_22984_33_lut (.I0(GND_net), .I1(n66[31]), .I2(n7064[0]), 
            .I3(n37216), .O(\PID_CONTROLLER.result_31__N_2994 [31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_8 (.CI(n38524), .I0(n8432[5]), .I1(n746_adj_3482), 
            .CO(n38525));
    SB_LUT4 add_3206_10_lut (.I0(GND_net), .I1(n11534[7]), .I2(GND_net), 
            .I3(n38067), .O(n10855[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3198_2_lut (.I0(GND_net), .I1(n20_adj_3484), .I2(n113_adj_3485), 
            .I3(GND_net), .O(n10674[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_32_lut (.I0(GND_net), .I1(n66[30]), .I2(n191[30]), 
            .I3(n37215), .O(\PID_CONTROLLER.result_31__N_2994 [30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_2 (.CI(GND_net), .I0(n20_adj_3484), .I1(n113_adj_3485), 
            .CO(n37429));
    SB_CARRY add_22984_32 (.CI(n37215), .I0(n66[30]), .I1(n191[30]), .CO(n37216));
    SB_LUT4 mult_14_add_1217_3_lut (.I0(GND_net), .I1(n1803[0]), .I2(n165_adj_3486), 
            .I3(n38798), .O(n1802[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_7_lut (.I0(GND_net), .I1(n8432[4]), .I2(n649_adj_3487), 
            .I3(n38523), .O(n8421[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_10 (.CI(n38067), .I0(n11534[7]), .I1(GND_net), .CO(n38068));
    SB_LUT4 add_3370_12_lut (.I0(GND_net), .I1(n14915[9]), .I2(GND_net), 
            .I3(n37428), .O(n14563[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_31_lut (.I0(GND_net), .I1(n66[29]), .I2(n191[29]), 
            .I3(n37214), .O(\PID_CONTROLLER.result_31__N_2994 [29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_11_lut (.I0(GND_net), .I1(n14915[8]), .I2(GND_net), 
            .I3(n37427), .O(n14563[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_31 (.CI(n37214), .I0(n66[29]), .I1(n191[29]), .CO(n37215));
    SB_CARRY add_3105_7 (.CI(n38523), .I0(n8432[4]), .I1(n649_adj_3487), 
            .CO(n38524));
    SB_LUT4 add_3206_9_lut (.I0(GND_net), .I1(n11534[6]), .I2(GND_net), 
            .I3(n38066), .O(n10855[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_11 (.CI(n37427), .I0(n14915[8]), .I1(GND_net), .CO(n37428));
    SB_LUT4 add_22984_30_lut (.I0(GND_net), .I1(n66[28]), .I2(n191[28]), 
            .I3(n37213), .O(\PID_CONTROLLER.result_31__N_2994 [28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n57[7]), .I3(n37023), .O(n15_adj_3488)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3370_10_lut (.I0(GND_net), .I1(n14915[7]), .I2(GND_net), 
            .I3(n37426), .O(n14563[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1217_3 (.CI(n38798), .I0(n1803[0]), .I1(n165_adj_3486), 
            .CO(n38799));
    SB_CARRY add_22984_30 (.CI(n37213), .I0(n66[28]), .I1(n191[28]), .CO(n37214));
    SB_CARRY unary_minus_5_add_3_9 (.CI(n37023), .I0(GND_net), .I1(n57[7]), 
            .CO(n37024));
    SB_LUT4 mult_14_add_1217_2_lut (.I0(GND_net), .I1(n23_adj_3490), .I2(n92), 
            .I3(GND_net), .O(n1802[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1217_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_6_lut (.I0(GND_net), .I1(n8432[3]), .I2(n552_adj_3491), 
            .I3(n38522), .O(n8421[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_6 (.CI(n38522), .I0(n8432[3]), .I1(n552_adj_3491), 
            .CO(n38523));
    SB_CARRY add_3206_9 (.CI(n38066), .I0(n11534[6]), .I1(GND_net), .CO(n38067));
    SB_CARRY add_3370_10 (.CI(n37426), .I0(n14915[7]), .I1(GND_net), .CO(n37427));
    SB_LUT4 add_22984_29_lut (.I0(GND_net), .I1(n66[27]), .I2(n191[27]), 
            .I3(n37212), .O(\PID_CONTROLLER.result_31__N_2994 [27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n57[6]), .I3(n37022), .O(n13_adj_3492)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3206_8_lut (.I0(GND_net), .I1(n11534[5]), .I2(n545), .I3(n38065), 
            .O(n10855[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_29 (.CI(n37212), .I0(n66[27]), .I1(n191[27]), .CO(n37213));
    SB_LUT4 add_3370_9_lut (.I0(GND_net), .I1(n14915[6]), .I2(GND_net), 
            .I3(n37425), .O(n14563[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_28_lut (.I0(GND_net), .I1(n66[26]), .I2(n191[26]), 
            .I3(n37211), .O(\PID_CONTROLLER.result_31__N_2994 [26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n37022), .I0(GND_net), .I1(n57[6]), 
            .CO(n37023));
    SB_CARRY add_22984_28 (.CI(n37211), .I0(n66[26]), .I1(n191[26]), .CO(n37212));
    SB_LUT4 add_3105_5_lut (.I0(GND_net), .I1(n8432[2]), .I2(n455_adj_3494), 
            .I3(n38521), .O(n8421[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_8 (.CI(n38065), .I0(n11534[5]), .I1(n545), .CO(n38066));
    SB_CARRY add_3370_9 (.CI(n37425), .I0(n14915[6]), .I1(GND_net), .CO(n37426));
    SB_CARRY add_3077_25 (.CI(n37565), .I0(n9128[22]), .I1(GND_net), .CO(n37566));
    SB_LUT4 add_22984_27_lut (.I0(GND_net), .I1(n66[25]), .I2(n191[25]), 
            .I3(n37210), .O(\PID_CONTROLLER.result_31__N_2994 [25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n57[5]), .I3(n37021), .O(n11_adj_3495)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n37021), .I0(GND_net), .I1(n57[5]), 
            .CO(n37022));
    SB_CARRY add_22984_27 (.CI(n37210), .I0(n66[25]), .I1(n191[25]), .CO(n37211));
    SB_LUT4 add_3370_8_lut (.I0(GND_net), .I1(n14915[5]), .I2(n545), .I3(n37424), 
            .O(n14563[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_26_lut (.I0(GND_net), .I1(n66[24]), .I2(n191[24]), 
            .I3(n37209), .O(\PID_CONTROLLER.result_31__N_2994 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n57[4]), .I3(n37020), .O(n9_adj_3497)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n37020), .I0(GND_net), .I1(n57[4]), 
            .CO(n37021));
    SB_CARRY add_22984_26 (.CI(n37209), .I0(n66[24]), .I1(n191[24]), .CO(n37210));
    SB_CARRY mult_14_add_1217_2 (.CI(GND_net), .I0(n23_adj_3490), .I1(n92), 
            .CO(n38798));
    SB_CARRY add_3105_5 (.CI(n38521), .I0(n8432[2]), .I1(n455_adj_3494), 
            .CO(n38522));
    SB_LUT4 add_3206_7_lut (.I0(GND_net), .I1(n11534[4]), .I2(n472), .I3(n38064), 
            .O(n10855[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_8 (.CI(n37424), .I0(n14915[5]), .I1(n545), .CO(n37425));
    SB_LUT4 add_22984_25_lut (.I0(GND_net), .I1(n66[23]), .I2(n191[23]), 
            .I3(n37208), .O(\PID_CONTROLLER.result_31__N_2994 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_7_lut (.I0(GND_net), .I1(n14915[4]), .I2(n472), .I3(n37423), 
            .O(n14563[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_25 (.CI(n37208), .I0(n66[23]), .I1(n191[23]), .CO(n37209));
    SB_LUT4 add_3105_4_lut (.I0(GND_net), .I1(n8432[1]), .I2(n358_adj_3499), 
            .I3(n38520), .O(n8421[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_7 (.CI(n38064), .I0(n11534[4]), .I1(n472), .CO(n38065));
    SB_CARRY add_3370_7 (.CI(n37423), .I0(n14915[4]), .I1(n472), .CO(n37424));
    SB_LUT4 add_22984_24_lut (.I0(GND_net), .I1(n66[22]), .I2(n191[22]), 
            .I3(n37207), .O(\PID_CONTROLLER.result_31__N_2994 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n57[3]), .I3(n37019), .O(n7_adj_3500)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_14_add_1216_24_lut (.I0(GND_net), .I1(n1802[21]), .I2(GND_net), 
            .I3(n38796), .O(n1801[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_4 (.CI(n38520), .I0(n8432[1]), .I1(n358_adj_3499), 
            .CO(n38521));
    SB_LUT4 add_3206_6_lut (.I0(GND_net), .I1(n11534[3]), .I2(n399), .I3(n38063), 
            .O(n10855[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_6_lut (.I0(GND_net), .I1(n14915[3]), .I2(n399), .I3(n37422), 
            .O(n14563[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_24 (.CI(n37207), .I0(n66[22]), .I1(n191[22]), .CO(n37208));
    SB_CARRY unary_minus_5_add_3_5 (.CI(n37019), .I0(GND_net), .I1(n57[3]), 
            .CO(n37020));
    SB_LUT4 add_22984_23_lut (.I0(GND_net), .I1(n66[21]), .I2(n191[21]), 
            .I3(n37206), .O(\PID_CONTROLLER.result_31__N_2994 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_6 (.CI(n37422), .I0(n14915[3]), .I1(n399), .CO(n37423));
    SB_CARRY add_22984_23 (.CI(n37206), .I0(n66[21]), .I1(n191[21]), .CO(n37207));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n57[2]), .I3(n37018), .O(n5_adj_3502)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_22984_22_lut (.I0(GND_net), .I1(n66[20]), .I2(n191[20]), 
            .I3(n37205), .O(\PID_CONTROLLER.result_31__N_2994 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_3_lut (.I0(GND_net), .I1(n8432[0]), .I2(n261_adj_3504), 
            .I3(n38519), .O(n8421[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_6 (.CI(n38063), .I0(n11534[3]), .I1(n399), .CO(n38064));
    SB_LUT4 add_3370_5_lut (.I0(GND_net), .I1(n14915[2]), .I2(n326), .I3(n37421), 
            .O(n14563[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_22 (.CI(n37205), .I0(n66[20]), .I1(n191[20]), .CO(n37206));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n37018), .I0(GND_net), .I1(n57[2]), 
            .CO(n37019));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n57[1]), .I3(n37017), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_22984_21_lut (.I0(GND_net), .I1(n66[19]), .I2(n191[19]), 
            .I3(n37204), .O(\PID_CONTROLLER.result_31__N_2994 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3206_5_lut (.I0(GND_net), .I1(n11534[2]), .I2(n326), .I3(n38062), 
            .O(n10855[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_24_lut (.I0(GND_net), .I1(n9128[21]), .I2(GND_net), 
            .I3(n37564), .O(n7763[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1216_24 (.CI(n38796), .I0(n1802[21]), .I1(GND_net), 
            .CO(n1703));
    SB_CARRY add_3105_3 (.CI(n38519), .I0(n8432[0]), .I1(n261_adj_3504), 
            .CO(n38520));
    SB_CARRY add_3206_5 (.CI(n38062), .I0(n11534[2]), .I1(n326), .CO(n38063));
    SB_LUT4 add_3206_4_lut (.I0(GND_net), .I1(n11534[1]), .I2(n253), .I3(n38061), 
            .O(n10855[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3105_2_lut (.I0(GND_net), .I1(n71_adj_3506), .I2(n164_adj_3507), 
            .I3(GND_net), .O(n8421[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3105_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_4 (.CI(n38061), .I0(n11534[1]), .I1(n253), .CO(n38062));
    SB_LUT4 add_3206_3_lut (.I0(GND_net), .I1(n11534[0]), .I2(n180), .I3(n38060), 
            .O(n10855[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_23_lut (.I0(GND_net), .I1(n1802[20]), .I2(GND_net), 
            .I3(n38795), .O(n1801[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3105_2 (.CI(GND_net), .I0(n71_adj_3506), .I1(n164_adj_3507), 
            .CO(n38519));
    SB_CARRY add_3206_3 (.CI(n38060), .I0(n11534[0]), .I1(n180), .CO(n38061));
    SB_CARRY add_3077_24 (.CI(n37564), .I0(n9128[21]), .I1(GND_net), .CO(n37565));
    SB_CARRY add_3370_5 (.CI(n37421), .I0(n14915[2]), .I1(n326), .CO(n37422));
    SB_LUT4 add_3206_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n10855[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3206_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3370_4_lut (.I0(GND_net), .I1(n14915[1]), .I2(n253), .I3(n37420), 
            .O(n14563[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_11_lut (.I0(GND_net), .I1(n8421[8]), .I2(GND_net), 
            .I3(n38518), .O(n8409[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3206_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n38060));
    SB_LUT4 add_3077_23_lut (.I0(GND_net), .I1(n9128[20]), .I2(GND_net), 
            .I3(n37563), .O(n7763[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_18_lut (.I0(GND_net), .I1(n12160[15]), .I2(GND_net), 
            .I3(n38059), .O(n11534[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3370_4 (.CI(n37420), .I0(n14915[1]), .I1(n253), .CO(n37421));
    SB_CARRY add_3077_23 (.CI(n37563), .I0(n9128[20]), .I1(GND_net), .CO(n37564));
    SB_LUT4 add_3077_22_lut (.I0(GND_net), .I1(n9128[19]), .I2(GND_net), 
            .I3(n37562), .O(n7763[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_23 (.CI(n38795), .I0(n1802[20]), .I1(GND_net), 
            .CO(n38796));
    SB_LUT4 add_3370_3_lut (.I0(GND_net), .I1(n14915[0]), .I2(n180), .I3(n37419), 
            .O(n14563[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_17_lut (.I0(GND_net), .I1(n12160[14]), .I2(GND_net), 
            .I3(n38058), .O(n11534[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_10_lut (.I0(GND_net), .I1(n8421[7]), .I2(GND_net), 
            .I3(n38517), .O(n8409[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_17 (.CI(n38058), .I0(n12160[14]), .I1(GND_net), 
            .CO(n38059));
    SB_LUT4 add_3233_16_lut (.I0(GND_net), .I1(n12160[13]), .I2(GND_net), 
            .I3(n38057), .O(n11534[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_16 (.CI(n38057), .I0(n12160[13]), .I1(GND_net), 
            .CO(n38058));
    SB_CARRY add_3104_10 (.CI(n38517), .I0(n8421[7]), .I1(GND_net), .CO(n38518));
    SB_LUT4 mult_10_i288_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n428));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3233_15_lut (.I0(GND_net), .I1(n12160[12]), .I2(GND_net), 
            .I3(n38056), .O(n11534[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_15 (.CI(n38056), .I0(n12160[12]), .I1(GND_net), 
            .CO(n38057));
    SB_CARRY add_22984_21 (.CI(n37204), .I0(n66[19]), .I1(n191[19]), .CO(n37205));
    SB_LUT4 mult_14_add_1216_22_lut (.I0(GND_net), .I1(n1802[19]), .I2(GND_net), 
            .I3(n38794), .O(n1801[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_9_lut (.I0(GND_net), .I1(n8421[6]), .I2(GND_net), 
            .I3(n38516), .O(n8409[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_14_lut (.I0(GND_net), .I1(n12160[11]), .I2(GND_net), 
            .I3(n38055), .O(n11534[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_22 (.CI(n37562), .I0(n9128[19]), .I1(GND_net), .CO(n37563));
    SB_CARRY add_3233_14 (.CI(n38055), .I0(n12160[11]), .I1(GND_net), 
            .CO(n38056));
    SB_CARRY add_3370_3 (.CI(n37419), .I0(n14915[0]), .I1(n180), .CO(n37420));
    SB_CARRY add_3104_9 (.CI(n38516), .I0(n8421[6]), .I1(GND_net), .CO(n38517));
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n701));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3233_13_lut (.I0(GND_net), .I1(n12160[10]), .I2(GND_net), 
            .I3(n38054), .O(n11534[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n525));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3077_21_lut (.I0(GND_net), .I1(n9128[18]), .I2(GND_net), 
            .I3(n37561), .O(n7763[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_13 (.CI(n38054), .I0(n12160[10]), .I1(GND_net), 
            .CO(n38055));
    SB_LUT4 add_3370_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n14563[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3370_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_22 (.CI(n38794), .I0(n1802[19]), .I1(GND_net), 
            .CO(n38795));
    SB_LUT4 add_3104_8_lut (.I0(GND_net), .I1(n8421[5]), .I2(n743), .I3(n38515), 
            .O(n8409[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_12_lut (.I0(GND_net), .I1(n12160[9]), .I2(GND_net), 
            .I3(n38053), .O(n11534[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_12 (.CI(n38053), .I0(n12160[9]), .I1(GND_net), .CO(n38054));
    SB_CARRY add_3104_8 (.CI(n38515), .I0(n8421[5]), .I1(n743), .CO(n38516));
    SB_LUT4 mult_14_add_1216_21_lut (.I0(GND_net), .I1(n1802[18]), .I2(GND_net), 
            .I3(n38793), .O(n1801[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_7_lut (.I0(GND_net), .I1(n8421[4]), .I2(n646), .I3(n38514), 
            .O(n8409[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_11_lut (.I0(GND_net), .I1(n12160[8]), .I2(GND_net), 
            .I3(n38052), .O(n11534[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_21 (.CI(n37561), .I0(n9128[18]), .I1(GND_net), .CO(n37562));
    SB_LUT4 add_22984_20_lut (.I0(GND_net), .I1(n66[18]), .I2(n191[18]), 
            .I3(n37203), .O(\PID_CONTROLLER.result_31__N_2994 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_20_lut (.I0(GND_net), .I1(n9128[17]), .I2(GND_net), 
            .I3(n37560), .O(n7763[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n622));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3077_20 (.CI(n37560), .I0(n9128[17]), .I1(GND_net), .CO(n37561));
    SB_CARRY add_3233_11 (.CI(n38052), .I0(n12160[8]), .I1(GND_net), .CO(n38053));
    SB_CARRY add_3370_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n37419));
    SB_CARRY mult_14_add_1216_21 (.CI(n38793), .I0(n1802[18]), .I1(GND_net), 
            .CO(n38794));
    SB_LUT4 add_3077_19_lut (.I0(GND_net), .I1(n9128[16]), .I2(GND_net), 
            .I3(n37559), .O(n7763[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_10_lut (.I0(GND_net), .I1(n12160[7]), .I2(GND_net), 
            .I3(n38051), .O(n11534[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_10 (.CI(n38051), .I0(n12160[7]), .I1(GND_net), .CO(n38052));
    SB_LUT4 mult_14_add_1216_20_lut (.I0(GND_net), .I1(n1802[17]), .I2(GND_net), 
            .I3(n38792), .O(n1801[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3104_7 (.CI(n38514), .I0(n8421[4]), .I1(n646), .CO(n38515));
    SB_LUT4 add_3233_9_lut (.I0(GND_net), .I1(n12160[6]), .I2(GND_net), 
            .I3(n38050), .O(n11534[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_19 (.CI(n37559), .I0(n9128[16]), .I1(GND_net), .CO(n37560));
    SB_CARRY add_3233_9 (.CI(n38050), .I0(n12160[6]), .I1(GND_net), .CO(n38051));
    SB_LUT4 add_3225_26_lut (.I0(GND_net), .I1(n11995[23]), .I2(GND_net), 
            .I3(n37418), .O(n11361[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_6_lut (.I0(GND_net), .I1(n8421[3]), .I2(n549), .I3(n38513), 
            .O(n8409[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_8_lut (.I0(GND_net), .I1(n12160[5]), .I2(n545), .I3(n38049), 
            .O(n11534[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_18_lut (.I0(GND_net), .I1(n9128[15]), .I2(GND_net), 
            .I3(n37558), .O(n7763[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_8 (.CI(n38049), .I0(n12160[5]), .I1(n545), .CO(n38050));
    SB_CARRY add_3077_18 (.CI(n37558), .I0(n9128[15]), .I1(GND_net), .CO(n37559));
    SB_CARRY add_3104_6 (.CI(n38513), .I0(n8421[3]), .I1(n549), .CO(n38514));
    SB_LUT4 add_3233_7_lut (.I0(GND_net), .I1(n12160[4]), .I2(n472), .I3(n38048), 
            .O(n11534[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_7 (.CI(n38048), .I0(n12160[4]), .I1(n472), .CO(n38049));
    SB_LUT4 add_3225_25_lut (.I0(GND_net), .I1(n11995[22]), .I2(GND_net), 
            .I3(n37417), .O(n11361[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_25 (.CI(n37417), .I0(n11995[22]), .I1(GND_net), 
            .CO(n37418));
    SB_LUT4 add_3104_5_lut (.I0(GND_net), .I1(n8421[2]), .I2(n452), .I3(n38512), 
            .O(n8409[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_20 (.CI(n37203), .I0(n66[18]), .I1(n191[18]), .CO(n37204));
    SB_LUT4 mult_10_i483_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n719));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i483_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n37017), .I0(GND_net), .I1(n57[1]), 
            .CO(n37018));
    SB_CARRY mult_14_add_1216_20 (.CI(n38792), .I0(n1802[17]), .I1(GND_net), 
            .CO(n38793));
    SB_CARRY add_3104_5 (.CI(n38512), .I0(n8421[2]), .I1(n452), .CO(n38513));
    SB_LUT4 add_3233_6_lut (.I0(GND_net), .I1(n12160[3]), .I2(n399), .I3(n38047), 
            .O(n11534[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_6 (.CI(n38047), .I0(n12160[3]), .I1(n399), .CO(n38048));
    SB_LUT4 add_3104_4_lut (.I0(GND_net), .I1(n8421[1]), .I2(n355), .I3(n38511), 
            .O(n8409[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_5_lut (.I0(GND_net), .I1(n12160[2]), .I2(n326), .I3(n38046), 
            .O(n11534[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_5 (.CI(n38046), .I0(n12160[2]), .I1(n326), .CO(n38047));
    SB_LUT4 add_3077_17_lut (.I0(GND_net), .I1(n9128[14]), .I2(GND_net), 
            .I3(n37557), .O(n7763[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_19_lut (.I0(GND_net), .I1(n66[17]), .I2(n191[17]), 
            .I3(n37202), .O(\PID_CONTROLLER.result_31__N_2994 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_19_lut (.I0(GND_net), .I1(n1802[16]), .I2(GND_net), 
            .I3(n38791), .O(n1801[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3104_4 (.CI(n38511), .I0(n8421[1]), .I1(n355), .CO(n38512));
    SB_CARRY add_3077_17 (.CI(n37557), .I0(n9128[14]), .I1(GND_net), .CO(n37558));
    SB_LUT4 add_3233_4_lut (.I0(GND_net), .I1(n12160[1]), .I2(n253), .I3(n38045), 
            .O(n11534[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3233_4 (.CI(n38045), .I0(n12160[1]), .I1(n253), .CO(n38046));
    SB_LUT4 add_3225_24_lut (.I0(GND_net), .I1(n11995[21]), .I2(GND_net), 
            .I3(n37416), .O(n11361[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_3_lut (.I0(GND_net), .I1(n12160[0]), .I2(n180), .I3(n38044), 
            .O(n11534[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_19 (.CI(n38791), .I0(n1802[16]), .I1(GND_net), 
            .CO(n38792));
    SB_LUT4 mult_14_add_1216_18_lut (.I0(GND_net), .I1(n1802[15]), .I2(GND_net), 
            .I3(n38790), .O(n1801[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_19 (.CI(n37202), .I0(n66[17]), .I1(n191[17]), .CO(n37203));
    SB_LUT4 add_3104_3_lut (.I0(GND_net), .I1(n8421[0]), .I2(n258), .I3(n38510), 
            .O(n8409[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3104_3 (.CI(n38510), .I0(n8421[0]), .I1(n258), .CO(n38511));
    SB_LUT4 add_22984_18_lut (.I0(GND_net), .I1(n66[16]), .I2(n191[16]), 
            .I3(n37201), .O(\PID_CONTROLLER.result_31__N_2994 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i95_2_lut (.I0(\Kd[1] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n140_adj_3508));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i32_2_lut (.I0(\Kd[0] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3233_3 (.CI(n38044), .I0(n12160[0]), .I1(n180), .CO(n38045));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n57[0]), 
            .I3(VCC_net), .O(n67[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_24 (.CI(n37416), .I0(n11995[21]), .I1(GND_net), 
            .CO(n37417));
    SB_LUT4 add_3077_16_lut (.I0(GND_net), .I1(n9128[13]), .I2(GND_net), 
            .I3(n37556), .O(n7763[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3233_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n11534[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3233_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_16 (.CI(n37556), .I0(n9128[13]), .I1(GND_net), .CO(n37557));
    SB_CARRY add_3233_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n38044));
    SB_LUT4 add_3077_15_lut (.I0(GND_net), .I1(n9128[12]), .I2(GND_net), 
            .I3(n37555), .O(n7763[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3259_17_lut (.I0(GND_net), .I1(n12735[14]), .I2(GND_net), 
            .I3(n38043), .O(n12160[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_18 (.CI(n38790), .I0(n1802[15]), .I1(GND_net), 
            .CO(n38791));
    SB_LUT4 add_3225_23_lut (.I0(GND_net), .I1(n11995[20]), .I2(GND_net), 
            .I3(n37415), .O(n11361[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3104_2_lut (.I0(GND_net), .I1(n68), .I2(n161), .I3(GND_net), 
            .O(n8409[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3104_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_16_lut (.I0(GND_net), .I1(n12735[13]), .I2(GND_net), 
            .I3(n38042), .O(n12160[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_15 (.CI(n37555), .I0(n9128[12]), .I1(GND_net), .CO(n37556));
    SB_CARRY add_3259_16 (.CI(n38042), .I0(n12735[13]), .I1(GND_net), 
            .CO(n38043));
    SB_CARRY add_3225_23 (.CI(n37415), .I0(n11995[20]), .I1(GND_net), 
            .CO(n37416));
    SB_LUT4 mult_14_add_1216_17_lut (.I0(GND_net), .I1(n1802[14]), .I2(GND_net), 
            .I3(n38789), .O(n1801[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3104_2 (.CI(GND_net), .I0(n68), .I1(n161), .CO(n38510));
    SB_LUT4 add_3259_15_lut (.I0(GND_net), .I1(n12735[12]), .I2(GND_net), 
            .I3(n38041), .O(n12160[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_15 (.CI(n38041), .I0(n12735[12]), .I1(GND_net), 
            .CO(n38042));
    SB_LUT4 add_3103_12_lut (.I0(GND_net), .I1(n8409[9]), .I2(GND_net), 
            .I3(n38509), .O(n8396[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_14_lut (.I0(GND_net), .I1(n12735[11]), .I2(GND_net), 
            .I3(n38040), .O(n12160[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_14 (.CI(n38040), .I0(n12735[11]), .I1(GND_net), 
            .CO(n38041));
    SB_CARRY mult_14_add_1216_17 (.CI(n38789), .I0(n1802[14]), .I1(GND_net), 
            .CO(n38790));
    SB_LUT4 add_3103_11_lut (.I0(GND_net), .I1(n8409[8]), .I2(GND_net), 
            .I3(n38508), .O(n8396[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_13_lut (.I0(GND_net), .I1(n12735[10]), .I2(GND_net), 
            .I3(n38039), .O(n12160[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_14_lut (.I0(GND_net), .I1(n9128[11]), .I2(GND_net), 
            .I3(n37554), .O(n7763[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_13 (.CI(n38039), .I0(n12735[10]), .I1(GND_net), 
            .CO(n38040));
    SB_LUT4 add_3225_22_lut (.I0(GND_net), .I1(n11995[19]), .I2(GND_net), 
            .I3(n37414), .O(n11361[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_11 (.CI(n38508), .I0(n8409[8]), .I1(GND_net), .CO(n38509));
    SB_LUT4 add_3259_12_lut (.I0(GND_net), .I1(n12735[9]), .I2(GND_net), 
            .I3(n38038), .O(n12160[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_14 (.CI(n37554), .I0(n9128[11]), .I1(GND_net), .CO(n37555));
    SB_CARRY add_3259_12 (.CI(n38038), .I0(n12735[9]), .I1(GND_net), .CO(n38039));
    SB_CARRY add_3225_22 (.CI(n37414), .I0(n11995[19]), .I1(GND_net), 
            .CO(n37415));
    SB_LUT4 mult_14_add_1216_16_lut (.I0(GND_net), .I1(n1802[13]), .I2(GND_net), 
            .I3(n38788), .O(n1801[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_10_lut (.I0(GND_net), .I1(n8409[7]), .I2(GND_net), 
            .I3(n38507), .O(n8396[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_11_lut (.I0(GND_net), .I1(n12735[8]), .I2(GND_net), 
            .I3(n38037), .O(n12160[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_11 (.CI(n38037), .I0(n12735[8]), .I1(GND_net), .CO(n38038));
    SB_CARRY add_3103_10 (.CI(n38507), .I0(n8409[7]), .I1(GND_net), .CO(n38508));
    SB_LUT4 add_3259_10_lut (.I0(GND_net), .I1(n12735[7]), .I2(GND_net), 
            .I3(n38036), .O(n12160[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_10 (.CI(n38036), .I0(n12735[7]), .I1(GND_net), .CO(n38037));
    SB_CARRY mult_14_add_1216_16 (.CI(n38788), .I0(n1802[13]), .I1(GND_net), 
            .CO(n38789));
    SB_LUT4 add_3103_9_lut (.I0(GND_net), .I1(n8409[6]), .I2(GND_net), 
            .I3(n38506), .O(n8396[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_9_lut (.I0(GND_net), .I1(n12735[6]), .I2(GND_net), 
            .I3(n38035), .O(n12160[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_13_lut (.I0(GND_net), .I1(n9128[10]), .I2(GND_net), 
            .I3(n37553), .O(n7763[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_9 (.CI(n38035), .I0(n12735[6]), .I1(GND_net), .CO(n38036));
    SB_LUT4 add_3225_21_lut (.I0(GND_net), .I1(n11995[18]), .I2(GND_net), 
            .I3(n37413), .O(n11361[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_9 (.CI(n38506), .I0(n8409[6]), .I1(GND_net), .CO(n38507));
    SB_LUT4 add_3259_8_lut (.I0(GND_net), .I1(n12735[5]), .I2(n545), .I3(n38034), 
            .O(n12160[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_13 (.CI(n37553), .I0(n9128[10]), .I1(GND_net), .CO(n37554));
    SB_CARRY add_3259_8 (.CI(n38034), .I0(n12735[5]), .I1(n545), .CO(n38035));
    SB_CARRY add_3225_21 (.CI(n37413), .I0(n11995[18]), .I1(GND_net), 
            .CO(n37414));
    SB_LUT4 mult_14_add_1216_15_lut (.I0(GND_net), .I1(n1802[12]), .I2(GND_net), 
            .I3(n38787), .O(n1801[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_8_lut (.I0(GND_net), .I1(n8409[5]), .I2(n740), .I3(n38505), 
            .O(n8396[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_7_lut (.I0(GND_net), .I1(n12735[4]), .I2(n472), .I3(n38033), 
            .O(n12160[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_7 (.CI(n38033), .I0(n12735[4]), .I1(n472), .CO(n38034));
    SB_CARRY add_3103_8 (.CI(n38505), .I0(n8409[5]), .I1(n740), .CO(n38506));
    SB_LUT4 add_3259_6_lut (.I0(GND_net), .I1(n12735[3]), .I2(n399), .I3(n38032), 
            .O(n12160[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_6 (.CI(n38032), .I0(n12735[3]), .I1(n399), .CO(n38033));
    SB_CARRY mult_14_add_1216_15 (.CI(n38787), .I0(n1802[12]), .I1(GND_net), 
            .CO(n38788));
    SB_LUT4 add_3103_7_lut (.I0(GND_net), .I1(n8409[4]), .I2(n643), .I3(n38504), 
            .O(n8396[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_5_lut (.I0(GND_net), .I1(n12735[2]), .I2(n326), .I3(n38031), 
            .O(n12160[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_12_lut (.I0(GND_net), .I1(n9128[9]), .I2(GND_net), 
            .I3(n37552), .O(n7763[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_5 (.CI(n38031), .I0(n12735[2]), .I1(n326), .CO(n38032));
    SB_LUT4 add_3225_20_lut (.I0(GND_net), .I1(n11995[17]), .I2(GND_net), 
            .I3(n37412), .O(n11361[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_7 (.CI(n38504), .I0(n8409[4]), .I1(n643), .CO(n38505));
    SB_LUT4 add_3259_4_lut (.I0(GND_net), .I1(n12735[1]), .I2(n253), .I3(n38030), 
            .O(n12160[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_12 (.CI(n37552), .I0(n9128[9]), .I1(GND_net), .CO(n37553));
    SB_CARRY add_3259_4 (.CI(n38030), .I0(n12735[1]), .I1(n253), .CO(n38031));
    SB_CARRY add_3225_20 (.CI(n37412), .I0(n11995[17]), .I1(GND_net), 
            .CO(n37413));
    SB_LUT4 mult_14_add_1216_14_lut (.I0(GND_net), .I1(n1802[11]), .I2(GND_net), 
            .I3(n38786), .O(n1801[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_6_lut (.I0(GND_net), .I1(n8409[3]), .I2(n546), .I3(n38503), 
            .O(n8396[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3259_3_lut (.I0(GND_net), .I1(n12735[0]), .I2(n180), .I3(n38029), 
            .O(n12160[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_3 (.CI(n38029), .I0(n12735[0]), .I1(n180), .CO(n38030));
    SB_CARRY add_3103_6 (.CI(n38503), .I0(n8409[3]), .I1(n546), .CO(n38504));
    SB_LUT4 add_3259_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n12160[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3259_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3259_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n38029));
    SB_CARRY mult_14_add_1216_14 (.CI(n38786), .I0(n1802[11]), .I1(GND_net), 
            .CO(n38787));
    SB_LUT4 add_3103_5_lut (.I0(GND_net), .I1(n8409[2]), .I2(n449), .I3(n38502), 
            .O(n8396[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_11_lut (.I0(GND_net), .I1(n9128[8]), .I2(GND_net), 
            .I3(n37551), .O(n7763[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_19_lut (.I0(GND_net), .I1(n11995[16]), .I2(GND_net), 
            .I3(n37411), .O(n11361[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_5 (.CI(n38502), .I0(n8409[2]), .I1(n449), .CO(n38503));
    SB_CARRY add_3077_11 (.CI(n37551), .I0(n9128[8]), .I1(GND_net), .CO(n37552));
    SB_CARRY add_3225_19 (.CI(n37411), .I0(n11995[16]), .I1(GND_net), 
            .CO(n37412));
    SB_LUT4 mult_10_i333_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n495_adj_3511));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1216_13_lut (.I0(GND_net), .I1(n1802[10]), .I2(GND_net), 
            .I3(n38785), .O(n1801[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_4_lut (.I0(GND_net), .I1(n8409[1]), .I2(n352), .I3(n38501), 
            .O(n8396[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_4 (.CI(n38501), .I0(n8409[1]), .I1(n352), .CO(n38502));
    SB_CARRY mult_14_add_1216_13 (.CI(n38785), .I0(n1802[10]), .I1(GND_net), 
            .CO(n38786));
    SB_LUT4 add_3103_3_lut (.I0(GND_net), .I1(n8409[0]), .I2(n255), .I3(n38500), 
            .O(n8396[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_10_lut (.I0(GND_net), .I1(n9128[7]), .I2(GND_net), 
            .I3(n37550), .O(n7763[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_18_lut (.I0(GND_net), .I1(n11995[15]), .I2(GND_net), 
            .I3(n37410), .O(n11361[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_3 (.CI(n38500), .I0(n8409[0]), .I1(n255), .CO(n38501));
    SB_CARRY add_3077_10 (.CI(n37550), .I0(n9128[7]), .I1(GND_net), .CO(n37551));
    SB_CARRY add_3225_18 (.CI(n37410), .I0(n11995[15]), .I1(GND_net), 
            .CO(n37411));
    SB_LUT4 mult_14_add_1216_12_lut (.I0(GND_net), .I1(n1802[9]), .I2(GND_net), 
            .I3(n38784), .O(n1801[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3103_2_lut (.I0(GND_net), .I1(n65), .I2(n158), .I3(GND_net), 
            .O(n8396[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3103_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3103_2 (.CI(GND_net), .I0(n65), .I1(n158), .CO(n38500));
    SB_CARRY mult_14_add_1216_12 (.CI(n38784), .I0(n1802[9]), .I1(GND_net), 
            .CO(n38785));
    SB_LUT4 add_3102_13_lut (.I0(GND_net), .I1(n8396[10]), .I2(GND_net), 
            .I3(n38499), .O(n8382[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_9_lut (.I0(GND_net), .I1(n9128[6]), .I2(GND_net), 
            .I3(n37549), .O(n7763[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_17_lut (.I0(GND_net), .I1(n11995[14]), .I2(GND_net), 
            .I3(n37409), .O(n11361[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_12_lut (.I0(GND_net), .I1(n8396[9]), .I2(GND_net), 
            .I3(n38498), .O(n8382[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_12 (.CI(n38498), .I0(n8396[9]), .I1(GND_net), .CO(n38499));
    SB_CARRY add_22984_18 (.CI(n37201), .I0(n66[16]), .I1(n191[16]), .CO(n37202));
    SB_CARRY add_3077_9 (.CI(n37549), .I0(n9128[6]), .I1(GND_net), .CO(n37550));
    SB_CARRY add_3225_17 (.CI(n37409), .I0(n11995[14]), .I1(GND_net), 
            .CO(n37410));
    SB_LUT4 mult_14_add_1216_11_lut (.I0(GND_net), .I1(n1802[8]), .I2(GND_net), 
            .I3(n38783), .O(n1801[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_11_lut (.I0(GND_net), .I1(n8396[8]), .I2(GND_net), 
            .I3(n38497), .O(n8382[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_11 (.CI(n38497), .I0(n8396[8]), .I1(GND_net), .CO(n38498));
    SB_LUT4 mult_12_i160_2_lut (.I0(\Kd[2] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n237_adj_3512));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i160_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1216_11 (.CI(n38783), .I0(n1802[8]), .I1(GND_net), 
            .CO(n38784));
    SB_LUT4 add_3102_10_lut (.I0(GND_net), .I1(n8396[7]), .I2(GND_net), 
            .I3(n38496), .O(n8382[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i225_2_lut (.I0(\Kd[3] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n334));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1216_10_lut (.I0(GND_net), .I1(n1802[7]), .I2(GND_net), 
            .I3(n38782), .O(n1801[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_10 (.CI(n38782), .I0(n1802[7]), .I1(GND_net), 
            .CO(n38783));
    SB_LUT4 add_22984_17_lut (.I0(GND_net), .I1(n66[15]), .I2(n191[15]), 
            .I3(n37200), .O(\PID_CONTROLLER.result_31__N_2994 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_8_lut (.I0(GND_net), .I1(n9128[5]), .I2(n686_adj_3513), 
            .I3(n37548), .O(n7763[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_16_lut (.I0(GND_net), .I1(n11995[13]), .I2(GND_net), 
            .I3(n37408), .O(n11361[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_8 (.CI(n37548), .I0(n9128[5]), .I1(n686_adj_3513), 
            .CO(n37549));
    SB_LUT4 add_3077_7_lut (.I0(GND_net), .I1(n9128[4]), .I2(n589_adj_3514), 
            .I3(n37547), .O(n7763[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_9_lut (.I0(GND_net), .I1(n1802[6]), .I2(GND_net), 
            .I3(n38781), .O(n1801[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_17 (.CI(n37200), .I0(n66[15]), .I1(n191[15]), .CO(n37201));
    SB_CARRY add_3102_10 (.CI(n38496), .I0(n8396[7]), .I1(GND_net), .CO(n38497));
    SB_CARRY add_3077_7 (.CI(n37547), .I0(n9128[4]), .I1(n589_adj_3514), 
            .CO(n37548));
    SB_CARRY mult_14_add_1216_9 (.CI(n38781), .I0(n1802[6]), .I1(GND_net), 
            .CO(n38782));
    SB_LUT4 add_3077_6_lut (.I0(GND_net), .I1(n9128[3]), .I2(n492_adj_3515), 
            .I3(n37546), .O(n7763[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_9_lut (.I0(GND_net), .I1(n8396[6]), .I2(GND_net), 
            .I3(n38495), .O(n8382[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_6 (.CI(n37546), .I0(n9128[3]), .I1(n492_adj_3515), 
            .CO(n37547));
    SB_LUT4 add_3077_5_lut (.I0(GND_net), .I1(n9128[2]), .I2(n395_adj_3516), 
            .I3(n37545), .O(n7763[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_8_lut (.I0(GND_net), .I1(n1802[5]), .I2(n527), 
            .I3(n38780), .O(n1801[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_9 (.CI(n38495), .I0(n8396[6]), .I1(GND_net), .CO(n38496));
    SB_CARRY add_3077_5 (.CI(n37545), .I0(n9128[2]), .I1(n395_adj_3516), 
            .CO(n37546));
    SB_LUT4 add_3102_8_lut (.I0(GND_net), .I1(n8396[5]), .I2(n737_adj_3517), 
            .I3(n38494), .O(n8382[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_8 (.CI(n38494), .I0(n8396[5]), .I1(n737_adj_3517), 
            .CO(n38495));
    SB_LUT4 mult_12_i290_2_lut (.I0(\Kd[4] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n431));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3102_7_lut (.I0(GND_net), .I1(n8396[4]), .I2(n640_adj_3518), 
            .I3(n38493), .O(n8382[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_4_lut (.I0(GND_net), .I1(n9128[1]), .I2(n298_adj_3519), 
            .I3(n37544), .O(n7763[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_16 (.CI(n37408), .I0(n11995[13]), .I1(GND_net), 
            .CO(n37409));
    SB_LUT4 add_3225_15_lut (.I0(GND_net), .I1(n11995[12]), .I2(GND_net), 
            .I3(n37407), .O(n11361[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_7 (.CI(n38493), .I0(n8396[4]), .I1(n640_adj_3518), 
            .CO(n38494));
    SB_CARRY mult_14_add_1216_8 (.CI(n38780), .I0(n1802[5]), .I1(n527), 
            .CO(n38781));
    SB_LUT4 mult_14_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3102_6_lut (.I0(GND_net), .I1(n8396[3]), .I2(n543_adj_3520), 
            .I3(n38492), .O(n8382[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_6 (.CI(n38492), .I0(n8396[3]), .I1(n543_adj_3520), 
            .CO(n38493));
    SB_LUT4 mult_14_add_1216_7_lut (.I0(GND_net), .I1(n1802[4]), .I2(n454), 
            .I3(n38779), .O(n1801[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_5_lut (.I0(GND_net), .I1(n8396[2]), .I2(n446_adj_3522), 
            .I3(n38491), .O(n8382[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_5 (.CI(n38491), .I0(n8396[2]), .I1(n446_adj_3522), 
            .CO(n38492));
    SB_CARRY add_3077_4 (.CI(n37544), .I0(n9128[1]), .I1(n298_adj_3519), 
            .CO(n37545));
    SB_CARRY add_3225_15 (.CI(n37407), .I0(n11995[12]), .I1(GND_net), 
            .CO(n37408));
    SB_LUT4 add_3102_4_lut (.I0(GND_net), .I1(n8396[1]), .I2(n349_adj_3523), 
            .I3(n38490), .O(n8382[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_16_lut (.I0(GND_net), .I1(n66[14]), .I2(n191[14]), 
            .I3(n37199), .O(\PID_CONTROLLER.result_31__N_2994 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3077_3_lut (.I0(GND_net), .I1(n9128[0]), .I2(n201_adj_3524), 
            .I3(n37543), .O(n7763[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3077_3 (.CI(n37543), .I0(n9128[0]), .I1(n201_adj_3524), 
            .CO(n37544));
    SB_LUT4 add_3077_2_lut (.I0(GND_net), .I1(n11_adj_3525), .I2(n104_adj_3526), 
            .I3(GND_net), .O(n7763[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3077_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_4 (.CI(n38490), .I0(n8396[1]), .I1(n349_adj_3523), 
            .CO(n38491));
    SB_LUT4 add_3225_14_lut (.I0(GND_net), .I1(n11995[11]), .I2(GND_net), 
            .I3(n37406), .O(n11361[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_14 (.CI(n37406), .I0(n11995[11]), .I1(GND_net), 
            .CO(n37407));
    SB_CARRY add_3077_2 (.CI(GND_net), .I0(n11_adj_3525), .I1(n104_adj_3526), 
            .CO(n37543));
    SB_LUT4 add_3307_15_lut (.I0(GND_net), .I1(n13737[12]), .I2(GND_net), 
            .I3(n37542), .O(n13259[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_7 (.CI(n38779), .I0(n1802[4]), .I1(n454), 
            .CO(n38780));
    SB_CARRY add_22984_16 (.CI(n37199), .I0(n66[14]), .I1(n191[14]), .CO(n37200));
    SB_LUT4 add_3102_3_lut (.I0(GND_net), .I1(n8396[0]), .I2(n252_adj_3527), 
            .I3(n38489), .O(n8382[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n57[0]), 
            .CO(n37017));
    SB_CARRY add_3102_3 (.CI(n38489), .I0(n8396[0]), .I1(n252_adj_3527), 
            .CO(n38490));
    SB_LUT4 unary_minus_17_inv_0_i2_1_lut (.I0(\deadband[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[1]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3225_13_lut (.I0(GND_net), .I1(n11995[10]), .I2(GND_net), 
            .I3(n37405), .O(n11361[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3102_2_lut (.I0(GND_net), .I1(n62_adj_3529), .I2(n155_adj_3530), 
            .I3(GND_net), .O(n8382[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3102_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1216_6_lut (.I0(GND_net), .I1(n1802[3]), .I2(n381), 
            .I3(n38778), .O(n1801[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n64[31]), 
            .I3(n37016), .O(pwm_23__N_2951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_6 (.CI(n38778), .I0(n1802[3]), .I1(n381), 
            .CO(n38779));
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n592_adj_3531));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i355_2_lut (.I0(\Kd[5] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n528_adj_3532));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i420_2_lut (.I0(\Kd[6] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n625));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n689_adj_3533));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i485_2_lut (.I0(\Kd[7] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n722));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n58[0]));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n282[0]));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i3_1_lut (.I0(\deadband[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[2]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_17_inv_0_i4_1_lut (.I0(\deadband[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[3]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i2_2_lut (.I0(\Kd[0] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n191[0]));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1216_5_lut (.I0(GND_net), .I1(n1802[2]), .I2(n308), 
            .I3(n38777), .O(n1801[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i97_2_lut (.I0(\Kd[1] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n143_adj_3536));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i97_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1216_5 (.CI(n38777), .I0(n1802[2]), .I1(n308), 
            .CO(n38778));
    SB_LUT4 mult_14_add_1216_4_lut (.I0(GND_net), .I1(n1802[1]), .I2(n235_adj_3538), 
            .I3(n38776), .O(n1801[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i34_2_lut (.I0(\Kd[0] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_3539));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1216_4 (.CI(n38776), .I0(n1802[1]), .I1(n235_adj_3538), 
            .CO(n38777));
    SB_LUT4 mult_14_add_1216_3_lut (.I0(GND_net), .I1(n1802[0]), .I2(n162), 
            .I3(n38775), .O(n1801[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3102_2 (.CI(GND_net), .I0(n62_adj_3529), .I1(n155_adj_3530), 
            .CO(n38489));
    SB_LUT4 mult_12_i162_2_lut (.I0(\Kd[2] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n240_adj_3540));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i227_2_lut (.I0(\Kd[3] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n337));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i227_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1216_3 (.CI(n38775), .I0(n1802[0]), .I1(n162), 
            .CO(n38776));
    SB_LUT4 mult_14_add_1216_2_lut (.I0(GND_net), .I1(n20_adj_3541), .I2(n89), 
            .I3(GND_net), .O(n1801[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1216_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1216_2 (.CI(GND_net), .I0(n20_adj_3541), .I1(n89), 
            .CO(n38775));
    SB_LUT4 mult_14_add_1215_24_lut (.I0(GND_net), .I1(n1801[21]), .I2(GND_net), 
            .I3(n38773), .O(n1800[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i292_2_lut (.I0(\Kd[4] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n434));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i357_2_lut (.I0(\Kd[5] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n531_adj_3542));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i357_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1215_24 (.CI(n38773), .I0(n1801[21]), .I1(GND_net), 
            .CO(n1699));
    SB_LUT4 mult_14_add_1215_23_lut (.I0(GND_net), .I1(n1801[20]), .I2(GND_net), 
            .I3(n38772), .O(n1800[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_14_lut (.I0(GND_net), .I1(n8382[11]), .I2(GND_net), 
            .I3(n38488), .O(n8367[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_14_lut (.I0(GND_net), .I1(n13737[11]), .I2(GND_net), 
            .I3(n37541), .O(n13259[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_13_lut (.I0(GND_net), .I1(n8382[10]), .I2(GND_net), 
            .I3(n38487), .O(n8367[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_13 (.CI(n38487), .I0(n8382[10]), .I1(GND_net), .CO(n38488));
    SB_LUT4 add_22984_15_lut (.I0(GND_net), .I1(n66[13]), .I2(n191[13]), 
            .I3(n37198), .O(\PID_CONTROLLER.result_31__N_2994 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_14 (.CI(n37541), .I0(n13737[11]), .I1(GND_net), 
            .CO(n37542));
    SB_LUT4 add_3307_13_lut (.I0(GND_net), .I1(n13737[10]), .I2(GND_net), 
            .I3(n37540), .O(n13259[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_12_lut (.I0(GND_net), .I1(n8382[9]), .I2(GND_net), 
            .I3(n38486), .O(n8367[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_13 (.CI(n37540), .I0(n13737[10]), .I1(GND_net), 
            .CO(n37541));
    SB_LUT4 add_3307_12_lut (.I0(GND_net), .I1(n13737[9]), .I2(GND_net), 
            .I3(n37539), .O(n13259[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_13 (.CI(n37405), .I0(n11995[10]), .I1(GND_net), 
            .CO(n37406));
    SB_LUT4 mult_12_i422_2_lut (.I0(\Kd[6] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n628));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1215_23 (.CI(n38772), .I0(n1801[20]), .I1(GND_net), 
            .CO(n38773));
    SB_LUT4 mult_14_add_1215_22_lut (.I0(GND_net), .I1(n1801[19]), .I2(GND_net), 
            .I3(n38771), .O(n1800[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_12 (.CI(n38486), .I0(n8382[9]), .I1(GND_net), .CO(n38487));
    SB_CARRY add_3307_12 (.CI(n37539), .I0(n13737[9]), .I1(GND_net), .CO(n37540));
    SB_LUT4 mult_12_i487_2_lut (.I0(\Kd[7] ), .I1(n61[15]), .I2(GND_net), 
            .I3(GND_net), .O(n725));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3101_11_lut (.I0(GND_net), .I1(n8382[8]), .I2(GND_net), 
            .I3(n38485), .O(n8367[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF Kd_delay_counter_1046__i0 (.Q(Kd_delay_counter[0]), .C(clk32MHz), 
           .D(n69[0]));   // verilog/motorControl.v(48[27:47])
    SB_CARRY add_3101_11 (.CI(n38485), .I0(n8382[8]), .I1(GND_net), .CO(n38486));
    SB_LUT4 add_3101_10_lut (.I0(GND_net), .I1(n8382[7]), .I2(GND_net), 
            .I3(n38484), .O(n8367[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_11_lut (.I0(GND_net), .I1(n13737[8]), .I2(GND_net), 
            .I3(n37538), .O(n13259[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_10 (.CI(n38484), .I0(n8382[7]), .I1(GND_net), .CO(n38485));
    SB_LUT4 add_3101_9_lut (.I0(GND_net), .I1(n8382[6]), .I2(GND_net), 
            .I3(n38483), .O(n8367[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_9 (.CI(n38483), .I0(n8382[6]), .I1(GND_net), .CO(n38484));
    SB_LUT4 add_3101_8_lut (.I0(GND_net), .I1(n8382[5]), .I2(n734_adj_3543), 
            .I3(n38482), .O(n8367[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_22 (.CI(n38771), .I0(n1801[19]), .I1(GND_net), 
            .CO(n38772));
    SB_LUT4 mult_14_add_1215_21_lut (.I0(GND_net), .I1(n1801[18]), .I2(GND_net), 
            .I3(n38770), .O(n1800[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_12_lut (.I0(GND_net), .I1(n11995[9]), .I2(GND_net), 
            .I3(n37404), .O(n11361[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_21 (.CI(n38770), .I0(n1801[18]), .I1(GND_net), 
            .CO(n38771));
    SB_CARRY add_3101_8 (.CI(n38482), .I0(n8382[5]), .I1(n734_adj_3543), 
            .CO(n38483));
    SB_CARRY add_3225_12 (.CI(n37404), .I0(n11995[9]), .I1(GND_net), .CO(n37405));
    SB_LUT4 mult_14_add_1215_20_lut (.I0(GND_net), .I1(n1801[17]), .I2(GND_net), 
            .I3(n38769), .O(n1800[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_20 (.CI(n38769), .I0(n1801[17]), .I1(GND_net), 
            .CO(n38770));
    SB_LUT4 add_3101_7_lut (.I0(GND_net), .I1(n8382[4]), .I2(n637_adj_3544), 
            .I3(n38481), .O(n8367[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_15 (.CI(n37198), .I0(n66[13]), .I1(n191[13]), .CO(n37199));
    SB_CARRY add_3101_7 (.CI(n38481), .I0(n8382[4]), .I1(n637_adj_3544), 
            .CO(n38482));
    SB_LUT4 add_3101_6_lut (.I0(GND_net), .I1(n8382[3]), .I2(n540_adj_3545), 
            .I3(n38480), .O(n8367[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_11_lut (.I0(GND_net), .I1(n11995[8]), .I2(GND_net), 
            .I3(n37403), .O(n11361[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_14_lut (.I0(GND_net), .I1(n66[12]), .I2(n191[12]), 
            .I3(n37197), .O(\PID_CONTROLLER.result_31__N_2994 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n64[31]), 
            .I3(n37015), .O(pwm_23__N_2951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_6 (.CI(n38480), .I0(n8382[3]), .I1(n540_adj_3545), 
            .CO(n38481));
    SB_CARRY add_3225_11 (.CI(n37403), .I0(n11995[8]), .I1(GND_net), .CO(n37404));
    SB_LUT4 unary_minus_17_inv_0_i5_1_lut (.I0(\deadband[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[4]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3101_5_lut (.I0(GND_net), .I1(n8382[2]), .I2(n443_adj_3547), 
            .I3(n38479), .O(n8367[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_19_lut (.I0(GND_net), .I1(n1801[16]), .I2(GND_net), 
            .I3(n38768), .O(n1800[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_5 (.CI(n38479), .I0(n8382[2]), .I1(n443_adj_3547), 
            .CO(n38480));
    SB_CARRY add_3307_11 (.CI(n37538), .I0(n13737[8]), .I1(GND_net), .CO(n37539));
    SB_LUT4 add_3101_4_lut (.I0(GND_net), .I1(n8382[1]), .I2(n346_adj_3548), 
            .I3(n38478), .O(n8367[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_10_lut (.I0(GND_net), .I1(n11995[7]), .I2(GND_net), 
            .I3(n37402), .O(n11361[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_4 (.CI(n38478), .I0(n8382[1]), .I1(n346_adj_3548), 
            .CO(n38479));
    SB_LUT4 add_3307_10_lut (.I0(GND_net), .I1(n13737[7]), .I2(GND_net), 
            .I3(n37537), .O(n13259[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_10 (.CI(n37402), .I0(n11995[7]), .I1(GND_net), .CO(n37403));
    SB_CARRY mult_14_add_1215_19 (.CI(n38768), .I0(n1801[16]), .I1(GND_net), 
            .CO(n38769));
    SB_LUT4 add_3101_3_lut (.I0(GND_net), .I1(n8382[0]), .I2(n249_adj_3549), 
            .I3(n38477), .O(n8367[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_3 (.CI(n38477), .I0(n8382[0]), .I1(n249_adj_3549), 
            .CO(n38478));
    SB_LUT4 mult_14_add_1215_18_lut (.I0(GND_net), .I1(n1801[15]), .I2(GND_net), 
            .I3(n38767), .O(n1800[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3101_2_lut (.I0(GND_net), .I1(n59_adj_3550), .I2(n152_adj_3551), 
            .I3(GND_net), .O(n8367[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_10 (.CI(n37537), .I0(n13737[7]), .I1(GND_net), .CO(n37538));
    SB_LUT4 add_3307_9_lut (.I0(GND_net), .I1(n13737[6]), .I2(GND_net), 
            .I3(n37536), .O(n13259[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_9 (.CI(n37536), .I0(n13737[6]), .I1(GND_net), .CO(n37537));
    SB_LUT4 add_3225_9_lut (.I0(GND_net), .I1(n11995[6]), .I2(GND_net), 
            .I3(n37401), .O(n11361[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3101_2 (.CI(GND_net), .I0(n59_adj_3550), .I1(n152_adj_3551), 
            .CO(n38477));
    SB_CARRY mult_14_add_1215_18 (.CI(n38767), .I0(n1801[15]), .I1(GND_net), 
            .CO(n38768));
    SB_LUT4 add_3307_8_lut (.I0(GND_net), .I1(n13737[5]), .I2(n545), .I3(n37535), 
            .O(n13259[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_9 (.CI(n37401), .I0(n11995[6]), .I1(GND_net), .CO(n37402));
    SB_LUT4 mult_14_add_1215_17_lut (.I0(GND_net), .I1(n1801[14]), .I2(GND_net), 
            .I3(n38766), .O(n1800[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_15_lut (.I0(GND_net), .I1(n8367[12]), .I2(GND_net), 
            .I3(n38476), .O(n8351[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_14_lut (.I0(GND_net), .I1(n8367[11]), .I2(GND_net), 
            .I3(n38475), .O(n8351[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_17 (.CI(n38766), .I0(n1801[14]), .I1(GND_net), 
            .CO(n38767));
    SB_CARRY add_3100_14 (.CI(n38475), .I0(n8367[11]), .I1(GND_net), .CO(n38476));
    SB_CARRY add_3307_8 (.CI(n37535), .I0(n13737[5]), .I1(n545), .CO(n37536));
    SB_LUT4 add_3225_8_lut (.I0(GND_net), .I1(n11995[5]), .I2(n698), .I3(n37400), 
            .O(n11361[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_13_lut (.I0(GND_net), .I1(n8367[10]), .I2(GND_net), 
            .I3(n38474), .O(n8351[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_8 (.CI(n37400), .I0(n11995[5]), .I1(n698), .CO(n37401));
    SB_LUT4 add_3307_7_lut (.I0(GND_net), .I1(n13737[4]), .I2(n472), .I3(n37534), 
            .O(n13259[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_7_lut (.I0(GND_net), .I1(n11995[4]), .I2(n601_adj_3552), 
            .I3(n37399), .O(n11361[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3553));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1215_16_lut (.I0(GND_net), .I1(n1801[13]), .I2(GND_net), 
            .I3(n38765), .O(n1800[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_13 (.CI(n38474), .I0(n8367[10]), .I1(GND_net), .CO(n38475));
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n37982), .O(n70[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_12_lut (.I0(GND_net), .I1(n8367[9]), .I2(GND_net), 
            .I3(n38473), .O(n8351[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n37981), .O(n70[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_7 (.CI(n37534), .I0(n13737[4]), .I1(n472), .CO(n37535));
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_10  (.CI(n37981), .I0(\PID_CONTROLLER.err[8] ), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n37982));
    SB_CARRY mult_14_add_1215_16 (.CI(n38765), .I0(n1801[13]), .I1(GND_net), 
            .CO(n38766));
    SB_CARRY add_3100_12 (.CI(n38473), .I0(n8367[9]), .I1(GND_net), .CO(n38474));
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n37980), .O(n70[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_6_lut (.I0(GND_net), .I1(n13737[3]), .I2(n399), .I3(n37533), 
            .O(n13259[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_9  (.CI(n37980), .I0(\PID_CONTROLLER.err[7] ), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n37981));
    SB_LUT4 mult_14_add_1215_15_lut (.I0(GND_net), .I1(n1801[12]), .I2(GND_net), 
            .I3(n38764), .O(n1800[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_7 (.CI(n37399), .I0(n11995[4]), .I1(n601_adj_3552), 
            .CO(n37400));
    SB_LUT4 add_3100_11_lut (.I0(GND_net), .I1(n8367[8]), .I2(GND_net), 
            .I3(n38472), .O(n8351[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_6_lut (.I0(GND_net), .I1(n11995[3]), .I2(n504), .I3(n37398), 
            .O(n11361[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n37979), .O(n70[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_6 (.CI(n37533), .I0(n13737[3]), .I1(n399), .CO(n37534));
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_8  (.CI(n37979), .I0(\PID_CONTROLLER.err[6] ), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n37980));
    SB_CARRY add_3225_6 (.CI(n37398), .I0(n11995[3]), .I1(n504), .CO(n37399));
    SB_CARRY mult_14_add_1215_15 (.CI(n38764), .I0(n1801[12]), .I1(GND_net), 
            .CO(n38765));
    SB_CARRY add_3100_11 (.CI(n38472), .I0(n8367[8]), .I1(GND_net), .CO(n38473));
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n37978), .O(n70[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_7  (.CI(n37978), .I0(\PID_CONTROLLER.err[5] ), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n37979));
    SB_LUT4 add_3100_10_lut (.I0(GND_net), .I1(n8367[7]), .I2(GND_net), 
            .I3(n38471), .O(n8351[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n37977), .O(n70[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_6  (.CI(n37977), .I0(\PID_CONTROLLER.err[4] ), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n37978));
    SB_CARRY add_22984_14 (.CI(n37197), .I0(n66[12]), .I1(n191[12]), .CO(n37198));
    SB_LUT4 mult_14_add_1215_14_lut (.I0(GND_net), .I1(n1801[11]), .I2(GND_net), 
            .I3(n38763), .O(n1800[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3557));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n37976), .O(n70[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_10 (.CI(n38471), .I0(n8367[7]), .I1(GND_net), .CO(n38472));
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_5  (.CI(n37976), .I0(\PID_CONTROLLER.err[3] ), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n37977));
    SB_CARRY mult_14_add_1215_14 (.CI(n38763), .I0(n1801[11]), .I1(GND_net), 
            .CO(n38764));
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n37975), .O(n70[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3307_5_lut (.I0(GND_net), .I1(n13737[2]), .I2(n326), .I3(n37532), 
            .O(n13259[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_13_lut (.I0(GND_net), .I1(n66[11]), .I2(n191[11]), 
            .I3(n37196), .O(\PID_CONTROLLER.result_31__N_2994 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_4  (.CI(n37975), .I0(\PID_CONTROLLER.err[2] ), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n37976));
    SB_LUT4 add_3225_5_lut (.I0(GND_net), .I1(n11995[2]), .I2(n407), .I3(n37397), 
            .O(n11361[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_9_lut (.I0(GND_net), .I1(n8367[6]), .I2(GND_net), 
            .I3(n38470), .O(n8351[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n37974), .O(n70[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_11 (.CI(n37015), .I0(GND_net), .I1(n64[31]), 
            .CO(n37016));
    SB_CARRY add_3307_5 (.CI(n37532), .I0(n13737[2]), .I1(n326), .CO(n37533));
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_3  (.CI(n37974), .I0(\PID_CONTROLLER.err[1] ), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n37975));
    SB_CARRY add_3225_5 (.CI(n37397), .I0(n11995[2]), .I1(n407), .CO(n37398));
    SB_LUT4 mult_14_add_1215_13_lut (.I0(GND_net), .I1(n1801[10]), .I2(GND_net), 
            .I3(n38762), .O(n1800[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_9 (.CI(n38470), .I0(n8367[6]), .I1(GND_net), .CO(n38471));
    SB_LUT4 \PID_CONTROLLER.integral_1048_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n70[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1048_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_8_lut (.I0(GND_net), .I1(n8367[5]), .I2(n731_adj_3559), 
            .I3(n38469), .O(n8351[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1048_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err[0] ), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n37974));
    SB_LUT4 pwm_count_1047_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[8]), 
            .I3(n37973), .O(n73[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_8 (.CI(n38469), .I0(n8367[5]), .I1(n731_adj_3559), 
            .CO(n38470));
    SB_LUT4 add_3307_4_lut (.I0(GND_net), .I1(n13737[1]), .I2(n253), .I3(n37531), 
            .O(n13259[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1047_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[7]), 
            .I3(n37972), .O(n73[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_4_lut (.I0(GND_net), .I1(n11995[1]), .I2(n310), .I3(n37396), 
            .O(n11361[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1047_add_4_9 (.CI(n37972), .I0(GND_net), .I1(pwm_count[7]), 
            .CO(n37973));
    SB_CARRY add_22984_13 (.CI(n37196), .I0(n66[11]), .I1(n191[11]), .CO(n37197));
    SB_CARRY mult_14_add_1215_13 (.CI(n38762), .I0(n1801[10]), .I1(GND_net), 
            .CO(n38763));
    SB_LUT4 pwm_count_1047_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[6]), 
            .I3(n37971), .O(n73[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_12_lut (.I0(GND_net), .I1(n1801[9]), .I2(GND_net), 
            .I3(n38761), .O(n1800[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_7_lut (.I0(GND_net), .I1(n8367[4]), .I2(n634_adj_3561), 
            .I3(n38468), .O(n8351[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_7 (.CI(n38468), .I0(n8367[4]), .I1(n634_adj_3561), 
            .CO(n38469));
    SB_CARRY pwm_count_1047_add_4_8 (.CI(n37971), .I0(GND_net), .I1(pwm_count[6]), 
            .CO(n37972));
    SB_CARRY add_3307_4 (.CI(n37531), .I0(n13737[1]), .I1(n253), .CO(n37532));
    SB_LUT4 pwm_count_1047_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[5]), 
            .I3(n37970), .O(n73[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_12_lut (.I0(GND_net), .I1(n66[10]), .I2(n191[10]), 
            .I3(n37195), .O(\PID_CONTROLLER.result_31__N_2994 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_4 (.CI(n37396), .I0(n11995[1]), .I1(n310), .CO(n37397));
    SB_LUT4 add_3100_6_lut (.I0(GND_net), .I1(n8367[3]), .I2(n537_adj_3562), 
            .I3(n38467), .O(n8351[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1047_add_4_7 (.CI(n37970), .I0(GND_net), .I1(pwm_count[5]), 
            .CO(n37971));
    SB_LUT4 add_3307_3_lut (.I0(GND_net), .I1(n13737[0]), .I2(n180), .I3(n37530), 
            .O(n13259[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_12 (.CI(n37195), .I0(n66[10]), .I1(n191[10]), .CO(n37196));
    SB_LUT4 pwm_count_1047_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[4]), 
            .I3(n37969), .O(n73[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3225_3_lut (.I0(GND_net), .I1(n11995[0]), .I2(n213), .I3(n37395), 
            .O(n11361[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_12 (.CI(n38761), .I0(n1801[9]), .I1(GND_net), 
            .CO(n38762));
    SB_CARRY add_3100_6 (.CI(n38467), .I0(n8367[3]), .I1(n537_adj_3562), 
            .CO(n38468));
    SB_CARRY pwm_count_1047_add_4_6 (.CI(n37969), .I0(GND_net), .I1(pwm_count[4]), 
            .CO(n37970));
    SB_LUT4 add_22984_11_lut (.I0(GND_net), .I1(n66[9]), .I2(n191[9]), 
            .I3(n37194), .O(\PID_CONTROLLER.result_31__N_2994 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_5_lut (.I0(GND_net), .I1(n8367[2]), .I2(n440_adj_3564), 
            .I3(n38466), .O(n8351[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1047_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[3]), 
            .I3(n37968), .O(n73[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n64[8]), 
            .I3(n37014), .O(pwm_23__N_2951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_5 (.CI(n38466), .I0(n8367[2]), .I1(n440_adj_3564), 
            .CO(n38467));
    SB_CARRY pwm_count_1047_add_4_5 (.CI(n37968), .I0(GND_net), .I1(pwm_count[3]), 
            .CO(n37969));
    SB_LUT4 mult_14_add_1215_11_lut (.I0(GND_net), .I1(n1801[8]), .I2(GND_net), 
            .I3(n38760), .O(n1800[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1047_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[2]), 
            .I3(n37967), .O(n73[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3100_4_lut (.I0(GND_net), .I1(n8367[1]), .I2(n343_adj_3568), 
            .I3(n38465), .O(n8351[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_11 (.CI(n38760), .I0(n1801[8]), .I1(GND_net), 
            .CO(n38761));
    SB_LUT4 mult_12_i99_2_lut (.I0(\Kd[1] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n146_adj_3569));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i99_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY pwm_count_1047_add_4_4 (.CI(n37967), .I0(GND_net), .I1(pwm_count[2]), 
            .CO(n37968));
    SB_CARRY add_3100_4 (.CI(n38465), .I0(n8367[1]), .I1(n343_adj_3568), 
            .CO(n38466));
    SB_LUT4 pwm_count_1047_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[1]), 
            .I3(n37966), .O(n73[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_3 (.CI(n37530), .I0(n13737[0]), .I1(n180), .CO(n37531));
    SB_LUT4 add_3307_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n13259[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3307_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1047_add_4_3 (.CI(n37966), .I0(GND_net), .I1(pwm_count[1]), 
            .CO(n37967));
    SB_CARRY add_3225_3 (.CI(n37395), .I0(n11995[0]), .I1(n213), .CO(n37396));
    SB_LUT4 add_3100_3_lut (.I0(GND_net), .I1(n8367[0]), .I2(n246_adj_3571), 
            .I3(n38464), .O(n8351[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_count_1047_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_count[0]), 
            .I3(VCC_net), .O(n73[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_count_1047_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3307_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n37530));
    SB_LUT4 add_3131_29_lut (.I0(GND_net), .I1(n9932[26]), .I2(GND_net), 
            .I3(n37529), .O(n9128[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_count_1047_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_count[0]), 
            .CO(n37966));
    SB_LUT4 add_3225_2_lut (.I0(GND_net), .I1(n23_adj_3573), .I2(n116), 
            .I3(GND_net), .O(n11361[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_31_lut (.I0(GND_net), .I1(n7991[28]), .I2(GND_net), 
            .I3(n37965), .O(n7959[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_10_lut (.I0(GND_net), .I1(n1801[7]), .I2(GND_net), 
            .I3(n38759), .O(n1800[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_30_lut (.I0(GND_net), .I1(n7991[27]), .I2(GND_net), 
            .I3(n37964), .O(n7959[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3100_3 (.CI(n38464), .I0(n8367[0]), .I1(n246_adj_3571), 
            .CO(n38465));
    SB_CARRY unary_minus_17_add_3_10 (.CI(n37014), .I0(GND_net), .I1(n64[8]), 
            .CO(n37015));
    SB_CARRY add_3084_30 (.CI(n37964), .I0(n7991[27]), .I1(GND_net), .CO(n37965));
    SB_LUT4 add_3100_2_lut (.I0(GND_net), .I1(n56_adj_3574), .I2(n149_adj_3575), 
            .I3(GND_net), .O(n8351[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3100_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i36_2_lut (.I0(\Kd[0] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_3576));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3084_29_lut (.I0(GND_net), .I1(n7991[26]), .I2(GND_net), 
            .I3(n37963), .O(n7959[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_29 (.CI(n37963), .I0(n7991[26]), .I1(GND_net), .CO(n37964));
    SB_LUT4 add_3084_28_lut (.I0(GND_net), .I1(n7991[25]), .I2(GND_net), 
            .I3(n37962), .O(n7959[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_28 (.CI(n37962), .I0(n7991[25]), .I1(GND_net), .CO(n37963));
    SB_CARRY add_3100_2 (.CI(GND_net), .I0(n56_adj_3574), .I1(n149_adj_3575), 
            .CO(n38464));
    SB_LUT4 add_3084_27_lut (.I0(GND_net), .I1(n7991[24]), .I2(GND_net), 
            .I3(n37961), .O(n7959[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_16_lut (.I0(GND_net), .I1(n8351[13]), .I2(GND_net), 
            .I3(n38463), .O(n8334[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_27 (.CI(n37961), .I0(n7991[24]), .I1(GND_net), .CO(n37962));
    SB_CARRY mult_14_add_1215_10 (.CI(n38759), .I0(n1801[7]), .I1(GND_net), 
            .CO(n38760));
    SB_LUT4 add_3099_15_lut (.I0(GND_net), .I1(n8351[12]), .I2(GND_net), 
            .I3(n38462), .O(n8334[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_26_lut (.I0(GND_net), .I1(n7991[23]), .I2(GND_net), 
            .I3(n37960), .O(n7959[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_28_lut (.I0(GND_net), .I1(n9932[25]), .I2(GND_net), 
            .I3(n37528), .O(n9128[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_26 (.CI(n37960), .I0(n7991[23]), .I1(GND_net), .CO(n37961));
    SB_LUT4 add_3084_25_lut (.I0(GND_net), .I1(n7991[22]), .I2(GND_net), 
            .I3(n37959), .O(n7959[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3225_2 (.CI(GND_net), .I0(n23_adj_3573), .I1(n116), .CO(n37395));
    SB_CARRY add_3099_15 (.CI(n38462), .I0(n8351[12]), .I1(GND_net), .CO(n38463));
    SB_CARRY add_3084_25 (.CI(n37959), .I0(n7991[22]), .I1(GND_net), .CO(n37960));
    SB_CARRY add_3131_28 (.CI(n37528), .I0(n9932[25]), .I1(GND_net), .CO(n37529));
    SB_LUT4 add_3084_24_lut (.I0(GND_net), .I1(n7991[21]), .I2(GND_net), 
            .I3(n37958), .O(n7959[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_11_lut (.I0(GND_net), .I1(n15229[8]), .I2(GND_net), 
            .I3(n37394), .O(n14915[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_9_lut (.I0(GND_net), .I1(n1801[6]), .I2(GND_net), 
            .I3(n38758), .O(n1800[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n64[7]), 
            .I3(n37013), .O(\pwm_23__N_2951[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_10_lut (.I0(GND_net), .I1(n15229[7]), .I2(GND_net), 
            .I3(n37393), .O(n14915[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_14_lut (.I0(GND_net), .I1(n8351[11]), .I2(GND_net), 
            .I3(n38461), .O(n8334[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i69_2_lut (.I0(\Kd[1] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_3579));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i69_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1215_9 (.CI(n38758), .I0(n1801[6]), .I1(GND_net), 
            .CO(n38759));
    SB_CARRY add_3084_24 (.CI(n37958), .I0(n7991[21]), .I1(GND_net), .CO(n37959));
    SB_CARRY add_3099_14 (.CI(n38461), .I0(n8351[11]), .I1(GND_net), .CO(n38462));
    SB_LUT4 add_3084_23_lut (.I0(GND_net), .I1(n7991[20]), .I2(GND_net), 
            .I3(n37957), .O(n7959[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_23 (.CI(n37957), .I0(n7991[20]), .I1(GND_net), .CO(n37958));
    SB_LUT4 add_3084_22_lut (.I0(GND_net), .I1(n7991[19]), .I2(GND_net), 
            .I3(n37956), .O(n7959[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_13_lut (.I0(GND_net), .I1(n8351[10]), .I2(GND_net), 
            .I3(n38460), .O(n8334[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_13 (.CI(n38460), .I0(n8351[10]), .I1(GND_net), .CO(n38461));
    SB_LUT4 add_3131_27_lut (.I0(GND_net), .I1(n9932[24]), .I2(GND_net), 
            .I3(n37527), .O(n9128[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_22 (.CI(n37956), .I0(n7991[19]), .I1(GND_net), .CO(n37957));
    SB_CARRY add_3389_10 (.CI(n37393), .I0(n15229[7]), .I1(GND_net), .CO(n37394));
    SB_LUT4 add_3084_21_lut (.I0(GND_net), .I1(n7991[18]), .I2(GND_net), 
            .I3(n37955), .O(n7959[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_11 (.CI(n37194), .I0(n66[9]), .I1(n191[9]), .CO(n37195));
    SB_CARRY unary_minus_17_add_3_9 (.CI(n37013), .I0(GND_net), .I1(n64[7]), 
            .CO(n37014));
    SB_LUT4 mult_14_add_1215_8_lut (.I0(GND_net), .I1(n1801[5]), .I2(n524), 
            .I3(n38757), .O(n1800[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i6_2_lut (.I0(\Kd[0] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_3581));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i6_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1215_8 (.CI(n38757), .I0(n1801[5]), .I1(n524), 
            .CO(n38758));
    SB_LUT4 add_3099_12_lut (.I0(GND_net), .I1(n8351[9]), .I2(GND_net), 
            .I3(n38459), .O(n8334[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_21 (.CI(n37955), .I0(n7991[18]), .I1(GND_net), .CO(n37956));
    SB_CARRY add_3131_27 (.CI(n37527), .I0(n9932[24]), .I1(GND_net), .CO(n37528));
    SB_LUT4 add_3084_20_lut (.I0(GND_net), .I1(n7991[17]), .I2(GND_net), 
            .I3(n37954), .O(n7959[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_9_lut (.I0(GND_net), .I1(n15229[6]), .I2(GND_net), 
            .I3(n37392), .O(n14915[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_12 (.CI(n38459), .I0(n8351[9]), .I1(GND_net), .CO(n38460));
    SB_CARRY add_3084_20 (.CI(n37954), .I0(n7991[17]), .I1(GND_net), .CO(n37955));
    SB_LUT4 add_3131_26_lut (.I0(GND_net), .I1(n9932[23]), .I2(GND_net), 
            .I3(n37526), .O(n9128[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_19_lut (.I0(GND_net), .I1(n7991[16]), .I2(GND_net), 
            .I3(n37953), .O(n7959[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_9 (.CI(n37392), .I0(n15229[6]), .I1(GND_net), .CO(n37393));
    SB_LUT4 mult_14_add_1215_7_lut (.I0(GND_net), .I1(n1801[4]), .I2(n451), 
            .I3(n38756), .O(n1800[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_11_lut (.I0(GND_net), .I1(n8351[8]), .I2(GND_net), 
            .I3(n38458), .O(n8334[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_19 (.CI(n37953), .I0(n7991[16]), .I1(GND_net), .CO(n37954));
    SB_LUT4 add_3084_18_lut (.I0(GND_net), .I1(n7991[15]), .I2(GND_net), 
            .I3(n37952), .O(n7959[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_11 (.CI(n38458), .I0(n8351[8]), .I1(GND_net), .CO(n38459));
    SB_CARRY add_3084_18 (.CI(n37952), .I0(n7991[15]), .I1(GND_net), .CO(n37953));
    SB_LUT4 unary_minus_17_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n64[6]), 
            .I3(n37012), .O(\pwm_23__N_2951[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_10_lut (.I0(GND_net), .I1(n8351[7]), .I2(GND_net), 
            .I3(n38457), .O(n8334[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_17_lut (.I0(GND_net), .I1(n7991[14]), .I2(GND_net), 
            .I3(n37951), .O(n7959[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i134_2_lut (.I0(\Kd[2] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_3584));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1215_7 (.CI(n38756), .I0(n1801[4]), .I1(n451), 
            .CO(n38757));
    SB_CARRY add_3084_17 (.CI(n37951), .I0(n7991[14]), .I1(GND_net), .CO(n37952));
    SB_CARRY add_3099_10 (.CI(n38457), .I0(n8351[7]), .I1(GND_net), .CO(n38458));
    SB_CARRY add_3131_26 (.CI(n37526), .I0(n9932[23]), .I1(GND_net), .CO(n37527));
    SB_LUT4 add_3084_16_lut (.I0(GND_net), .I1(n7991[13]), .I2(GND_net), 
            .I3(n37950), .O(n7959[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_8_lut (.I0(GND_net), .I1(n15229[5]), .I2(n545), .I3(n37391), 
            .O(n14915[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_25_lut (.I0(GND_net), .I1(n9932[22]), .I2(GND_net), 
            .I3(n37525), .O(n9128[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_22984_10_lut (.I0(GND_net), .I1(n66[8]), .I2(n191[8]), 
            .I3(n37193), .O(\PID_CONTROLLER.result_31__N_2994 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_16 (.CI(n37950), .I0(n7991[13]), .I1(GND_net), .CO(n37951));
    SB_CARRY unary_minus_17_add_3_8 (.CI(n37012), .I0(GND_net), .I1(n64[6]), 
            .CO(n37013));
    SB_LUT4 unary_minus_17_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n64[5]), 
            .I3(n37011), .O(\pwm_23__N_2951[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_8 (.CI(n37391), .I0(n15229[5]), .I1(n545), .CO(n37392));
    SB_LUT4 add_3099_9_lut (.I0(GND_net), .I1(n8351[6]), .I2(GND_net), 
            .I3(n38456), .O(n8334[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_15_lut (.I0(GND_net), .I1(n7991[12]), .I2(GND_net), 
            .I3(n37949), .O(n7959[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_25 (.CI(n37525), .I0(n9932[22]), .I1(GND_net), .CO(n37526));
    SB_CARRY add_3084_15 (.CI(n37949), .I0(n7991[12]), .I1(GND_net), .CO(n37950));
    SB_LUT4 add_3389_7_lut (.I0(GND_net), .I1(n15229[4]), .I2(n472), .I3(n37390), 
            .O(n14915[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_6_lut (.I0(GND_net), .I1(n1801[3]), .I2(n378), 
            .I3(n38755), .O(n1800[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_9 (.CI(n38456), .I0(n8351[6]), .I1(GND_net), .CO(n38457));
    SB_LUT4 add_3084_14_lut (.I0(GND_net), .I1(n7991[11]), .I2(GND_net), 
            .I3(n37948), .O(n7959[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_14 (.CI(n37948), .I0(n7991[11]), .I1(GND_net), .CO(n37949));
    SB_LUT4 add_3099_8_lut (.I0(GND_net), .I1(n8351[5]), .I2(n728_adj_3586), 
            .I3(n38455), .O(n8334[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_13_lut (.I0(GND_net), .I1(n7991[10]), .I2(GND_net), 
            .I3(n37947), .O(n7959[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_13 (.CI(n37947), .I0(n7991[10]), .I1(GND_net), .CO(n37948));
    SB_CARRY mult_14_add_1215_6 (.CI(n38755), .I0(n1801[3]), .I1(n378), 
            .CO(n38756));
    SB_CARRY add_3099_8 (.CI(n38455), .I0(n8351[5]), .I1(n728_adj_3586), 
            .CO(n38456));
    SB_LUT4 add_3084_12_lut (.I0(GND_net), .I1(n7991[9]), .I2(GND_net), 
            .I3(n37946), .O(n7959[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_24_lut (.I0(GND_net), .I1(n9932[21]), .I2(GND_net), 
            .I3(n37524), .O(n9128[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_12 (.CI(n37946), .I0(n7991[9]), .I1(GND_net), .CO(n37947));
    SB_LUT4 mult_12_i199_2_lut (.I0(\Kd[3] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n295_adj_3587));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i199_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3389_7 (.CI(n37390), .I0(n15229[4]), .I1(n472), .CO(n37391));
    SB_LUT4 add_3099_7_lut (.I0(GND_net), .I1(n8351[4]), .I2(n631_adj_3588), 
            .I3(n38454), .O(n8334[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1215_5_lut (.I0(GND_net), .I1(n1801[2]), .I2(n305), 
            .I3(n38754), .O(n1800[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_11_lut (.I0(GND_net), .I1(n7991[8]), .I2(GND_net), 
            .I3(n37945), .O(n7959[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_7 (.CI(n38454), .I0(n8351[4]), .I1(n631_adj_3588), 
            .CO(n38455));
    SB_LUT4 mult_12_i164_2_lut (.I0(\Kd[2] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n243_adj_3589));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i164_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1215_5 (.CI(n38754), .I0(n1801[2]), .I1(n305), 
            .CO(n38755));
    SB_CARRY add_3084_11 (.CI(n37945), .I0(n7991[8]), .I1(GND_net), .CO(n37946));
    SB_CARRY add_3131_24 (.CI(n37524), .I0(n9932[21]), .I1(GND_net), .CO(n37525));
    SB_LUT4 add_3084_10_lut (.I0(GND_net), .I1(n7991[7]), .I2(GND_net), 
            .I3(n37944), .O(n7959[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_10 (.CI(n37944), .I0(n7991[7]), .I1(GND_net), .CO(n37945));
    SB_LUT4 mult_14_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3099_6_lut (.I0(GND_net), .I1(n8351[3]), .I2(n534_adj_3590), 
            .I3(n38453), .O(n8334[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_6_lut (.I0(GND_net), .I1(n15229[3]), .I2(n399), .I3(n37389), 
            .O(n14915[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_9_lut (.I0(GND_net), .I1(n7991[6]), .I2(GND_net), 
            .I3(n37943), .O(n7959[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i264_2_lut (.I0(\Kd[4] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n392_adj_3591));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i264_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3099_6 (.CI(n38453), .I0(n8351[3]), .I1(n534_adj_3590), 
            .CO(n38454));
    SB_CARRY add_3084_9 (.CI(n37943), .I0(n7991[6]), .I1(GND_net), .CO(n37944));
    SB_LUT4 add_3131_23_lut (.I0(GND_net), .I1(n9932[20]), .I2(GND_net), 
            .I3(n37523), .O(n9128[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_23 (.CI(n37523), .I0(n9932[20]), .I1(GND_net), .CO(n37524));
    SB_LUT4 add_3084_8_lut (.I0(GND_net), .I1(n7991[5]), .I2(n683_adj_3592), 
            .I3(n37942), .O(n7959[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_8 (.CI(n37942), .I0(n7991[5]), .I1(n683_adj_3592), 
            .CO(n37943));
    SB_LUT4 mult_12_i229_2_lut (.I0(\Kd[3] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n340_adj_3593));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1215_4_lut (.I0(GND_net), .I1(n1801[1]), .I2(n232_adj_3595), 
            .I3(n38753), .O(n1800[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3099_5_lut (.I0(GND_net), .I1(n8351[2]), .I2(n437_adj_3596), 
            .I3(n38452), .O(n8334[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_7_lut (.I0(GND_net), .I1(n7991[4]), .I2(n586_adj_3597), 
            .I3(n37941), .O(n7959[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_7 (.CI(n37941), .I0(n7991[4]), .I1(n586_adj_3597), 
            .CO(n37942));
    SB_CARRY add_3099_5 (.CI(n38452), .I0(n8351[2]), .I1(n437_adj_3596), 
            .CO(n38453));
    SB_LUT4 add_3084_6_lut (.I0(GND_net), .I1(n7991[3]), .I2(n489_adj_3598), 
            .I3(n37940), .O(n7959[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_6 (.CI(n37940), .I0(n7991[3]), .I1(n489_adj_3598), 
            .CO(n37941));
    SB_CARRY mult_14_add_1215_4 (.CI(n38753), .I0(n1801[1]), .I1(n232_adj_3595), 
            .CO(n38754));
    SB_LUT4 add_3099_4_lut (.I0(GND_net), .I1(n8351[1]), .I2(n340_adj_3593), 
            .I3(n38451), .O(n8334[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_5_lut (.I0(GND_net), .I1(n7991[2]), .I2(n392_adj_3591), 
            .I3(n37939), .O(n7959[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_22_lut (.I0(GND_net), .I1(n9932[19]), .I2(GND_net), 
            .I3(n37522), .O(n9128[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_5 (.CI(n37939), .I0(n7991[2]), .I1(n392_adj_3591), 
            .CO(n37940));
    SB_CARRY add_3389_6 (.CI(n37389), .I0(n15229[3]), .I1(n399), .CO(n37390));
    SB_LUT4 mult_14_add_1215_3_lut (.I0(GND_net), .I1(n1801[0]), .I2(n159), 
            .I3(n38752), .O(n1800[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_4 (.CI(n38451), .I0(n8351[1]), .I1(n340_adj_3593), 
            .CO(n38452));
    SB_LUT4 add_3099_3_lut (.I0(GND_net), .I1(n8351[0]), .I2(n243_adj_3589), 
            .I3(n38450), .O(n8334[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_4_lut (.I0(GND_net), .I1(n7991[1]), .I2(n295_adj_3587), 
            .I3(n37938), .O(n7959[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_4 (.CI(n37938), .I0(n7991[1]), .I1(n295_adj_3587), 
            .CO(n37939));
    SB_CARRY add_3131_22 (.CI(n37522), .I0(n9932[19]), .I1(GND_net), .CO(n37523));
    SB_LUT4 add_3131_21_lut (.I0(GND_net), .I1(n9932[18]), .I2(GND_net), 
            .I3(n37521), .O(n9128[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3084_3_lut (.I0(GND_net), .I1(n7991[0]), .I2(n198_adj_3584), 
            .I3(n37937), .O(n7959[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3084_3 (.CI(n37937), .I0(n7991[0]), .I1(n198_adj_3584), 
            .CO(n37938));
    SB_LUT4 add_3389_5_lut (.I0(GND_net), .I1(n15229[2]), .I2(n326), .I3(n37388), 
            .O(n14915[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_5 (.CI(n37388), .I0(n15229[2]), .I1(n326), .CO(n37389));
    SB_CARRY add_22984_10 (.CI(n37193), .I0(n66[8]), .I1(n191[8]), .CO(n37194));
    SB_LUT4 mult_12_i329_2_lut (.I0(\Kd[5] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n489_adj_3598));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i329_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1215_3 (.CI(n38752), .I0(n1801[0]), .I1(n159), 
            .CO(n38753));
    SB_LUT4 add_3084_2_lut (.I0(GND_net), .I1(n8_adj_3581), .I2(n101_adj_3579), 
            .I3(GND_net), .O(n7959[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3084_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_3 (.CI(n38450), .I0(n8351[0]), .I1(n243_adj_3589), 
            .CO(n38451));
    SB_LUT4 add_3099_2_lut (.I0(GND_net), .I1(n53_adj_3576), .I2(n146_adj_3569), 
            .I3(GND_net), .O(n8334[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3099_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_7 (.CI(n37011), .I0(GND_net), .I1(n64[5]), 
            .CO(n37012));
    SB_LUT4 add_3389_4_lut (.I0(GND_net), .I1(n15229[1]), .I2(n253), .I3(n37387), 
            .O(n14915[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3099_2 (.CI(GND_net), .I0(n53_adj_3576), .I1(n146_adj_3569), 
            .CO(n38450));
    SB_CARRY add_3084_2 (.CI(GND_net), .I0(n8_adj_3581), .I1(n101_adj_3579), 
            .CO(n37937));
    SB_LUT4 add_22984_9_lut (.I0(GND_net), .I1(n66[7]), .I2(n191[7]), 
            .I3(n37192), .O(\PID_CONTROLLER.result_31__N_2994 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_16_lut (.I0(GND_net), .I1(n13259[13]), .I2(GND_net), 
            .I3(n37936), .O(n12735[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_15_lut (.I0(GND_net), .I1(n13259[12]), .I2(GND_net), 
            .I3(n37935), .O(n12735[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_21 (.CI(n37521), .I0(n9932[18]), .I1(GND_net), .CO(n37522));
    SB_LUT4 add_3131_20_lut (.I0(GND_net), .I1(n9932[17]), .I2(GND_net), 
            .I3(n37520), .O(n9128[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_15 (.CI(n37935), .I0(n13259[12]), .I1(GND_net), 
            .CO(n37936));
    SB_LUT4 mult_14_add_1215_2_lut (.I0(GND_net), .I1(n17_adj_3557), .I2(n86_adj_3553), 
            .I3(GND_net), .O(n1800[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1215_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_14_lut (.I0(GND_net), .I1(n13259[11]), .I2(GND_net), 
            .I3(n37934), .O(n12735[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_17_lut (.I0(GND_net), .I1(n8334[14]), .I2(GND_net), 
            .I3(n38449), .O(n8316[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_14 (.CI(n37934), .I0(n13259[11]), .I1(GND_net), 
            .CO(n37935));
    SB_LUT4 add_3284_13_lut (.I0(GND_net), .I1(n13259[10]), .I2(GND_net), 
            .I3(n37933), .O(n12735[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1215_2 (.CI(GND_net), .I0(n17_adj_3557), .I1(n86_adj_3553), 
            .CO(n38752));
    SB_LUT4 add_3098_16_lut (.I0(GND_net), .I1(n8334[13]), .I2(GND_net), 
            .I3(n38448), .O(n8316[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_13 (.CI(n37933), .I0(n13259[10]), .I1(GND_net), 
            .CO(n37934));
    SB_CARRY add_3131_20 (.CI(n37520), .I0(n9932[17]), .I1(GND_net), .CO(n37521));
    SB_LUT4 add_3284_12_lut (.I0(GND_net), .I1(n13259[9]), .I2(GND_net), 
            .I3(n37932), .O(n12735[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_4 (.CI(n37387), .I0(n15229[1]), .I1(n253), .CO(n37388));
    SB_CARRY add_3098_16 (.CI(n38448), .I0(n8334[13]), .I1(GND_net), .CO(n38449));
    SB_CARRY add_3284_12 (.CI(n37932), .I0(n13259[9]), .I1(GND_net), .CO(n37933));
    SB_LUT4 add_3131_19_lut (.I0(GND_net), .I1(n9932[16]), .I2(GND_net), 
            .I3(n37519), .O(n9128[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_11_lut (.I0(GND_net), .I1(n13259[8]), .I2(GND_net), 
            .I3(n37931), .O(n12735[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_15_lut (.I0(GND_net), .I1(n8334[12]), .I2(GND_net), 
            .I3(n38447), .O(n8316[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n64[4]), 
            .I3(n37010), .O(pwm_23__N_2951[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_3_lut (.I0(GND_net), .I1(n15229[0]), .I2(n180), .I3(n37386), 
            .O(n14915[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_15 (.CI(n38447), .I0(n8334[12]), .I1(GND_net), .CO(n38448));
    SB_CARRY add_22984_9 (.CI(n37192), .I0(n66[7]), .I1(n191[7]), .CO(n37193));
    SB_CARRY add_3284_11 (.CI(n37931), .I0(n13259[8]), .I1(GND_net), .CO(n37932));
    SB_LUT4 mult_14_add_1214_24_lut (.I0(GND_net), .I1(n1800[21]), .I2(GND_net), 
            .I3(n38750), .O(n1799[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_3 (.CI(n37386), .I0(n15229[0]), .I1(n180), .CO(n37387));
    SB_CARRY add_3131_19 (.CI(n37519), .I0(n9932[16]), .I1(GND_net), .CO(n37520));
    SB_LUT4 add_3098_14_lut (.I0(GND_net), .I1(n8334[11]), .I2(GND_net), 
            .I3(n38446), .O(n8316[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_18_lut (.I0(GND_net), .I1(n9932[15]), .I2(GND_net), 
            .I3(n37518), .O(n9128[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_10_lut (.I0(GND_net), .I1(n13259[7]), .I2(GND_net), 
            .I3(n37930), .O(n12735[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_10 (.CI(n37930), .I0(n13259[7]), .I1(GND_net), .CO(n37931));
    SB_LUT4 add_22984_8_lut (.I0(GND_net), .I1(n66[6]), .I2(n191[6]), 
            .I3(n37191), .O(\PID_CONTROLLER.result_31__N_2994 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3389_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n14915[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3389_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3389_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n37386));
    SB_CARRY mult_14_add_1214_24 (.CI(n38750), .I0(n1800[21]), .I1(GND_net), 
            .CO(n1695));
    SB_CARRY add_3098_14 (.CI(n38446), .I0(n8334[11]), .I1(GND_net), .CO(n38447));
    SB_LUT4 mult_12_i394_2_lut (.I0(\Kd[6] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n586_adj_3597));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3098_13_lut (.I0(GND_net), .I1(n8334[10]), .I2(GND_net), 
            .I3(n38445), .O(n8316[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_9_lut (.I0(GND_net), .I1(n13259[6]), .I2(GND_net), 
            .I3(n37929), .O(n12735[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_13 (.CI(n38445), .I0(n8334[10]), .I1(GND_net), .CO(n38446));
    SB_CARRY add_3284_9 (.CI(n37929), .I0(n13259[6]), .I1(GND_net), .CO(n37930));
    SB_LUT4 add_3098_12_lut (.I0(GND_net), .I1(n8334[9]), .I2(GND_net), 
            .I3(n38444), .O(n8316[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_18 (.CI(n37518), .I0(n9932[15]), .I1(GND_net), .CO(n37519));
    SB_LUT4 add_3284_8_lut (.I0(GND_net), .I1(n13259[5]), .I2(n545), .I3(n37928), 
            .O(n12735[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_17_lut (.I0(GND_net), .I1(n9932[14]), .I2(GND_net), 
            .I3(n37517), .O(n9128[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_8 (.CI(n37928), .I0(n13259[5]), .I1(n545), .CO(n37929));
    SB_LUT4 add_3284_7_lut (.I0(GND_net), .I1(n13259[4]), .I2(n472), .I3(n37927), 
            .O(n12735[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_23_lut (.I0(GND_net), .I1(n1800[20]), .I2(GND_net), 
            .I3(n38749), .O(n1799[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_12 (.CI(n38444), .I0(n8334[9]), .I1(GND_net), .CO(n38445));
    SB_CARRY add_3284_7 (.CI(n37927), .I0(n13259[4]), .I1(n472), .CO(n37928));
    SB_CARRY add_3131_17 (.CI(n37517), .I0(n9932[14]), .I1(GND_net), .CO(n37518));
    SB_LUT4 add_3284_6_lut (.I0(GND_net), .I1(n13259[3]), .I2(n399), .I3(n37926), 
            .O(n12735[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_11_lut (.I0(GND_net), .I1(n8334[8]), .I2(GND_net), 
            .I3(n38443), .O(n8316[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_6 (.CI(n37926), .I0(n13259[3]), .I1(n399), .CO(n37927));
    SB_LUT4 add_3131_16_lut (.I0(GND_net), .I1(n9932[13]), .I2(GND_net), 
            .I3(n37516), .O(n9128[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_5_lut (.I0(GND_net), .I1(n13259[2]), .I2(n326), .I3(n37925), 
            .O(n12735[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_23 (.CI(n38749), .I0(n1800[20]), .I1(GND_net), 
            .CO(n38750));
    SB_CARRY add_3098_11 (.CI(n38443), .I0(n8334[8]), .I1(GND_net), .CO(n38444));
    SB_CARRY add_3284_5 (.CI(n37925), .I0(n13259[2]), .I1(n326), .CO(n37926));
    SB_LUT4 add_3284_4_lut (.I0(GND_net), .I1(n13259[1]), .I2(n253), .I3(n37924), 
            .O(n12735[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_4 (.CI(n37924), .I0(n13259[1]), .I1(n253), .CO(n37925));
    SB_LUT4 add_3098_10_lut (.I0(GND_net), .I1(n8334[7]), .I2(GND_net), 
            .I3(n38442), .O(n8316[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i294_2_lut (.I0(\Kd[4] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n437_adj_3596));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3284_3_lut (.I0(GND_net), .I1(n13259[0]), .I2(n180), .I3(n37923), 
            .O(n12735[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_3 (.CI(n37923), .I0(n13259[0]), .I1(n180), .CO(n37924));
    SB_LUT4 mult_14_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_3595));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_22_lut (.I0(GND_net), .I1(n1800[19]), .I2(GND_net), 
            .I3(n38748), .O(n1799[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_22 (.CI(n38748), .I0(n1800[19]), .I1(GND_net), 
            .CO(n38749));
    SB_CARRY add_3098_10 (.CI(n38442), .I0(n8334[7]), .I1(GND_net), .CO(n38443));
    SB_LUT4 mult_14_add_1214_21_lut (.I0(GND_net), .I1(n1800[18]), .I2(GND_net), 
            .I3(n38747), .O(n1799[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_9_lut (.I0(GND_net), .I1(n8334[6]), .I2(GND_net), 
            .I3(n38441), .O(n8316[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3284_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n12735[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3284_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3284_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n37923));
    SB_CARRY add_3131_16 (.CI(n37516), .I0(n9932[13]), .I1(GND_net), .CO(n37517));
    SB_LUT4 add_13_add_1_22984_add_1_33_lut (.I0(GND_net), .I1(n7068[8]), 
            .I2(n5789[0]), .I3(n37922), .O(n66[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_9 (.CI(n38441), .I0(n8334[6]), .I1(GND_net), .CO(n38442));
    SB_LUT4 add_13_add_1_22984_add_1_32_lut (.I0(GND_net), .I1(n7068[7]), 
            .I2(n58[30]), .I3(n37921), .O(n66[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_15_lut (.I0(GND_net), .I1(n9932[12]), .I2(GND_net), 
            .I3(n37515), .O(n9128[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_32 (.CI(n37921), .I0(n7068[7]), .I1(n58[30]), 
            .CO(n37922));
    SB_CARRY mult_14_add_1214_21 (.CI(n38747), .I0(n1800[18]), .I1(GND_net), 
            .CO(n38748));
    SB_LUT4 add_3098_8_lut (.I0(GND_net), .I1(n8334[5]), .I2(n725), .I3(n38440), 
            .O(n8316[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i440_2_lut (.I0(\Kd[6] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n655));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i440_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_22984_add_1_31_lut (.I0(GND_net), .I1(n7068[6]), 
            .I2(n58[29]), .I3(n37920), .O(n66[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_31 (.CI(n37920), .I0(n7068[6]), .I1(n58[29]), 
            .CO(n37921));
    SB_LUT4 mult_12_i459_2_lut (.I0(\Kd[7] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n683_adj_3592));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3098_8 (.CI(n38440), .I0(n8334[5]), .I1(n725), .CO(n38441));
    SB_LUT4 add_3098_7_lut (.I0(GND_net), .I1(n8334[4]), .I2(n628), .I3(n38439), 
            .O(n8316[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_30_lut (.I0(GND_net), .I1(n7068[5]), 
            .I2(n58[28]), .I3(n37919), .O(n66[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_30 (.CI(n37919), .I0(n7068[5]), .I1(n58[28]), 
            .CO(n37920));
    SB_LUT4 add_13_add_1_22984_add_1_29_lut (.I0(GND_net), .I1(n7068[4]), 
            .I2(n58[27]), .I3(n37918), .O(n66[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i505_2_lut (.I0(\Kd[7] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_3420));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_20_lut (.I0(GND_net), .I1(n1800[17]), .I2(GND_net), 
            .I3(n38746), .O(n1799[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i95_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3418));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i95_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3098_7 (.CI(n38439), .I0(n8334[4]), .I1(n628), .CO(n38440));
    SB_CARRY add_13_add_1_22984_add_1_29 (.CI(n37918), .I0(n7068[4]), .I1(n58[27]), 
            .CO(n37919));
    SB_CARRY mult_14_add_1214_20 (.CI(n38746), .I0(n1800[17]), .I1(GND_net), 
            .CO(n38747));
    SB_CARRY add_3131_15 (.CI(n37515), .I0(n9932[12]), .I1(GND_net), .CO(n37516));
    SB_LUT4 add_13_add_1_22984_add_1_28_lut (.I0(GND_net), .I1(n7068[3]), 
            .I2(n58[26]), .I3(n37917), .O(n66[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_6_lut (.I0(GND_net), .I1(n8334[3]), .I2(n531_adj_3542), 
            .I3(n38438), .O(n8316[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_28 (.CI(n37917), .I0(n7068[3]), .I1(n58[26]), 
            .CO(n37918));
    SB_LUT4 add_3131_14_lut (.I0(GND_net), .I1(n9932[11]), .I2(GND_net), 
            .I3(n37514), .O(n9128[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_27_lut (.I0(GND_net), .I1(n7068[2]), 
            .I2(n58[25]), .I3(n37916), .O(n66[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_19_lut (.I0(GND_net), .I1(n1800[16]), .I2(GND_net), 
            .I3(n38745), .O(n1799[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_6 (.CI(n38438), .I0(n8334[3]), .I1(n531_adj_3542), 
            .CO(n38439));
    SB_CARRY add_13_add_1_22984_add_1_27 (.CI(n37916), .I0(n7068[2]), .I1(n58[25]), 
            .CO(n37917));
    SB_LUT4 add_13_add_1_22984_add_1_26_lut (.I0(GND_net), .I1(n7068[1]), 
            .I2(n58[24]), .I3(n37915), .O(n66[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_5_lut (.I0(GND_net), .I1(n8334[2]), .I2(n434), .I3(n38437), 
            .O(n8316[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_8 (.CI(n37191), .I0(n66[6]), .I1(n191[6]), .CO(n37192));
    SB_CARRY add_13_add_1_22984_add_1_26 (.CI(n37915), .I0(n7068[1]), .I1(n58[24]), 
            .CO(n37916));
    SB_CARRY mult_14_add_1214_19 (.CI(n38745), .I0(n1800[16]), .I1(GND_net), 
            .CO(n38746));
    SB_LUT4 add_13_add_1_22984_add_1_25_lut (.I0(GND_net), .I1(n7068[0]), 
            .I2(n58[23]), .I3(n37914), .O(n66[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_5 (.CI(n38437), .I0(n8334[2]), .I1(n434), .CO(n38438));
    SB_LUT4 mult_14_add_1214_18_lut (.I0(GND_net), .I1(n1800[15]), .I2(GND_net), 
            .I3(n38744), .O(n1799[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_4_lut (.I0(GND_net), .I1(n8334[1]), .I2(n337), .I3(n38436), 
            .O(n8316[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i144_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i144_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3098_4 (.CI(n38436), .I0(n8334[1]), .I1(n337), .CO(n38437));
    SB_LUT4 mult_14_i193_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i193_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_13_add_1_22984_add_1_25 (.CI(n37914), .I0(n7068[0]), .I1(n58[23]), 
            .CO(n37915));
    SB_LUT4 mult_14_i242_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i242_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i291_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i291_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_22984_add_1_24_lut (.I0(GND_net), .I1(n282[22]), 
            .I2(n58[22]), .I3(n37913), .O(n66[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_14 (.CI(n37514), .I0(n9932[11]), .I1(GND_net), .CO(n37515));
    SB_CARRY add_13_add_1_22984_add_1_24 (.CI(n37913), .I0(n282[22]), .I1(n58[22]), 
            .CO(n37914));
    SB_LUT4 add_22984_7_lut (.I0(GND_net), .I1(n66[5]), .I2(n191[5]), 
            .I3(n37190), .O(\PID_CONTROLLER.result_31__N_2994 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_25_lut (.I0(GND_net), .I1(n12578[22]), .I2(GND_net), 
            .I3(n37379), .O(n11995[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3098_3_lut (.I0(GND_net), .I1(n8334[0]), .I2(n240_adj_3540), 
            .I3(n38435), .O(n8316[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_7 (.CI(n37190), .I0(n66[5]), .I1(n191[5]), .CO(n37191));
    SB_LUT4 add_13_add_1_22984_add_1_23_lut (.I0(GND_net), .I1(n282[21]), 
            .I2(n58[21]), .I3(n37912), .O(n66[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_13_lut (.I0(GND_net), .I1(n9932[10]), .I2(GND_net), 
            .I3(n37513), .O(n9128[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_23 (.CI(n37912), .I0(n282[21]), .I1(n58[21]), 
            .CO(n37913));
    SB_LUT4 add_3251_24_lut (.I0(GND_net), .I1(n12578[21]), .I2(GND_net), 
            .I3(n37378), .O(n11995[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_18 (.CI(n38744), .I0(n1800[15]), .I1(GND_net), 
            .CO(n38745));
    SB_CARRY add_3098_3 (.CI(n38435), .I0(n8334[0]), .I1(n240_adj_3540), 
            .CO(n38436));
    SB_LUT4 add_13_add_1_22984_add_1_22_lut (.I0(GND_net), .I1(n282[20]), 
            .I2(n58[20]), .I3(n37911), .O(n66[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_22 (.CI(n37911), .I0(n282[20]), .I1(n58[20]), 
            .CO(n37912));
    SB_LUT4 add_3098_2_lut (.I0(GND_net), .I1(n50_adj_3539), .I2(n143_adj_3536), 
            .I3(GND_net), .O(n8316[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3098_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_21_lut (.I0(GND_net), .I1(n282[19]), 
            .I2(n58[19]), .I3(n37910), .O(n66[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_21 (.CI(n37910), .I0(n282[19]), .I1(n58[19]), 
            .CO(n37911));
    SB_LUT4 mult_14_add_1214_17_lut (.I0(GND_net), .I1(n1800[14]), .I2(GND_net), 
            .I3(n38743), .O(n1799[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3098_2 (.CI(GND_net), .I0(n50_adj_3539), .I1(n143_adj_3536), 
            .CO(n38435));
    SB_LUT4 add_13_add_1_22984_add_1_20_lut (.I0(GND_net), .I1(n282[18]), 
            .I2(n58[18]), .I3(n37909), .O(n66[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_13 (.CI(n37513), .I0(n9932[10]), .I1(GND_net), .CO(n37514));
    SB_LUT4 add_22984_6_lut (.I0(GND_net), .I1(n66[4]), .I2(n191[4]), 
            .I3(n37189), .O(\PID_CONTROLLER.result_31__N_2994 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_20 (.CI(n37909), .I0(n282[18]), .I1(n58[18]), 
            .CO(n37910));
    SB_CARRY add_3251_24 (.CI(n37378), .I0(n12578[21]), .I1(GND_net), 
            .CO(n37379));
    SB_CARRY mult_14_add_1214_17 (.CI(n38743), .I0(n1800[14]), .I1(GND_net), 
            .CO(n38744));
    SB_LUT4 mult_14_i340_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i340_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i389_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i389_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3097_18_lut (.I0(GND_net), .I1(n8316[15]), .I2(GND_net), 
            .I3(n38434), .O(n8297[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_19_lut (.I0(GND_net), .I1(n282[17]), 
            .I2(n58[17]), .I3(n37908), .O(n66[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_12_lut (.I0(GND_net), .I1(n9932[9]), .I2(GND_net), 
            .I3(n37512), .O(n9128[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_19 (.CI(n37908), .I0(n282[17]), .I1(n58[17]), 
            .CO(n37909));
    SB_LUT4 add_3251_23_lut (.I0(GND_net), .I1(n12578[20]), .I2(GND_net), 
            .I3(n37377), .O(n11995[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_16_lut (.I0(GND_net), .I1(n1800[13]), .I2(GND_net), 
            .I3(n38742), .O(n1799[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_17_lut (.I0(GND_net), .I1(n8316[14]), .I2(GND_net), 
            .I3(n38433), .O(n8297[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_18_lut (.I0(GND_net), .I1(n282[16]), 
            .I2(n58[16]), .I3(n37907), .O(n66[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_18 (.CI(n37907), .I0(n282[16]), .I1(n58[16]), 
            .CO(n37908));
    SB_CARRY add_3097_17 (.CI(n38433), .I0(n8316[14]), .I1(GND_net), .CO(n38434));
    SB_LUT4 add_13_add_1_22984_add_1_17_lut (.I0(GND_net), .I1(n282[15]), 
            .I2(n58[15]), .I3(n37906), .O(n66[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_17 (.CI(n37906), .I0(n282[15]), .I1(n58[15]), 
            .CO(n37907));
    SB_CARRY mult_14_add_1214_16 (.CI(n38742), .I0(n1800[13]), .I1(GND_net), 
            .CO(n38743));
    SB_LUT4 add_3097_16_lut (.I0(GND_net), .I1(n8316[13]), .I2(GND_net), 
            .I3(n38432), .O(n8297[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_16_lut (.I0(GND_net), .I1(n282[14]), 
            .I2(n58[14]), .I3(n37905), .O(n66[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_23 (.CI(n37377), .I0(n12578[20]), .I1(GND_net), 
            .CO(n37378));
    SB_CARRY add_13_add_1_22984_add_1_16 (.CI(n37905), .I0(n282[14]), .I1(n58[14]), 
            .CO(n37906));
    SB_LUT4 add_13_add_1_22984_add_1_15_lut (.I0(GND_net), .I1(n282[13]), 
            .I2(n58[13]), .I3(n37904), .O(n66[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_12 (.CI(n37512), .I0(n9932[9]), .I1(GND_net), .CO(n37513));
    SB_LUT4 mult_12_i67_2_lut (.I0(\Kd[1] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_3415));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_13_add_1_22984_add_1_15 (.CI(n37904), .I0(n282[13]), .I1(n58[13]), 
            .CO(n37905));
    SB_LUT4 mult_12_i359_2_lut (.I0(\Kd[5] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n534_adj_3590));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3251_22_lut (.I0(GND_net), .I1(n12578[19]), .I2(GND_net), 
            .I3(n37376), .O(n11995[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i4_2_lut (.I0(\Kd[0] ), .I1(n61[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_3414));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_15_lut (.I0(GND_net), .I1(n1800[12]), .I2(GND_net), 
            .I3(n38741), .O(n1799[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_16 (.CI(n38432), .I0(n8316[13]), .I1(GND_net), .CO(n38433));
    SB_LUT4 add_13_add_1_22984_add_1_14_lut (.I0(GND_net), .I1(n282[12]), 
            .I2(n58[12]), .I3(n37903), .O(n66[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_11_lut (.I0(GND_net), .I1(n9932[8]), .I2(GND_net), 
            .I3(n37511), .O(n9128[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_14 (.CI(n37903), .I0(n282[12]), .I1(n58[12]), 
            .CO(n37904));
    SB_CARRY add_3251_22 (.CI(n37376), .I0(n12578[19]), .I1(GND_net), 
            .CO(n37377));
    SB_CARRY mult_14_add_1214_15 (.CI(n38741), .I0(n1800[12]), .I1(GND_net), 
            .CO(n38742));
    SB_LUT4 add_3097_15_lut (.I0(GND_net), .I1(n8316[12]), .I2(GND_net), 
            .I3(n38431), .O(n8297[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_15 (.CI(n38431), .I0(n8316[12]), .I1(GND_net), .CO(n38432));
    SB_LUT4 mult_12_i132_2_lut (.I0(\Kd[2] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_3412));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3097_14_lut (.I0(GND_net), .I1(n8316[11]), .I2(GND_net), 
            .I3(n38430), .O(n8297[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i197_2_lut (.I0(\Kd[3] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n292_adj_3410));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3408));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_22984_add_1_13_lut (.I0(GND_net), .I1(n282[11]), 
            .I2(n58[11]), .I3(n37902), .O(n66[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_13 (.CI(n37902), .I0(n282[11]), .I1(n58[11]), 
            .CO(n37903));
    SB_CARRY add_3097_14 (.CI(n38430), .I0(n8316[11]), .I1(GND_net), .CO(n38431));
    SB_LUT4 add_13_add_1_22984_add_1_12_lut (.I0(GND_net), .I1(n282[10]), 
            .I2(n58[10]), .I3(n37901), .O(n66[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_12 (.CI(n37901), .I0(n282[10]), .I1(n58[10]), 
            .CO(n37902));
    SB_LUT4 mult_14_add_1214_14_lut (.I0(GND_net), .I1(n1800[11]), .I2(GND_net), 
            .I3(n38740), .O(n1799[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_13_lut (.I0(GND_net), .I1(n8316[10]), .I2(GND_net), 
            .I3(n38429), .O(n8297[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_11_lut (.I0(GND_net), .I1(n282[9]), 
            .I2(n58[9]), .I3(n37900), .O(n66[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_11 (.CI(n37511), .I0(n9932[8]), .I1(GND_net), .CO(n37512));
    SB_LUT4 add_3251_21_lut (.I0(GND_net), .I1(n12578[18]), .I2(GND_net), 
            .I3(n37375), .O(n11995[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_6 (.CI(n37189), .I0(n66[4]), .I1(n191[4]), .CO(n37190));
    SB_CARRY add_13_add_1_22984_add_1_11 (.CI(n37900), .I0(n282[9]), .I1(n58[9]), 
            .CO(n37901));
    SB_LUT4 add_13_add_1_22984_add_1_10_lut (.I0(GND_net), .I1(n282[8]), 
            .I2(n58[8]), .I3(n37899), .O(n66[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_21 (.CI(n37375), .I0(n12578[18]), .I1(GND_net), 
            .CO(n37376));
    SB_LUT4 add_22984_5_lut (.I0(GND_net), .I1(n66[3]), .I2(n191[3]), 
            .I3(n37188), .O(\PID_CONTROLLER.result_31__N_2994 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_22984_5 (.CI(n37188), .I0(n66[3]), .I1(n191[3]), .CO(n37189));
    SB_CARRY add_3097_13 (.CI(n38429), .I0(n8316[10]), .I1(GND_net), .CO(n38430));
    SB_CARRY add_13_add_1_22984_add_1_10 (.CI(n37899), .I0(n282[8]), .I1(n58[8]), 
            .CO(n37900));
    SB_LUT4 add_3251_20_lut (.I0(GND_net), .I1(n12578[17]), .I2(GND_net), 
            .I3(n37374), .O(n11995[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3131_10_lut (.I0(GND_net), .I1(n9932[7]), .I2(GND_net), 
            .I3(n37510), .O(n9128[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_9_lut (.I0(GND_net), .I1(n282[7]), 
            .I2(n58[7]), .I3(n37898), .O(n66[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i262_2_lut (.I0(\Kd[4] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n389_adj_3407));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i327_2_lut (.I0(\Kd[5] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n486_adj_3404));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_22984_4_lut (.I0(GND_net), .I1(n66[2]), .I2(n191[2]), 
            .I3(n37187), .O(\PID_CONTROLLER.result_31__N_2994 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_20 (.CI(n37374), .I0(n12578[17]), .I1(GND_net), 
            .CO(n37375));
    SB_CARRY add_22984_4 (.CI(n37187), .I0(n66[2]), .I1(n191[2]), .CO(n37188));
    SB_CARRY add_13_add_1_22984_add_1_9 (.CI(n37898), .I0(n282[7]), .I1(n58[7]), 
            .CO(n37899));
    SB_LUT4 add_22984_3_lut (.I0(GND_net), .I1(n66[1]), .I2(n191[1]), 
            .I3(n37186), .O(\PID_CONTROLLER.result_31__N_2994 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_14 (.CI(n38740), .I0(n1800[11]), .I1(GND_net), 
            .CO(n38741));
    SB_LUT4 add_3097_12_lut (.I0(GND_net), .I1(n8316[9]), .I2(GND_net), 
            .I3(n38428), .O(n8297[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_8_lut (.I0(GND_net), .I1(n282[6]), 
            .I2(n58[6]), .I3(n37897), .O(n66[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_8 (.CI(n37897), .I0(n282[6]), .I1(n58[6]), 
            .CO(n37898));
    SB_CARRY add_3097_12 (.CI(n38428), .I0(n8316[9]), .I1(GND_net), .CO(n38429));
    SB_LUT4 mult_14_add_1214_13_lut (.I0(GND_net), .I1(n1800[10]), .I2(GND_net), 
            .I3(n38739), .O(n1799[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_13 (.CI(n38739), .I0(n1800[10]), .I1(GND_net), 
            .CO(n38740));
    SB_LUT4 add_13_add_1_22984_add_1_7_lut (.I0(GND_net), .I1(n282[5]), 
            .I2(n58[5]), .I3(n37896), .O(n66[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_7 (.CI(n37896), .I0(n282[5]), .I1(n58[5]), 
            .CO(n37897));
    SB_LUT4 add_3251_19_lut (.I0(GND_net), .I1(n12578[16]), .I2(GND_net), 
            .I3(n37373), .O(n11995[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_12_lut (.I0(GND_net), .I1(n1800[9]), .I2(GND_net), 
            .I3(n38738), .O(n1799[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_12 (.CI(n38738), .I0(n1800[9]), .I1(GND_net), 
            .CO(n38739));
    SB_CARRY add_22984_3 (.CI(n37186), .I0(n66[1]), .I1(n191[1]), .CO(n37187));
    SB_LUT4 add_3097_11_lut (.I0(GND_net), .I1(n8316[8]), .I2(GND_net), 
            .I3(n38427), .O(n8297[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_6 (.CI(n37010), .I0(GND_net), .I1(n64[4]), 
            .CO(n37011));
    SB_LUT4 mult_10_i197_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n292));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i197_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_13_add_1_22984_add_1_6_lut (.I0(GND_net), .I1(n282[4]), 
            .I2(n58[4]), .I3(n37895), .O(n66[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i392_2_lut (.I0(\Kd[6] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n583_adj_3402));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i392_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3131_10 (.CI(n37510), .I0(n9932[7]), .I1(GND_net), .CO(n37511));
    SB_CARRY add_3251_19 (.CI(n37373), .I0(n12578[16]), .I1(GND_net), 
            .CO(n37374));
    SB_LUT4 add_22984_2_lut (.I0(GND_net), .I1(n66[0]), .I2(n191[0]), 
            .I3(GND_net), .O(\PID_CONTROLLER.result_31__N_2994 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_22984_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n64[3]), 
            .I3(n37009), .O(pwm_23__N_2951[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_6 (.CI(n37895), .I0(n282[4]), .I1(n58[4]), 
            .CO(n37896));
    SB_CARRY add_22984_2 (.CI(GND_net), .I0(n66[0]), .I1(n191[0]), .CO(n37186));
    SB_CARRY unary_minus_17_add_3_5 (.CI(n37009), .I0(GND_net), .I1(n64[3]), 
            .CO(n37010));
    SB_LUT4 mult_14_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i206_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3097_11 (.CI(n38427), .I0(n8316[8]), .I1(GND_net), .CO(n38428));
    SB_LUT4 add_13_add_1_22984_add_1_5_lut (.I0(GND_net), .I1(n282[3]), 
            .I2(n58[3]), .I3(n37894), .O(n66[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_9_lut (.I0(GND_net), .I1(n9932[6]), .I2(GND_net), 
            .I3(n37509), .O(n9128[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_18_lut (.I0(GND_net), .I1(n12578[15]), .I2(GND_net), 
            .I3(n37372), .O(n11995[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i424_2_lut (.I0(\Kd[6] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n631_adj_3588));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i489_2_lut (.I0(\Kd[7] ), .I1(n61[16]), .I2(GND_net), 
            .I3(GND_net), .O(n728_adj_3586));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_17_inv_0_i6_1_lut (.I0(\deadband[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[5]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i262_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n389));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i262_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_11_lut (.I0(GND_net), .I1(n1800[8]), .I2(GND_net), 
            .I3(n38737), .O(n1799[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_19_lut (.I0(GND_net), .I1(n15117[16]), .I2(GND_net), 
            .I3(n37185), .O(n14796[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_5 (.CI(n37894), .I0(n282[3]), .I1(n58[3]), 
            .CO(n37895));
    SB_LUT4 add_3382_18_lut (.I0(GND_net), .I1(n15117[15]), .I2(GND_net), 
            .I3(n37184), .O(n14796[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n64[2]), 
            .I3(n37008), .O(pwm_23__N_2951[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_11 (.CI(n38737), .I0(n1800[8]), .I1(GND_net), 
            .CO(n38738));
    SB_LUT4 mult_14_add_1214_10_lut (.I0(GND_net), .I1(n1800[7]), .I2(GND_net), 
            .I3(n38736), .O(n1799[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_10_lut (.I0(GND_net), .I1(n8316[7]), .I2(GND_net), 
            .I3(n38426), .O(n8297[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i7_1_lut (.I0(\deadband[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[6]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_13_add_1_22984_add_1_4_lut (.I0(GND_net), .I1(n282[2]), 
            .I2(n58[2]), .I3(n37893), .O(n66[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i457_2_lut (.I0(\Kd[7] ), .I1(n61[0]), .I2(GND_net), 
            .I3(GND_net), .O(n680_adj_3400));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i327_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n486));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i327_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i392_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n583));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n680_adj_3398));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_13_add_1_22984_add_1_4 (.CI(n37893), .I0(n282[2]), .I1(n58[2]), 
            .CO(n37894));
    SB_CARRY add_3097_10 (.CI(n38426), .I0(n8316[7]), .I1(GND_net), .CO(n38427));
    SB_CARRY add_3251_18 (.CI(n37372), .I0(n12578[15]), .I1(GND_net), 
            .CO(n37373));
    SB_LUT4 add_13_add_1_22984_add_1_3_lut (.I0(GND_net), .I1(n282[1]), 
            .I2(n58[1]), .I3(n37892), .O(n66[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_3 (.CI(n37892), .I0(n282[1]), .I1(n58[1]), 
            .CO(n37893));
    SB_CARRY mult_14_add_1214_10 (.CI(n38736), .I0(n1800[7]), .I1(GND_net), 
            .CO(n38737));
    SB_LUT4 add_3097_9_lut (.I0(GND_net), .I1(n8316[6]), .I2(GND_net), 
            .I3(n38425), .O(n8297[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_add_1_22984_add_1_2_lut (.I0(GND_net), .I1(n282[0]), 
            .I2(n58[0]), .I3(GND_net), .O(n66[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_add_1_22984_add_1_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_18 (.CI(n37184), .I0(n15117[15]), .I1(GND_net), 
            .CO(n37185));
    SB_CARRY add_3097_9 (.CI(n38425), .I0(n8316[6]), .I1(GND_net), .CO(n38426));
    SB_LUT4 add_3382_17_lut (.I0(GND_net), .I1(n15117[14]), .I2(GND_net), 
            .I3(n37183), .O(n14796[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_17 (.CI(n37183), .I0(n15117[14]), .I1(GND_net), 
            .CO(n37184));
    SB_CARRY add_3131_9 (.CI(n37509), .I0(n9932[6]), .I1(GND_net), .CO(n37510));
    SB_LUT4 add_3251_17_lut (.I0(GND_net), .I1(n12578[14]), .I2(GND_net), 
            .I3(n37371), .O(n11995[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_add_1_22984_add_1_2 (.CI(GND_net), .I0(n282[0]), .I1(n58[0]), 
            .CO(n37892));
    SB_LUT4 Kd_delay_counter_1046_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[6]), .I3(n37891), .O(n69[6])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1046_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_16_lut (.I0(GND_net), .I1(n15117[13]), .I2(GND_net), 
            .I3(n37182), .O(n14796[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_8_lut (.I0(GND_net), .I1(n8316[5]), .I2(n722), .I3(n38424), 
            .O(n8297[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1046_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[5]), .I3(n37890), .O(n69[5])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1046_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_8_lut (.I0(GND_net), .I1(n9932[5]), .I2(n689_adj_3533), 
            .I3(n37508), .O(n9128[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_17 (.CI(n37371), .I0(n12578[14]), .I1(GND_net), 
            .CO(n37372));
    SB_CARRY Kd_delay_counter_1046_add_4_7 (.CI(n37890), .I0(GND_net), .I1(Kd_delay_counter[5]), 
            .CO(n37891));
    SB_CARRY add_3382_16 (.CI(n37182), .I0(n15117[13]), .I1(GND_net), 
            .CO(n37183));
    SB_LUT4 mult_14_add_1214_9_lut (.I0(GND_net), .I1(n1800[6]), .I2(GND_net), 
            .I3(n38735), .O(n1799[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_8 (.CI(n38424), .I0(n8316[5]), .I1(n722), .CO(n38425));
    SB_LUT4 Kd_delay_counter_1046_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[4]), .I3(n37889), .O(n69[4])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1046_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1046_add_4_6 (.CI(n37889), .I0(GND_net), .I1(Kd_delay_counter[4]), 
            .CO(n37890));
    SB_LUT4 add_3097_7_lut (.I0(GND_net), .I1(n8316[4]), .I2(n625), .I3(n38423), 
            .O(n8297[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1046_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[3]), .I3(n37888), .O(n69[3])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1046_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1046_add_4_5 (.CI(n37888), .I0(GND_net), .I1(Kd_delay_counter[3]), 
            .CO(n37889));
    SB_CARRY mult_14_add_1214_9 (.CI(n38735), .I0(n1800[6]), .I1(GND_net), 
            .CO(n38736));
    SB_CARRY add_3097_7 (.CI(n38423), .I0(n8316[4]), .I1(n625), .CO(n38424));
    SB_LUT4 Kd_delay_counter_1046_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[2]), .I3(n37887), .O(n69[2])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1046_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_8 (.CI(n37508), .I0(n9932[5]), .I1(n689_adj_3533), 
            .CO(n37509));
    SB_LUT4 add_3251_16_lut (.I0(GND_net), .I1(n12578[13]), .I2(GND_net), 
            .I3(n37370), .O(n11995[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_15_lut (.I0(GND_net), .I1(n15117[12]), .I2(GND_net), 
            .I3(n37181), .O(n14796[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY Kd_delay_counter_1046_add_4_4 (.CI(n37887), .I0(GND_net), .I1(Kd_delay_counter[2]), 
            .CO(n37888));
    SB_CARRY add_3382_15 (.CI(n37181), .I0(n15117[12]), .I1(GND_net), 
            .CO(n37182));
    SB_CARRY unary_minus_17_add_3_4 (.CI(n37008), .I0(GND_net), .I1(n64[2]), 
            .CO(n37009));
    SB_LUT4 add_3097_6_lut (.I0(GND_net), .I1(n8316[3]), .I2(n528_adj_3532), 
            .I3(n38422), .O(n8297[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_14_lut (.I0(GND_net), .I1(n15117[11]), .I2(GND_net), 
            .I3(n37180), .O(n14796[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1046_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[1]), .I3(n37886), .O(n69[1])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1046_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_7_lut (.I0(GND_net), .I1(n9932[4]), .I2(n592_adj_3531), 
            .I3(n37507), .O(n9128[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_16 (.CI(n37370), .I0(n12578[13]), .I1(GND_net), 
            .CO(n37371));
    SB_CARRY add_3382_14 (.CI(n37180), .I0(n15117[11]), .I1(GND_net), 
            .CO(n37181));
    SB_CARRY Kd_delay_counter_1046_add_4_3 (.CI(n37886), .I0(GND_net), .I1(Kd_delay_counter[1]), 
            .CO(n37887));
    SB_LUT4 add_3382_13_lut (.I0(GND_net), .I1(n15117[10]), .I2(GND_net), 
            .I3(n37179), .O(n14796[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1047__i0 (.Q(pwm_count[0]), .C(clk32MHz), .D(n73[0]));   // verilog/motorControl.v(99[18:29])
    SB_CARRY add_3382_13 (.CI(n37179), .I0(n15117[10]), .I1(GND_net), 
            .CO(n37180));
    SB_LUT4 unary_minus_17_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n64[1]), 
            .I3(n37007), .O(pwm_23__N_2951[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_15_lut (.I0(GND_net), .I1(n12578[12]), .I2(GND_net), 
            .I3(n37369), .O(n11995[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_15 (.CI(n37369), .I0(n12578[12]), .I1(GND_net), 
            .CO(n37370));
    SB_CARRY add_3097_6 (.CI(n38422), .I0(n8316[3]), .I1(n528_adj_3532), 
            .CO(n38423));
    SB_LUT4 add_3251_14_lut (.I0(GND_net), .I1(n12578[11]), .I2(GND_net), 
            .I3(n37368), .O(n11995[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1214_8_lut (.I0(GND_net), .I1(n1800[5]), .I2(n521), 
            .I3(n38734), .O(n1799[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 Kd_delay_counter_1046_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(Kd_delay_counter[0]), .I3(VCC_net), .O(n69[0])) /* synthesis syn_instantiated=1 */ ;
    defparam Kd_delay_counter_1046_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3097_5_lut (.I0(GND_net), .I1(n8316[2]), .I2(n431), .I3(n38421), 
            .O(n8297[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_14 (.CI(n37368), .I0(n12578[11]), .I1(GND_net), 
            .CO(n37369));
    SB_CARRY Kd_delay_counter_1046_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(Kd_delay_counter[0]), .CO(n37886));
    SB_LUT4 add_3251_13_lut (.I0(GND_net), .I1(n12578[10]), .I2(GND_net), 
            .I3(n37367), .O(n11995[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_13 (.CI(n37367), .I0(n12578[10]), .I1(GND_net), 
            .CO(n37368));
    SB_CARRY add_3097_5 (.CI(n38421), .I0(n8316[2]), .I1(n431), .CO(n38422));
    SB_LUT4 add_3097_4_lut (.I0(GND_net), .I1(n8316[1]), .I2(n334), .I3(n38420), 
            .O(n8297[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_12_lut (.I0(GND_net), .I1(n15117[9]), .I2(GND_net), 
            .I3(n37178), .O(n14796[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_12 (.CI(n37178), .I0(n15117[9]), .I1(GND_net), .CO(n37179));
    SB_LUT4 add_3382_11_lut (.I0(GND_net), .I1(n15117[8]), .I2(GND_net), 
            .I3(n37177), .O(n14796[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_8 (.CI(n38734), .I0(n1800[5]), .I1(n521), 
            .CO(n38735));
    SB_CARRY add_3097_4 (.CI(n38420), .I0(n8316[1]), .I1(n334), .CO(n38421));
    SB_LUT4 unary_minus_17_inv_0_i8_1_lut (.I0(\deadband[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[7]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3382_11 (.CI(n37177), .I0(n15117[8]), .I1(GND_net), .CO(n37178));
    SB_LUT4 add_3097_3_lut (.I0(GND_net), .I1(n8316[0]), .I2(n237_adj_3512), 
            .I3(n38419), .O(n8297[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_12_lut (.I0(GND_net), .I1(n12578[9]), .I2(GND_net), 
            .I3(n37366), .O(n11995[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i101_2_lut (.I0(\Kd[1] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n149_adj_3575));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i101_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3131_7 (.CI(n37507), .I0(n9932[4]), .I1(n592_adj_3531), 
            .CO(n37508));
    SB_LUT4 add_3131_6_lut (.I0(GND_net), .I1(n9932[3]), .I2(n495_adj_3511), 
            .I3(n37506), .O(n9128[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_12 (.CI(n37366), .I0(n12578[9]), .I1(GND_net), .CO(n37367));
    SB_LUT4 add_3382_10_lut (.I0(GND_net), .I1(n15117[7]), .I2(GND_net), 
            .I3(n37176), .O(n14796[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_10 (.CI(n37176), .I0(n15117[7]), .I1(GND_net), .CO(n37177));
    SB_LUT4 add_3382_9_lut (.I0(GND_net), .I1(n15117[6]), .I2(GND_net), 
            .I3(n37175), .O(n14796[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_11_lut (.I0(GND_net), .I1(n12578[8]), .I2(GND_net), 
            .I3(n37365), .O(n11995[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i38_2_lut (.I0(\Kd[0] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_3574));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3393));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_7_lut (.I0(GND_net), .I1(n1800[4]), .I2(n448), 
            .I3(n38733), .O(n1799[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3097_3 (.CI(n38419), .I0(n8316[0]), .I1(n237_adj_3512), 
            .CO(n38420));
    SB_CARRY add_3251_11 (.CI(n37365), .I0(n12578[8]), .I1(GND_net), .CO(n37366));
    SB_LUT4 mult_14_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i163_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_9 (.CI(n37175), .I0(n15117[6]), .I1(GND_net), .CO(n37176));
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[7] ), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3573));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i166_2_lut (.I0(\Kd[2] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n246_adj_3571));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i231_2_lut (.I0(\Kd[3] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n343_adj_3568));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i71_2_lut (.I0(\Kd[1] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3097_2_lut (.I0(GND_net), .I1(n47), .I2(n140_adj_3508), 
            .I3(GND_net), .O(n8297[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3097_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_10_lut (.I0(GND_net), .I1(n12578[7]), .I2(GND_net), 
            .I3(n37364), .O(n11995[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3382_8_lut (.I0(GND_net), .I1(n15117[5]), .I2(n719), .I3(n37174), 
            .O(n14796[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_8 (.CI(n37174), .I0(n15117[5]), .I1(n719), .CO(n37175));
    SB_CARRY add_3097_2 (.CI(GND_net), .I0(n47), .I1(n140_adj_3508), .CO(n38419));
    SB_CARRY add_3251_10 (.CI(n37364), .I0(n12578[7]), .I1(GND_net), .CO(n37365));
    SB_CARRY add_3131_6 (.CI(n37506), .I0(n9932[3]), .I1(n495_adj_3511), 
            .CO(n37507));
    SB_LUT4 add_3382_7_lut (.I0(GND_net), .I1(n15117[4]), .I2(n622), .I3(n37173), 
            .O(n14796[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_9_lut (.I0(GND_net), .I1(n12578[6]), .I2(GND_net), 
            .I3(n37363), .O(n11995[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_19_lut (.I0(GND_net), .I1(n8297[16]), .I2(GND_net), 
            .I3(n38418), .O(n8277[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_7 (.CI(n37173), .I0(n15117[4]), .I1(n622), .CO(n37174));
    SB_CARRY add_3251_9 (.CI(n37363), .I0(n12578[6]), .I1(GND_net), .CO(n37364));
    SB_LUT4 add_3382_6_lut (.I0(GND_net), .I1(n15117[3]), .I2(n525), .I3(n37172), 
            .O(n14796[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i9_1_lut (.I0(\deadband[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[8]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_14_add_1214_7 (.CI(n38733), .I0(n1800[4]), .I1(n448), 
            .CO(n38734));
    SB_LUT4 add_3251_8_lut (.I0(GND_net), .I1(n12578[5]), .I2(n701), .I3(n37362), 
            .O(n11995[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_18_lut (.I0(GND_net), .I1(n8297[15]), .I2(GND_net), 
            .I3(n38417), .O(n8277[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3382_6 (.CI(n37172), .I0(n15117[3]), .I1(n525), .CO(n37173));
    SB_LUT4 add_3382_5_lut (.I0(GND_net), .I1(n15117[2]), .I2(n428), .I3(n37171), 
            .O(n14796[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i8_2_lut (.I0(\Kd[0] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3389));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i8_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3096_18 (.CI(n38417), .I0(n8297[15]), .I1(GND_net), .CO(n38418));
    SB_LUT4 mult_12_i296_2_lut (.I0(\Kd[4] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n440_adj_3564));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i105_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n155));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i105_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i144_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n213));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_6_lut (.I0(GND_net), .I1(n1800[3]), .I2(n375), 
            .I3(n38732), .O(n1799[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_17_lut (.I0(GND_net), .I1(n8297[14]), .I2(GND_net), 
            .I3(n38416), .O(n8277[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1214_6 (.CI(n38732), .I0(n1800[3]), .I1(n375), 
            .CO(n38733));
    SB_LUT4 mult_12_i136_2_lut (.I0(\Kd[2] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n201));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i201_2_lut (.I0(\Kd[3] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n298));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i201_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3096_17 (.CI(n38416), .I0(n8297[14]), .I1(GND_net), .CO(n38417));
    SB_LUT4 add_3131_5_lut (.I0(GND_net), .I1(n9932[2]), .I2(n398_adj_3475), 
            .I3(n37505), .O(n9128[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_8 (.CI(n37362), .I0(n12578[5]), .I1(n701), .CO(n37363));
    SB_LUT4 add_3251_7_lut (.I0(GND_net), .I1(n12578[4]), .I2(n604), .I3(n37361), 
            .O(n11995[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_7 (.CI(n37361), .I0(n12578[4]), .I1(n604), .CO(n37362));
    SB_LUT4 mult_12_i361_2_lut (.I0(\Kd[5] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n537_adj_3562));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3096_16_lut (.I0(GND_net), .I1(n8297[13]), .I2(GND_net), 
            .I3(n38415), .O(n8277[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3251_6_lut (.I0(GND_net), .I1(n12578[3]), .I2(n507), .I3(n37360), 
            .O(n11995[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i426_2_lut (.I0(\Kd[6] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n634_adj_3561));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i426_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3251_6 (.CI(n37360), .I0(n12578[3]), .I1(n507), .CO(n37361));
    SB_CARRY add_3382_5 (.CI(n37171), .I0(n15117[2]), .I1(n428), .CO(n37172));
    SB_LUT4 mult_14_add_1214_5_lut (.I0(GND_net), .I1(n1800[2]), .I2(n302), 
            .I3(n38731), .O(n1799[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i170_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n252));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3382_4_lut (.I0(GND_net), .I1(n15117[1]), .I2(n331), .I3(n37170), 
            .O(n14796[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i209_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n310));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i209_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3096_16 (.CI(n38415), .I0(n8297[13]), .I1(GND_net), .CO(n38416));
    SB_LUT4 mult_12_i491_2_lut (.I0(\Kd[7] ), .I1(n61[17]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_3559));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_17_add_3_3 (.CI(n37007), .I0(GND_net), .I1(n64[1]), 
            .CO(n37008));
    SB_LUT4 add_3251_5_lut (.I0(GND_net), .I1(n12578[2]), .I2(n410_adj_3469), 
            .I3(n37359), .O(n11995[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i266_2_lut (.I0(\Kd[4] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n395));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i331_2_lut (.I0(\Kd[5] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n492));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3096_15_lut (.I0(GND_net), .I1(n8297[12]), .I2(GND_net), 
            .I3(n38414), .O(n8277[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i274_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n407));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i235_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n349));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i235_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3382_4 (.CI(n37170), .I0(n15117[1]), .I1(n331), .CO(n37171));
    SB_CARRY add_3251_5 (.CI(n37359), .I0(n12578[2]), .I1(n410_adj_3469), 
            .CO(n37360));
    SB_LUT4 add_3382_3_lut (.I0(GND_net), .I1(n15117[0]), .I2(n234_adj_3460), 
            .I3(n37169), .O(n14796[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i396_2_lut (.I0(\Kd[6] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n589));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i396_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3131_5 (.CI(n37505), .I0(n9932[2]), .I1(n398_adj_3475), 
            .CO(n37506));
    SB_CARRY add_3096_15 (.CI(n38414), .I0(n8297[12]), .I1(GND_net), .CO(n38415));
    SB_CARRY add_3382_3 (.CI(n37169), .I0(n15117[0]), .I1(n234_adj_3460), 
            .CO(n37170));
    SB_LUT4 unary_minus_17_add_3_2_lut (.I0(n28729), .I1(GND_net), .I2(n64[0]), 
            .I3(VCC_net), .O(n47126)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_17_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3251_4_lut (.I0(GND_net), .I1(n12578[1]), .I2(n313), .I3(n37358), 
            .O(n11995[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_17_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n64[0]), 
            .CO(n37007));
    SB_LUT4 add_3382_2_lut (.I0(GND_net), .I1(n44), .I2(n137_adj_3447), 
            .I3(GND_net), .O(n14796[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3382_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i339_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n504));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i339_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3251_4 (.CI(n37358), .I0(n12578[1]), .I1(n313), .CO(n37359));
    SB_LUT4 add_3131_4_lut (.I0(GND_net), .I1(n9932[1]), .I2(n301_adj_3446), 
            .I3(n37504), .O(n9128[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i461_2_lut (.I0(\Kd[7] ), .I1(n61[2]), .I2(GND_net), 
            .I3(GND_net), .O(n686));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3096_14_lut (.I0(GND_net), .I1(n8297[11]), .I2(GND_net), 
            .I3(n38413), .O(n8277[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_5 (.CI(n38731), .I0(n1800[2]), .I1(n302), 
            .CO(n38732));
    SB_LUT4 add_3251_3_lut (.I0(GND_net), .I1(n12578[0]), .I2(n216), .I3(n37357), 
            .O(n11995[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_3 (.CI(n37357), .I0(n12578[0]), .I1(n216), .CO(n37358));
    SB_CARRY add_3096_14 (.CI(n38413), .I0(n8297[11]), .I1(GND_net), .CO(n38414));
    SB_LUT4 add_3251_2_lut (.I0(GND_net), .I1(n26_adj_3440), .I2(n119), 
            .I3(GND_net), .O(n11995[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3251_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3251_2 (.CI(GND_net), .I0(n26_adj_3440), .I1(n119), .CO(n37357));
    SB_CARRY add_3382_2 (.CI(GND_net), .I0(n44), .I1(n137_adj_3447), .CO(n37169));
    SB_LUT4 mult_14_add_1214_4_lut (.I0(GND_net), .I1(n1800[1]), .I2(n229_adj_3437), 
            .I3(n38730), .O(n1799[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_13_lut (.I0(GND_net), .I1(n8297[10]), .I2(GND_net), 
            .I3(n38412), .O(n8277[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(n37356), .O(n15229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n446));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_9_lut (.I0(GND_net), .I1(n583_adj_3436), .I2(GND_net), 
            .I3(n37355), .O(n15229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n601_adj_3552));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3096_13 (.CI(n38412), .I0(n8297[10]), .I1(GND_net), .CO(n38413));
    SB_LUT4 mult_14_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n698));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3096_12_lut (.I0(GND_net), .I1(n8297[9]), .I2(GND_net), 
            .I3(n38411), .O(n8277[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n543));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i430_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n640));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i430_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i495_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i103_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n152));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i103_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3131_4 (.CI(n37504), .I0(n9932[1]), .I1(n301_adj_3446), 
            .CO(n37505));
    SB_CARRY add_3407_9 (.CI(n37355), .I0(n583_adj_3436), .I1(GND_net), 
            .CO(n37356));
    SB_LUT4 mult_10_i40_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[19] ), 
            .I2(GND_net), .I3(GND_net), .O(n59));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i40_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1214_4 (.CI(n38730), .I0(n1800[1]), .I1(n229_adj_3437), 
            .CO(n38731));
    SB_CARRY add_3096_12 (.CI(n38411), .I0(n8297[9]), .I1(GND_net), .CO(n38412));
    SB_LUT4 mult_10_i168_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n249));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i168_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i233_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n346));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i233_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_8_lut (.I0(GND_net), .I1(n510), .I2(n545), .I3(n37354), 
            .O(n15229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_8 (.CI(n37354), .I0(n510), .I1(n545), .CO(n37355));
    SB_LUT4 mult_12_i73_2_lut (.I0(\Kd[1] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i10_2_lut (.I0(\Kd[0] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_3387));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i138_2_lut (.I0(\Kd[2] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n204));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n443));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i203_2_lut (.I0(\Kd[3] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n301));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i203_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i268_2_lut (.I0(\Kd[4] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n398));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i268_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n540));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i333_2_lut (.I0(\Kd[5] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n495));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i333_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_3_lut (.I0(GND_net), .I1(n1800[0]), .I2(n156_adj_3626), 
            .I3(n38729), .O(n1799[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i398_2_lut (.I0(\Kd[6] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n592));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3096_11_lut (.I0(GND_net), .I1(n8297[8]), .I2(GND_net), 
            .I3(n38410), .O(n8277[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i428_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n637));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i428_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3096_11 (.CI(n38410), .I0(n8297[8]), .I1(GND_net), .CO(n38411));
    SB_CARRY mult_14_add_1214_3 (.CI(n38729), .I0(n1800[0]), .I1(n156_adj_3626), 
            .CO(n38730));
    SB_LUT4 add_3096_10_lut (.I0(GND_net), .I1(n8297[7]), .I2(GND_net), 
            .I3(n38409), .O(n8277[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3131_3_lut (.I0(GND_net), .I1(n9932[0]), .I2(n204_adj_3627), 
            .I3(n37503), .O(n9128[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_7_lut (.I0(GND_net), .I1(n437_adj_3628), .I2(n472), 
            .I3(n37353), .O(n15229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_10 (.CI(n38409), .I0(n8297[7]), .I1(GND_net), .CO(n38410));
    SB_CARRY add_3131_3 (.CI(n37503), .I0(n9932[0]), .I1(n204_adj_3627), 
            .CO(n37504));
    SB_CARRY add_3407_7 (.CI(n37353), .I0(n437_adj_3628), .I1(n472), .CO(n37354));
    SB_LUT4 mult_12_i103_2_lut (.I0(\Kd[1] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n152_adj_3551));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i103_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1214_2_lut (.I0(GND_net), .I1(n14_adj_3629), .I2(n83), 
            .I3(GND_net), .O(n1799[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1214_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_9_lut (.I0(GND_net), .I1(n8297[6]), .I2(GND_net), 
            .I3(n38408), .O(n8277[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_6_lut (.I0(GND_net), .I1(n364_adj_3630), .I2(n399), 
            .I3(n37352), .O(n15229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i463_2_lut (.I0(\Kd[7] ), .I1(n61[3]), .I2(GND_net), 
            .I3(GND_net), .O(n689));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3407_6 (.CI(n37352), .I0(n364_adj_3630), .I1(n399), .CO(n37353));
    SB_LUT4 mult_10_i493_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i101_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n149));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i101_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[18] ), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i40_2_lut (.I0(\Kd[0] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n59_adj_3550));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i40_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[9]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i166_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n246));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i166_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i231_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n343));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n440));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i75_2_lut (.I0(\Kd[1] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i75_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3096_9 (.CI(n38408), .I0(n8297[6]), .I1(GND_net), .CO(n38409));
    SB_LUT4 mult_12_i12_2_lut (.I0(\Kd[0] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3380));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3407_5_lut (.I0(GND_net), .I1(n291), .I2(n326), .I3(n37351), 
            .O(n15229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n537_adj_3379));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i140_2_lut (.I0(\Kd[2] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n207));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3096_8_lut (.I0(GND_net), .I1(n8297[5]), .I2(n719_adj_3632), 
            .I3(n38407), .O(n8277[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1214_2 (.CI(GND_net), .I0(n14_adj_3629), .I1(n83), 
            .CO(n38729));
    SB_CARRY add_3096_8 (.CI(n38407), .I0(n8297[5]), .I1(n719_adj_3632), 
            .CO(n38408));
    SB_LUT4 add_3131_2_lut (.I0(GND_net), .I1(n14_adj_3633), .I2(n107_adj_3634), 
            .I3(GND_net), .O(n9128[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3131_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_5 (.CI(n37351), .I0(n291), .I1(n326), .CO(n37352));
    SB_LUT4 add_3096_7_lut (.I0(GND_net), .I1(n8297[4]), .I2(n622_adj_3635), 
            .I3(n38406), .O(n8277[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3131_2 (.CI(GND_net), .I0(n14_adj_3633), .I1(n107_adj_3634), 
            .CO(n37503));
    SB_LUT4 add_3407_4_lut (.I0(GND_net), .I1(n218_adj_3636), .I2(n253), 
            .I3(n37350), .O(n15229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i205_2_lut (.I0(\Kd[3] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n304));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i205_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3407_4 (.CI(n37350), .I0(n218_adj_3636), .I1(n253), .CO(n37351));
    SB_LUT4 mult_14_add_1213_24_lut (.I0(GND_net), .I1(n1799[21]), .I2(GND_net), 
            .I3(n38727), .O(n1798[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_24 (.CI(n38727), .I0(n1799[21]), .I1(GND_net), 
            .CO(n1691));
    SB_CARRY add_3096_7 (.CI(n38406), .I0(n8297[4]), .I1(n622_adj_3635), 
            .CO(n38407));
    SB_LUT4 add_3096_6_lut (.I0(GND_net), .I1(n8297[3]), .I2(n525_adj_3637), 
            .I3(n38405), .O(n8277[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_3_lut (.I0(GND_net), .I1(n145_adj_3638), .I2(n180), 
            .I3(n37349), .O(n15229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_6 (.CI(n38405), .I0(n8297[3]), .I1(n525_adj_3637), 
            .CO(n38406));
    SB_LUT4 mult_14_add_1213_23_lut (.I0(GND_net), .I1(n1799[20]), .I2(GND_net), 
            .I3(n38726), .O(n1798[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_5_lut (.I0(GND_net), .I1(n8297[2]), .I2(n428_adj_3639), 
            .I3(n38404), .O(n8277[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3407_3 (.CI(n37349), .I0(n145_adj_3638), .I1(n180), .CO(n37350));
    SB_LUT4 add_3329_14_lut (.I0(GND_net), .I1(n14171[11]), .I2(GND_net), 
            .I3(n37502), .O(n13737[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3407_2_lut (.I0(GND_net), .I1(n72), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n15229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3407_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_23 (.CI(n38726), .I0(n1799[20]), .I1(GND_net), 
            .CO(n38727));
    SB_CARRY add_3096_5 (.CI(n38404), .I0(n8297[2]), .I1(n428_adj_3639), 
            .CO(n38405));
    SB_LUT4 add_3329_13_lut (.I0(GND_net), .I1(n14171[10]), .I2(GND_net), 
            .I3(n37501), .O(n13737[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i168_2_lut (.I0(\Kd[2] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n249_adj_3549));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i168_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3329_13 (.CI(n37501), .I0(n14171[10]), .I1(GND_net), 
            .CO(n37502));
    SB_CARRY add_3407_2 (.CI(GND_net), .I0(n72), .I1(n107_adj_3418), .CO(n37349));
    SB_LUT4 mult_14_add_1213_22_lut (.I0(GND_net), .I1(n1799[19]), .I2(GND_net), 
            .I3(n38725), .O(n1798[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_4_lut (.I0(GND_net), .I1(n8297[1]), .I2(n331_adj_3640), 
            .I3(n38403), .O(n8277[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_4 (.CI(n38403), .I0(n8297[1]), .I1(n331_adj_3640), 
            .CO(n38404));
    SB_CARRY mult_14_add_1213_22 (.CI(n38725), .I0(n1799[19]), .I1(GND_net), 
            .CO(n38726));
    SB_LUT4 add_3276_24_lut (.I0(GND_net), .I1(n13112[21]), .I2(GND_net), 
            .I3(n37348), .O(n12578[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_3_lut (.I0(GND_net), .I1(n8297[0]), .I2(n234_adj_3641), 
            .I3(n38402), .O(n8277[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3329_12_lut (.I0(GND_net), .I1(n14171[9]), .I2(GND_net), 
            .I3(n37500), .O(n13737[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_3 (.CI(n38402), .I0(n8297[0]), .I1(n234_adj_3641), 
            .CO(n38403));
    SB_LUT4 add_3276_23_lut (.I0(GND_net), .I1(n13112[20]), .I2(GND_net), 
            .I3(n37347), .O(n12578[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_12 (.CI(n37500), .I0(n14171[9]), .I1(GND_net), .CO(n37501));
    SB_CARRY add_3276_23 (.CI(n37347), .I0(n13112[20]), .I1(GND_net), 
            .CO(n37348));
    SB_LUT4 add_3276_22_lut (.I0(GND_net), .I1(n13112[19]), .I2(GND_net), 
            .I3(n37346), .O(n12578[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3096_2_lut (.I0(GND_net), .I1(n44_adj_3642), .I2(n137_adj_3643), 
            .I3(GND_net), .O(n8277[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3096_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_21_lut (.I0(GND_net), .I1(n1799[18]), .I2(GND_net), 
            .I3(n38724), .O(n1798[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3096_2 (.CI(GND_net), .I0(n44_adj_3642), .I1(n137_adj_3643), 
            .CO(n38402));
    SB_CARRY add_3276_22 (.CI(n37346), .I0(n13112[19]), .I1(GND_net), 
            .CO(n37347));
    SB_LUT4 add_3329_11_lut (.I0(GND_net), .I1(n14171[8]), .I2(GND_net), 
            .I3(n37499), .O(n13737[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_21_lut (.I0(GND_net), .I1(n13112[18]), .I2(GND_net), 
            .I3(n37345), .O(n12578[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i233_2_lut (.I0(\Kd[3] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n346_adj_3548));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i233_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1213_21 (.CI(n38724), .I0(n1799[18]), .I1(GND_net), 
            .CO(n38725));
    SB_LUT4 mult_14_add_1213_20_lut (.I0(GND_net), .I1(n1799[17]), .I2(GND_net), 
            .I3(n38723), .O(n1798[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i426_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n634));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i426_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3329_11 (.CI(n37499), .I0(n14171[8]), .I1(GND_net), .CO(n37500));
    SB_LUT4 mult_12_i298_2_lut (.I0(\Kd[4] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n443_adj_3547));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1213_20 (.CI(n38723), .I0(n1799[17]), .I1(GND_net), 
            .CO(n38724));
    SB_LUT4 add_3095_20_lut (.I0(GND_net), .I1(n8277[17]), .I2(GND_net), 
            .I3(n38401), .O(n8256[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_21 (.CI(n37345), .I0(n13112[18]), .I1(GND_net), 
            .CO(n37346));
    SB_LUT4 add_3276_20_lut (.I0(GND_net), .I1(n13112[17]), .I2(GND_net), 
            .I3(n37344), .O(n12578[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_19_lut (.I0(GND_net), .I1(n8277[16]), .I2(GND_net), 
            .I3(n38400), .O(n8256[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_20 (.CI(n37344), .I0(n13112[17]), .I1(GND_net), 
            .CO(n37345));
    SB_LUT4 mult_12_i363_2_lut (.I0(\Kd[5] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n540_adj_3545));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i270_2_lut (.I0(\Kd[4] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n401));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3276_19_lut (.I0(GND_net), .I1(n13112[16]), .I2(GND_net), 
            .I3(n37343), .O(n12578[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_19 (.CI(n37343), .I0(n13112[16]), .I1(GND_net), 
            .CO(n37344));
    SB_LUT4 add_3276_18_lut (.I0(GND_net), .I1(n13112[15]), .I2(GND_net), 
            .I3(n37342), .O(n12578[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_19_lut (.I0(GND_net), .I1(n1799[16]), .I2(GND_net), 
            .I3(n38722), .O(n1798[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_19 (.CI(n38400), .I0(n8277[16]), .I1(GND_net), .CO(n38401));
    SB_LUT4 add_3095_18_lut (.I0(GND_net), .I1(n8277[15]), .I2(GND_net), 
            .I3(n38399), .O(n8256[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_19 (.CI(n38722), .I0(n1799[16]), .I1(GND_net), 
            .CO(n38723));
    SB_CARRY add_3095_18 (.CI(n38399), .I0(n8277[15]), .I1(GND_net), .CO(n38400));
    SB_LUT4 add_3329_10_lut (.I0(GND_net), .I1(n14171[7]), .I2(GND_net), 
            .I3(n37498), .O(n13737[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_18 (.CI(n37342), .I0(n13112[15]), .I1(GND_net), 
            .CO(n37343));
    SB_LUT4 add_3095_17_lut (.I0(GND_net), .I1(n8277[14]), .I2(GND_net), 
            .I3(n38398), .O(n8256[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_10 (.CI(n37498), .I0(n14171[7]), .I1(GND_net), .CO(n37499));
    SB_LUT4 add_3276_17_lut (.I0(GND_net), .I1(n13112[14]), .I2(GND_net), 
            .I3(n37341), .O(n12578[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_18_lut (.I0(GND_net), .I1(n1799[15]), .I2(GND_net), 
            .I3(n38721), .O(n1798[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_18 (.CI(n38721), .I0(n1799[15]), .I1(GND_net), 
            .CO(n38722));
    SB_CARRY add_3095_17 (.CI(n38398), .I0(n8277[14]), .I1(GND_net), .CO(n38399));
    SB_LUT4 add_3095_16_lut (.I0(GND_net), .I1(n8277[13]), .I2(GND_net), 
            .I3(n38397), .O(n8256[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_16 (.CI(n38397), .I0(n8277[13]), .I1(GND_net), .CO(n38398));
    SB_LUT4 mult_14_add_1213_17_lut (.I0(GND_net), .I1(n1799[14]), .I2(GND_net), 
            .I3(n38720), .O(n1798[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_15_lut (.I0(GND_net), .I1(n8277[12]), .I2(GND_net), 
            .I3(n38396), .O(n8256[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3329_9_lut (.I0(GND_net), .I1(n14171[6]), .I2(GND_net), 
            .I3(n37497), .O(n13737[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_17 (.CI(n37341), .I0(n13112[14]), .I1(GND_net), 
            .CO(n37342));
    SB_CARRY add_3095_15 (.CI(n38396), .I0(n8277[12]), .I1(GND_net), .CO(n38397));
    SB_CARRY add_3329_9 (.CI(n37497), .I0(n14171[6]), .I1(GND_net), .CO(n37498));
    SB_LUT4 add_3276_16_lut (.I0(GND_net), .I1(n13112[13]), .I2(GND_net), 
            .I3(n37340), .O(n12578[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_17 (.CI(n38720), .I0(n1799[14]), .I1(GND_net), 
            .CO(n38721));
    SB_LUT4 add_3095_14_lut (.I0(GND_net), .I1(n8277[11]), .I2(GND_net), 
            .I3(n38395), .O(n8256[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_16 (.CI(n37340), .I0(n13112[13]), .I1(GND_net), 
            .CO(n37341));
    SB_LUT4 add_3276_15_lut (.I0(GND_net), .I1(n13112[12]), .I2(GND_net), 
            .I3(n37339), .O(n12578[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_26_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n75[23]), .I3(n37145), .O(\PID_CONTROLLER.err_31__N_2816 [24])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_14 (.CI(n38395), .I0(n8277[11]), .I1(GND_net), .CO(n38396));
    SB_CARRY add_3276_15 (.CI(n37339), .I0(n13112[12]), .I1(GND_net), 
            .CO(n37340));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(\motor_state[23] ), 
            .I2(n75[23]), .I3(n37144), .O(\PID_CONTROLLER.err_31__N_2816 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_25 (.CI(n37144), .I0(\motor_state[23] ), 
            .I1(n75[23]), .CO(n37145));
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(\motor_state[22] ), 
            .I2(n75[22]), .I3(n37143), .O(\PID_CONTROLLER.err_31__N_2816 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n37143), .I0(\motor_state[22] ), 
            .I1(n75[22]), .CO(n37144));
    SB_DFFE \PID_CONTROLLER.integral_1048__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[0]));   // verilog/motorControl.v(34[21:33])
    SB_LUT4 add_3095_13_lut (.I0(GND_net), .I1(n8277[10]), .I2(GND_net), 
            .I3(n38394), .O(n8256[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_16_lut (.I0(GND_net), .I1(n1799[13]), .I2(GND_net), 
            .I3(n38719), .O(n1798[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i428_2_lut (.I0(\Kd[6] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n637_adj_3544));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i428_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3329_8_lut (.I0(GND_net), .I1(n14171[5]), .I2(n545), .I3(n37496), 
            .O(n13737[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i493_2_lut (.I0(\Kd[7] ), .I1(n61[18]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_3543));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i493_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3276_14_lut (.I0(GND_net), .I1(n13112[11]), .I2(GND_net), 
            .I3(n37338), .O(n12578[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(\motor_state[21] ), 
            .I2(n75[21]), .I3(n37142), .O(\PID_CONTROLLER.err_31__N_2816 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n37142), .I0(\motor_state[21] ), 
            .I1(n75[21]), .CO(n37143));
    SB_LUT4 mult_12_i335_2_lut (.I0(\Kd[5] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n498));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i335_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1213_16 (.CI(n38719), .I0(n1799[13]), .I1(GND_net), 
            .CO(n38720));
    SB_CARRY add_3095_13 (.CI(n38394), .I0(n8277[10]), .I1(GND_net), .CO(n38395));
    SB_CARRY add_3276_14 (.CI(n37338), .I0(n13112[11]), .I1(GND_net), 
            .CO(n37339));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(\motor_state[20] ), 
            .I2(n75[20]), .I3(n37141), .O(\PID_CONTROLLER.err_31__N_2816 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n37141), .I0(\motor_state[20] ), 
            .I1(n75[20]), .CO(n37142));
    SB_LUT4 add_3276_13_lut (.I0(GND_net), .I1(n13112[10]), .I2(GND_net), 
            .I3(n37337), .O(n12578[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(\motor_state[19] ), 
            .I2(n75[19]), .I3(n37140), .O(\PID_CONTROLLER.err_31__N_2816 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n37140), .I0(\motor_state[19] ), 
            .I1(n75[19]), .CO(n37141));
    SB_LUT4 add_3095_12_lut (.I0(GND_net), .I1(n8277[9]), .I2(GND_net), 
            .I3(n38393), .O(n8256[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_13 (.CI(n37337), .I0(n13112[10]), .I1(GND_net), 
            .CO(n37338));
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(\motor_state[18] ), 
            .I2(n75[18]), .I3(n37139), .O(\PID_CONTROLLER.err_31__N_2816 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n37139), .I0(\motor_state[18] ), 
            .I1(n75[18]), .CO(n37140));
    SB_LUT4 mult_14_add_1213_15_lut (.I0(GND_net), .I1(n1799[12]), .I2(GND_net), 
            .I3(n38718), .O(n1798[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_12 (.CI(n38393), .I0(n8277[9]), .I1(GND_net), .CO(n38394));
    SB_LUT4 add_3095_11_lut (.I0(GND_net), .I1(n8277[8]), .I2(GND_net), 
            .I3(n38392), .O(n8256[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_15 (.CI(n38718), .I0(n1799[12]), .I1(GND_net), 
            .CO(n38719));
    SB_LUT4 mult_10_i491_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i491_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i400_2_lut (.I0(\Kd[6] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n595));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3095_11 (.CI(n38392), .I0(n8277[8]), .I1(GND_net), .CO(n38393));
    SB_LUT4 add_3276_12_lut (.I0(GND_net), .I1(n13112[9]), .I2(GND_net), 
            .I3(n37336), .O(n12578[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(\motor_state[17] ), 
            .I2(n75[17]), .I3(n37138), .O(\PID_CONTROLLER.err_31__N_2816 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n37138), .I0(\motor_state[17] ), 
            .I1(n75[17]), .CO(n37139));
    SB_CARRY add_3329_8 (.CI(n37496), .I0(n14171[5]), .I1(n545), .CO(n37497));
    SB_LUT4 mult_14_add_1213_14_lut (.I0(GND_net), .I1(n1799[11]), .I2(GND_net), 
            .I3(n38717), .O(n1798[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_10_lut (.I0(GND_net), .I1(n8277[7]), .I2(GND_net), 
            .I3(n38391), .O(n8256[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_12 (.CI(n37336), .I0(n13112[9]), .I1(GND_net), .CO(n37337));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(\motor_state[16] ), 
            .I2(n75[16]), .I3(n37137), .O(\PID_CONTROLLER.err_31__N_2816 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_11_lut (.I0(GND_net), .I1(n13112[8]), .I2(GND_net), 
            .I3(n37335), .O(n12578[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_11 (.CI(n37335), .I0(n13112[8]), .I1(GND_net), .CO(n37336));
    SB_CARRY state_23__I_0_add_2_18 (.CI(n37137), .I0(\motor_state[16] ), 
            .I1(n75[16]), .CO(n37138));
    SB_CARRY add_3095_10 (.CI(n38391), .I0(n8277[7]), .I1(GND_net), .CO(n38392));
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(\motor_state[15] ), 
            .I2(n75[15]), .I3(n37136), .O(\PID_CONTROLLER.err_31__N_2816 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_9_lut (.I0(GND_net), .I1(n8277[6]), .I2(GND_net), 
            .I3(n38390), .O(n8256[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n37136), .I0(\motor_state[15] ), 
            .I1(n75[15]), .CO(n37137));
    SB_LUT4 add_3329_7_lut (.I0(GND_net), .I1(n14171[4]), .I2(n472), .I3(n37495), 
            .O(n13737[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_10_lut (.I0(GND_net), .I1(n13112[7]), .I2(GND_net), 
            .I3(n37334), .O(n12578[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(\motor_state[14] ), 
            .I2(n75[14]), .I3(n37135), .O(\PID_CONTROLLER.err_31__N_2816 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_16 (.CI(n37135), .I0(\motor_state[14] ), 
            .I1(n75[14]), .CO(n37136));
    SB_CARRY mult_14_add_1213_14 (.CI(n38717), .I0(n1799[11]), .I1(GND_net), 
            .CO(n38718));
    SB_CARRY add_3095_9 (.CI(n38390), .I0(n8277[6]), .I1(GND_net), .CO(n38391));
    SB_LUT4 add_3095_8_lut (.I0(GND_net), .I1(n8277[5]), .I2(n716), .I3(n38389), 
            .O(n8256[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_13_lut (.I0(GND_net), .I1(n1799[10]), .I2(GND_net), 
            .I3(n38716), .O(n1798[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_8 (.CI(n38389), .I0(n8277[5]), .I1(n716), .CO(n38390));
    SB_LUT4 mult_12_i465_2_lut (.I0(\Kd[7] ), .I1(n61[4]), .I2(GND_net), 
            .I3(GND_net), .O(n692));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1213_13 (.CI(n38716), .I0(n1799[10]), .I1(GND_net), 
            .CO(n38717));
    SB_LUT4 mult_10_i111_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3095_7_lut (.I0(GND_net), .I1(n8277[4]), .I2(n619_adj_3655), 
            .I3(n38388), .O(n8256[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i48_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n71));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i48_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3276_10 (.CI(n37334), .I0(n13112[7]), .I1(GND_net), .CO(n37335));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(\motor_state[13] ), 
            .I2(n75[13]), .I3(n37134), .O(\PID_CONTROLLER.err_31__N_2816 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_7 (.CI(n37495), .I0(n14171[4]), .I1(n472), .CO(n37496));
    SB_LUT4 add_3276_9_lut (.I0(GND_net), .I1(n13112[6]), .I2(GND_net), 
            .I3(n37333), .O(n12578[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n37134), .I0(\motor_state[13] ), 
            .I1(n75[13]), .CO(n37135));
    SB_CARRY add_3276_9 (.CI(n37333), .I0(n13112[6]), .I1(GND_net), .CO(n37334));
    SB_LUT4 mult_10_i176_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n261));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[10]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(\motor_state[12] ), 
            .I2(n75[12]), .I3(n37133), .O(\PID_CONTROLLER.err_31__N_2816 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i241_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n358));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n455_c));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n552));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3095_7 (.CI(n38388), .I0(n8277[4]), .I1(n619_adj_3655), 
            .CO(n38389));
    SB_LUT4 mult_14_add_1213_12_lut (.I0(GND_net), .I1(n1799[9]), .I2(GND_net), 
            .I3(n38715), .O(n1798[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i436_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n649));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3095_6_lut (.I0(GND_net), .I1(n8277[3]), .I2(n522_adj_3658), 
            .I3(n38387), .O(n8256[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3329_6_lut (.I0(GND_net), .I1(n14171[3]), .I2(n399), .I3(n37494), 
            .O(n13737[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[11]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3276_8_lut (.I0(GND_net), .I1(n13112[5]), .I2(n704), .I3(n37332), 
            .O(n12578[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n37133), .I0(\motor_state[12] ), 
            .I1(n75[12]), .CO(n37134));
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(\motor_state[11] ), 
            .I2(n75[11]), .I3(n37132), .O(\PID_CONTROLLER.err_31__N_2816 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_8 (.CI(n37332), .I0(n13112[5]), .I1(n704), .CO(n37333));
    SB_CARRY mult_14_add_1213_12 (.CI(n38715), .I0(n1799[9]), .I1(GND_net), 
            .CO(n38716));
    SB_LUT4 mult_10_i501_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3276_7_lut (.I0(GND_net), .I1(n13112[4]), .I2(n607_adj_3660), 
            .I3(n37331), .O(n12578[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n37132), .I0(\motor_state[11] ), 
            .I1(n75[11]), .CO(n37133));
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(\motor_state[10] ), 
            .I2(n75[10]), .I3(n37131), .O(\PID_CONTROLLER.err_31__N_2816 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_7 (.CI(n37331), .I0(n13112[4]), .I1(n607_adj_3660), 
            .CO(n37332));
    SB_CARRY state_23__I_0_add_2_12 (.CI(n37131), .I0(\motor_state[10] ), 
            .I1(n75[10]), .CO(n37132));
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(\motor_state[9] ), 
            .I2(n75[9]), .I3(n37130), .O(\PID_CONTROLLER.err_31__N_2816 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_6 (.CI(n38387), .I0(n8277[3]), .I1(n522_adj_3658), 
            .CO(n38388));
    SB_LUT4 mult_14_add_1213_11_lut (.I0(GND_net), .I1(n1799[8]), .I2(GND_net), 
            .I3(n38714), .O(n1798[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_6_lut (.I0(GND_net), .I1(n13112[3]), .I2(n510_adj_3663), 
            .I3(n37330), .O(n12578[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_5_lut (.I0(GND_net), .I1(n8277[2]), .I2(n425_adj_3664), 
            .I3(n38386), .O(n8256[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n37130), .I0(\motor_state[9] ), 
            .I1(n75[9]), .CO(n37131));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(\motor_state[8] ), 
            .I2(n75[8]), .I3(n37129), .O(\PID_CONTROLLER.err_31__N_2816 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_6 (.CI(n37330), .I0(n13112[3]), .I1(n510_adj_3663), 
            .CO(n37331));
    SB_CARRY mult_14_add_1213_11 (.CI(n38714), .I0(n1799[8]), .I1(GND_net), 
            .CO(n38715));
    SB_CARRY add_3095_5 (.CI(n38386), .I0(n8277[2]), .I1(n425_adj_3664), 
            .CO(n38387));
    SB_CARRY state_23__I_0_add_2_10 (.CI(n37129), .I0(\motor_state[8] ), 
            .I1(n75[8]), .CO(n37130));
    SB_LUT4 add_3276_5_lut (.I0(GND_net), .I1(n13112[2]), .I2(n413_adj_3666), 
            .I3(n37329), .O(n12578[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(\motor_state[7] ), 
            .I2(n75[7]), .I3(n37128), .O(\PID_CONTROLLER.err_31__N_2816 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_10_lut (.I0(GND_net), .I1(n1799[7]), .I2(GND_net), 
            .I3(n38713), .O(n1798[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_10 (.CI(n38713), .I0(n1799[7]), .I1(GND_net), 
            .CO(n38714));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n37128), .I0(\motor_state[7] ), 
            .I1(n75[7]), .CO(n37129));
    SB_LUT4 mult_14_add_1213_9_lut (.I0(GND_net), .I1(n1799[6]), .I2(GND_net), 
            .I3(n38712), .O(n1798[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3095_4_lut (.I0(GND_net), .I1(n8277[1]), .I2(n328_adj_3669), 
            .I3(n38385), .O(n8256[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3276_5 (.CI(n37329), .I0(n13112[2]), .I1(n413_adj_3666), 
            .CO(n37330));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(\motor_state[6] ), 
            .I2(n75[6]), .I3(n37127), .O(\PID_CONTROLLER.err_31__N_2816 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_4_lut (.I0(GND_net), .I1(n13112[1]), .I2(n316_adj_3671), 
            .I3(n37328), .O(n12578[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n37127), .I0(\motor_state[6] ), 
            .I1(n75[6]), .CO(n37128));
    SB_CARRY add_3095_4 (.CI(n38385), .I0(n8277[1]), .I1(n328_adj_3669), 
            .CO(n38386));
    SB_CARRY add_3276_4 (.CI(n37328), .I0(n13112[1]), .I1(n316_adj_3671), 
            .CO(n37329));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(\motor_state[5] ), 
            .I2(n75[5]), .I3(n37126), .O(\PID_CONTROLLER.err_31__N_2816 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_3_lut (.I0(GND_net), .I1(n13112[0]), .I2(n219_adj_3673), 
            .I3(n37327), .O(n12578[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n37126), .I0(\motor_state[5] ), 
            .I1(n75[5]), .CO(n37127));
    SB_CARRY mult_14_add_1213_9 (.CI(n38712), .I0(n1799[6]), .I1(GND_net), 
            .CO(n38713));
    SB_LUT4 add_3095_3_lut (.I0(GND_net), .I1(n8277[0]), .I2(n231_adj_3674), 
            .I3(n38384), .O(n8256[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(\motor_state[4] ), 
            .I2(n75[4]), .I3(n37125), .O(\PID_CONTROLLER.err_31__N_2816 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_8_lut (.I0(GND_net), .I1(n1799[5]), .I2(n518), 
            .I3(n38711), .O(n1798[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[12]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3276_3 (.CI(n37327), .I0(n13112[0]), .I1(n219_adj_3673), 
            .CO(n37328));
    SB_CARRY state_23__I_0_add_2_6 (.CI(n37125), .I0(\motor_state[4] ), 
            .I1(n75[4]), .CO(n37126));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(\motor_state[3] ), 
            .I2(n75[3]), .I3(n37124), .O(\PID_CONTROLLER.err_31__N_2816 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3276_2_lut (.I0(GND_net), .I1(n29_adj_3677), .I2(n122), 
            .I3(GND_net), .O(n12578[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3276_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n37124), .I0(\motor_state[3] ), 
            .I1(n75[3]), .CO(n37125));
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[13]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(\motor_state[2] ), 
            .I2(n75[2]), .I3(n37123), .O(\PID_CONTROLLER.err_31__N_2816 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3095_3 (.CI(n38384), .I0(n8277[0]), .I1(n231_adj_3674), 
            .CO(n38385));
    SB_CARRY add_3276_2 (.CI(GND_net), .I0(n29_adj_3677), .I1(n122), .CO(n37327));
    SB_CARRY state_23__I_0_add_2_4 (.CI(n37123), .I0(\motor_state[2] ), 
            .I1(n75[2]), .CO(n37124));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(\motor_state[1] ), 
            .I2(n75[1]), .I3(n37122), .O(\PID_CONTROLLER.err_31__N_2816 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i91_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n134));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[13] ), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[14]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i156_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n231));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3482_12_lut (.I0(GND_net), .I1(n16423[9]), .I2(GND_net), 
            .I3(n37326), .O(n16317[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n37122), .I0(\motor_state[1] ), 
            .I1(n75[1]), .CO(n37123));
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(\motor_state[0] ), 
            .I2(n75[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_31__N_2816 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_8 (.CI(n38711), .I0(n1799[5]), .I1(n518), 
            .CO(n38712));
    SB_LUT4 add_3095_2_lut (.I0(GND_net), .I1(n41_adj_3681), .I2(n134_adj_3682), 
            .I3(GND_net), .O(n8256[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3095_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3482_11_lut (.I0(GND_net), .I1(n16423[8]), .I2(GND_net), 
            .I3(n37325), .O(n16317[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(\motor_state[0] ), 
            .I1(n75[0]), .CO(n37122));
    SB_LUT4 mult_14_add_1213_7_lut (.I0(GND_net), .I1(n1799[4]), .I2(n445), 
            .I3(n38710), .O(n1798[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_11 (.CI(n37325), .I0(n16423[8]), .I1(GND_net), .CO(n37326));
    SB_LUT4 add_3482_10_lut (.I0(GND_net), .I1(n16423[7]), .I2(GND_net), 
            .I3(n37324), .O(n16317[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_10 (.CI(n37324), .I0(n16423[7]), .I1(GND_net), .CO(n37325));
    SB_CARRY add_3095_2 (.CI(GND_net), .I0(n41_adj_3681), .I1(n134_adj_3682), 
            .CO(n38384));
    SB_LUT4 add_3482_9_lut (.I0(GND_net), .I1(n16423[6]), .I2(GND_net), 
            .I3(n37323), .O(n16317[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_9 (.CI(n37323), .I0(n16423[6]), .I1(GND_net), .CO(n37324));
    SB_CARRY mult_14_add_1213_7 (.CI(n38710), .I0(n1799[4]), .I1(n445), 
            .CO(n38711));
    SB_LUT4 add_3094_21_lut (.I0(GND_net), .I1(n8256[18]), .I2(GND_net), 
            .I3(n38383), .O(n8234[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_20_lut (.I0(GND_net), .I1(n8256[17]), .I2(GND_net), 
            .I3(n38382), .O(n8234[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_20 (.CI(n38382), .I0(n8256[17]), .I1(GND_net), .CO(n38383));
    SB_LUT4 add_3094_19_lut (.I0(GND_net), .I1(n8256[16]), .I2(GND_net), 
            .I3(n38381), .O(n8234[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_19 (.CI(n38381), .I0(n8256[16]), .I1(GND_net), .CO(n38382));
    SB_LUT4 add_3482_8_lut (.I0(GND_net), .I1(n16423[5]), .I2(n740_adj_3684), 
            .I3(n37322), .O(n16317[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_8 (.CI(n37322), .I0(n16423[5]), .I1(n740_adj_3684), 
            .CO(n37323));
    SB_LUT4 add_3482_7_lut (.I0(GND_net), .I1(n16423[4]), .I2(n643_adj_3685), 
            .I3(n37321), .O(n16317[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_7 (.CI(n37321), .I0(n16423[4]), .I1(n643_adj_3685), 
            .CO(n37322));
    SB_LUT4 mult_14_add_1213_6_lut (.I0(GND_net), .I1(n1799[3]), .I2(n372), 
            .I3(n38709), .O(n1798[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_18_lut (.I0(GND_net), .I1(n8256[15]), .I2(GND_net), 
            .I3(n38380), .O(n8234[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3482_6_lut (.I0(GND_net), .I1(n16423[3]), .I2(n546_adj_3686), 
            .I3(n37320), .O(n16317[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3482_6 (.CI(n37320), .I0(n16423[3]), .I1(n546_adj_3686), 
            .CO(n37321));
    SB_CARRY mult_14_add_1213_6 (.CI(n38709), .I0(n1799[3]), .I1(n372), 
            .CO(n38710));
    SB_LUT4 mult_14_add_1213_5_lut (.I0(GND_net), .I1(n1799[2]), .I2(n299_adj_3688), 
            .I3(n38708), .O(n1798[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_18 (.CI(n38380), .I0(n8256[15]), .I1(GND_net), .CO(n38381));
    SB_LUT4 add_3482_5_lut (.I0(GND_net), .I1(n16423[2]), .I2(n449_adj_3689), 
            .I3(n37319), .O(n16317[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_5 (.CI(n38708), .I0(n1799[2]), .I1(n299_adj_3688), 
            .CO(n38709));
    SB_LUT4 add_3094_17_lut (.I0(GND_net), .I1(n8256[14]), .I2(GND_net), 
            .I3(n38379), .O(n8234[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_6 (.CI(n37494), .I0(n14171[3]), .I1(n399), .CO(n37495));
    SB_CARRY add_3482_5 (.CI(n37319), .I0(n16423[2]), .I1(n449_adj_3689), 
            .CO(n37320));
    SB_LUT4 add_3329_5_lut (.I0(GND_net), .I1(n14171[2]), .I2(n326), .I3(n37493), 
            .O(n13737[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1213_4_lut (.I0(GND_net), .I1(n1799[1]), .I2(n226_adj_3691), 
            .I3(n38707), .O(n1798[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3482_4_lut (.I0(GND_net), .I1(n16423[1]), .I2(n352_adj_3692), 
            .I3(n37318), .O(n16317[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_5 (.CI(n37493), .I0(n14171[2]), .I1(n326), .CO(n37494));
    SB_CARRY add_3094_17 (.CI(n38379), .I0(n8256[14]), .I1(GND_net), .CO(n38380));
    SB_CARRY mult_14_add_1213_4 (.CI(n38707), .I0(n1799[1]), .I1(n226_adj_3691), 
            .CO(n38708));
    SB_LUT4 mult_14_add_1213_3_lut (.I0(GND_net), .I1(n1799[0]), .I2(n153_adj_3694), 
            .I3(n38706), .O(n1798[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i221_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n328));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i115_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n182));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i50_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i50_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3482_4 (.CI(n37318), .I0(n16423[1]), .I1(n352_adj_3692), 
            .CO(n37319));
    SB_LUT4 add_3482_3_lut (.I0(GND_net), .I1(n16423[0]), .I2(n255_adj_3695), 
            .I3(n37317), .O(n16317[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_16_lut (.I0(GND_net), .I1(n8256[13]), .I2(GND_net), 
            .I3(n38378), .O(n8234[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_3 (.CI(n38706), .I0(n1799[0]), .I1(n153_adj_3694), 
            .CO(n38707));
    SB_CARRY add_3094_16 (.CI(n38378), .I0(n8256[13]), .I1(GND_net), .CO(n38379));
    SB_CARRY add_3482_3 (.CI(n37317), .I0(n16423[0]), .I1(n255_adj_3695), 
            .CO(n37318));
    SB_LUT4 add_3094_15_lut (.I0(GND_net), .I1(n8256[12]), .I2(GND_net), 
            .I3(n38377), .O(n8234[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3482_2_lut (.I0(GND_net), .I1(n65_adj_3696), .I2(n158_adj_3697), 
            .I3(GND_net), .O(n16317[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3482_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i180_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n276));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i46_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i245_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n370));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n464_adj_3377));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3482_2 (.CI(GND_net), .I0(n65_adj_3696), .I1(n158_adj_3697), 
            .CO(n37317));
    SB_LUT4 mult_14_add_1213_2_lut (.I0(GND_net), .I1(n11_adj_3698), .I2(n80), 
            .I3(GND_net), .O(n1798[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1213_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_15 (.CI(n38377), .I0(n8256[12]), .I1(GND_net), .CO(n38378));
    SB_LUT4 add_3300_23_lut (.I0(GND_net), .I1(n13597[20]), .I2(GND_net), 
            .I3(n37316), .O(n13112[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3300_22_lut (.I0(GND_net), .I1(n13597[19]), .I2(GND_net), 
            .I3(n37315), .O(n13112[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_14_lut (.I0(GND_net), .I1(n8256[11]), .I2(GND_net), 
            .I3(n38376), .O(n8234[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_22 (.CI(n37315), .I0(n13597[19]), .I1(GND_net), 
            .CO(n37316));
    SB_LUT4 add_3300_21_lut (.I0(GND_net), .I1(n13597[18]), .I2(GND_net), 
            .I3(n37314), .O(n13112[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1213_2 (.CI(GND_net), .I0(n11_adj_3698), .I1(n80), 
            .CO(n38706));
    SB_CARRY add_3094_14 (.CI(n38376), .I0(n8256[11]), .I1(GND_net), .CO(n38377));
    SB_CARRY add_3300_21 (.CI(n37314), .I0(n13597[18]), .I1(GND_net), 
            .CO(n37315));
    SB_LUT4 add_3300_20_lut (.I0(GND_net), .I1(n13597[17]), .I2(GND_net), 
            .I3(n37313), .O(n13112[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_13_lut (.I0(GND_net), .I1(n8256[10]), .I2(GND_net), 
            .I3(n38375), .O(n8234[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_20 (.CI(n37313), .I0(n13597[17]), .I1(GND_net), 
            .CO(n37314));
    SB_LUT4 add_3300_19_lut (.I0(GND_net), .I1(n13597[16]), .I2(GND_net), 
            .I3(n37312), .O(n13112[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i61_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3300_19 (.CI(n37312), .I0(n13597[16]), .I1(GND_net), 
            .CO(n37313));
    SB_LUT4 mult_14_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3541));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1212_24_lut (.I0(GND_net), .I1(n1798[21]), .I2(GND_net), 
            .I3(n38704), .O(n1797[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_13 (.CI(n38375), .I0(n8256[10]), .I1(GND_net), .CO(n38376));
    SB_LUT4 add_3300_18_lut (.I0(GND_net), .I1(n13597[15]), .I2(GND_net), 
            .I3(n37311), .O(n13112[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_18 (.CI(n37311), .I0(n13597[15]), .I1(GND_net), 
            .CO(n37312));
    SB_LUT4 add_3094_12_lut (.I0(GND_net), .I1(n8256[9]), .I2(GND_net), 
            .I3(n38374), .O(n8234[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3300_17_lut (.I0(GND_net), .I1(n13597[14]), .I2(GND_net), 
            .I3(n37310), .O(n13112[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_17 (.CI(n37310), .I0(n13597[14]), .I1(GND_net), 
            .CO(n37311));
    SB_CARRY mult_14_add_1212_24 (.CI(n38704), .I0(n1798[21]), .I1(GND_net), 
            .CO(n1687));
    SB_CARRY add_3094_12 (.CI(n38374), .I0(n8256[9]), .I1(GND_net), .CO(n38375));
    SB_LUT4 add_3300_16_lut (.I0(GND_net), .I1(n13597[13]), .I2(GND_net), 
            .I3(n37309), .O(n13112[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_16 (.CI(n37309), .I0(n13597[13]), .I1(GND_net), 
            .CO(n37310));
    SB_LUT4 add_3094_11_lut (.I0(GND_net), .I1(n8256[8]), .I2(GND_net), 
            .I3(n38373), .O(n8234[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3300_15_lut (.I0(GND_net), .I1(n13597[12]), .I2(GND_net), 
            .I3(n37308), .O(n13112[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_15 (.CI(n37308), .I0(n13597[12]), .I1(GND_net), 
            .CO(n37309));
    SB_LUT4 add_3300_14_lut (.I0(GND_net), .I1(n13597[11]), .I2(GND_net), 
            .I3(n37307), .O(n13112[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n558));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1212_23_lut (.I0(GND_net), .I1(n1798[20]), .I2(GND_net), 
            .I3(n38703), .O(n1797[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_11 (.CI(n38373), .I0(n8256[8]), .I1(GND_net), .CO(n38374));
    SB_CARRY add_3300_14 (.CI(n37307), .I0(n13597[11]), .I1(GND_net), 
            .CO(n37308));
    SB_LUT4 add_3300_13_lut (.I0(GND_net), .I1(n13597[10]), .I2(GND_net), 
            .I3(n37306), .O(n13112[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_10_lut (.I0(GND_net), .I1(n8256[7]), .I2(GND_net), 
            .I3(n38372), .O(n8234[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3329_4_lut (.I0(GND_net), .I1(n14171[1]), .I2(n253), .I3(n37492), 
            .O(n13737[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_13 (.CI(n37306), .I0(n13597[10]), .I1(GND_net), 
            .CO(n37307));
    SB_LUT4 mult_14_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_3538));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3300_12_lut (.I0(GND_net), .I1(n13597[9]), .I2(GND_net), 
            .I3(n37305), .O(n13112[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_12 (.CI(n37305), .I0(n13597[9]), .I1(GND_net), .CO(n37306));
    SB_LUT4 mult_14_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_14_add_1212_23 (.CI(n38703), .I0(n1798[20]), .I1(GND_net), 
            .CO(n38704));
    SB_CARRY add_3094_10 (.CI(n38372), .I0(n8256[7]), .I1(GND_net), .CO(n38373));
    SB_LUT4 add_3300_11_lut (.I0(GND_net), .I1(n13597[8]), .I2(GND_net), 
            .I3(n37304), .O(n13112[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_11 (.CI(n37304), .I0(n13597[8]), .I1(GND_net), .CO(n37305));
    SB_LUT4 mult_14_add_1212_22_lut (.I0(GND_net), .I1(n1798[19]), .I2(GND_net), 
            .I3(n38702), .O(n1797[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_9_lut (.I0(GND_net), .I1(n8256[6]), .I2(GND_net), 
            .I3(n38371), .O(n8234[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_9 (.CI(n38371), .I0(n8256[6]), .I1(GND_net), .CO(n38372));
    SB_CARRY mult_14_add_1212_22 (.CI(n38702), .I0(n1798[19]), .I1(GND_net), 
            .CO(n38703));
    SB_LUT4 add_3094_8_lut (.I0(GND_net), .I1(n8256[5]), .I2(n713), .I3(n38370), 
            .O(n8234[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_4 (.CI(n37492), .I0(n14171[1]), .I1(n253), .CO(n37493));
    SB_LUT4 add_3300_10_lut (.I0(GND_net), .I1(n13597[7]), .I2(GND_net), 
            .I3(n37303), .O(n13112[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_10 (.CI(n37303), .I0(n13597[7]), .I1(GND_net), .CO(n37304));
    SB_CARRY add_3094_8 (.CI(n38370), .I0(n8256[5]), .I1(n713), .CO(n38371));
    SB_LUT4 add_3329_3_lut (.I0(GND_net), .I1(n14171[0]), .I2(n180), .I3(n37491), 
            .O(n13737[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3300_9_lut (.I0(GND_net), .I1(n13597[6]), .I2(GND_net), 
            .I3(n37302), .O(n13112[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3094_7_lut (.I0(GND_net), .I1(n8256[4]), .I2(n616), .I3(n38369), 
            .O(n8234[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_21_lut (.I0(GND_net), .I1(n1798[18]), .I2(GND_net), 
            .I3(n38701), .O(n1797[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_7 (.CI(n38369), .I0(n8256[4]), .I1(n616), .CO(n38370));
    SB_LUT4 add_3094_6_lut (.I0(GND_net), .I1(n8256[3]), .I2(n519_adj_3699), 
            .I3(n38368), .O(n8234[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_21 (.CI(n38701), .I0(n1798[18]), .I1(GND_net), 
            .CO(n38702));
    SB_CARRY add_3094_6 (.CI(n38368), .I0(n8256[3]), .I1(n519_adj_3699), 
            .CO(n38369));
    SB_CARRY add_3300_9 (.CI(n37302), .I0(n13597[6]), .I1(GND_net), .CO(n37303));
    SB_LUT4 add_3094_5_lut (.I0(GND_net), .I1(n8256[2]), .I2(n422), .I3(n38367), 
            .O(n8234[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_20_lut (.I0(GND_net), .I1(n1798[17]), .I2(GND_net), 
            .I3(n38700), .O(n1797[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_5 (.CI(n38367), .I0(n8256[2]), .I1(n422), .CO(n38368));
    SB_LUT4 add_3094_4_lut (.I0(GND_net), .I1(n8256[1]), .I2(n325), .I3(n38366), 
            .O(n8234[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_3 (.CI(n37491), .I0(n14171[0]), .I1(n180), .CO(n37492));
    SB_LUT4 add_3300_8_lut (.I0(GND_net), .I1(n13597[5]), .I2(n707), .I3(n37301), 
            .O(n13112[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_4 (.CI(n38366), .I0(n8256[1]), .I1(n325), .CO(n38367));
    SB_LUT4 add_3094_3_lut (.I0(GND_net), .I1(n8256[0]), .I2(n228_adj_3700), 
            .I3(n38365), .O(n8234[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3329_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n13737[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3329_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_8 (.CI(n37301), .I0(n13597[5]), .I1(n707), .CO(n37302));
    SB_CARRY mult_14_add_1212_20 (.CI(n38700), .I0(n1798[17]), .I1(GND_net), 
            .CO(n38701));
    SB_CARRY add_3094_3 (.CI(n38365), .I0(n8256[0]), .I1(n228_adj_3700), 
            .CO(n38366));
    SB_LUT4 add_3094_2_lut (.I0(GND_net), .I1(n38_adj_3701), .I2(n131_adj_3702), 
            .I3(GND_net), .O(n8234[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3094_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_19_lut (.I0(GND_net), .I1(n1798[16]), .I2(GND_net), 
            .I3(n38699), .O(n1797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3094_2 (.CI(GND_net), .I0(n38_adj_3701), .I1(n131_adj_3702), 
            .CO(n38365));
    SB_LUT4 add_3093_22_lut (.I0(GND_net), .I1(n8234[19]), .I2(GND_net), 
            .I3(n38364), .O(n8211[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_19 (.CI(n38699), .I0(n1798[16]), .I1(GND_net), 
            .CO(n38700));
    SB_LUT4 add_3093_21_lut (.I0(GND_net), .I1(n8234[18]), .I2(GND_net), 
            .I3(n38363), .O(n8211[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_18_lut (.I0(GND_net), .I1(n1798[15]), .I2(GND_net), 
            .I3(n38698), .O(n1797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_21 (.CI(n38363), .I0(n8234[18]), .I1(GND_net), .CO(n38364));
    SB_LUT4 add_3093_20_lut (.I0(GND_net), .I1(n8234[17]), .I2(GND_net), 
            .I3(n38362), .O(n8211[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3300_7_lut (.I0(GND_net), .I1(n13597[4]), .I2(n610_adj_3703), 
            .I3(n37300), .O(n13112[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_18 (.CI(n38698), .I0(n1798[15]), .I1(GND_net), 
            .CO(n38699));
    SB_CARRY add_3093_20 (.CI(n38362), .I0(n8234[17]), .I1(GND_net), .CO(n38363));
    SB_CARRY add_3300_7 (.CI(n37300), .I0(n13597[4]), .I1(n610_adj_3703), 
            .CO(n37301));
    SB_LUT4 add_3300_6_lut (.I0(GND_net), .I1(n13597[3]), .I2(n513), .I3(n37299), 
            .O(n13112[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_17_lut (.I0(GND_net), .I1(n1798[14]), .I2(GND_net), 
            .I3(n38697), .O(n1797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_19_lut (.I0(GND_net), .I1(n8234[16]), .I2(GND_net), 
            .I3(n38361), .O(n8211[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_17 (.CI(n38697), .I0(n1798[14]), .I1(GND_net), 
            .CO(n38698));
    SB_CARRY add_3093_19 (.CI(n38361), .I0(n8234[16]), .I1(GND_net), .CO(n38362));
    SB_CARRY add_3300_6 (.CI(n37299), .I0(n13597[3]), .I1(n513), .CO(n37300));
    SB_LUT4 add_3300_5_lut (.I0(GND_net), .I1(n13597[2]), .I2(n416_adj_3704), 
            .I3(n37298), .O(n13112[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_5 (.CI(n37298), .I0(n13597[2]), .I1(n416_adj_3704), 
            .CO(n37299));
    SB_LUT4 add_3093_18_lut (.I0(GND_net), .I1(n8234[15]), .I2(GND_net), 
            .I3(n38360), .O(n8211[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3300_4_lut (.I0(GND_net), .I1(n13597[1]), .I2(n319), .I3(n37297), 
            .O(n13112[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_4 (.CI(n37297), .I0(n13597[1]), .I1(n319), .CO(n37298));
    SB_LUT4 sub_11_add_2_27_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n76[26]), .I3(n37097), .O(n61[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_26_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[31] ), 
            .I2(n76[26]), .I3(n37096), .O(n61[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_16_lut (.I0(GND_net), .I1(n1798[13]), .I2(GND_net), 
            .I3(n38696), .O(n1797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_18 (.CI(n38360), .I0(n8234[15]), .I1(GND_net), .CO(n38361));
    SB_LUT4 add_3300_3_lut (.I0(GND_net), .I1(n13597[0]), .I2(n222_adj_3706), 
            .I3(n37296), .O(n13112[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_26 (.CI(n37096), .I0(\PID_CONTROLLER.err_prev[31] ), 
            .I1(n76[26]), .CO(n37097));
    SB_LUT4 sub_11_add_2_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[23] ), 
            .I2(n76[23]), .I3(n37095), .O(n61[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_3 (.CI(n37296), .I0(n13597[0]), .I1(n222_adj_3706), 
            .CO(n37297));
    SB_CARRY sub_11_add_2_25 (.CI(n37095), .I0(\PID_CONTROLLER.err_prev[23] ), 
            .I1(n76[23]), .CO(n37096));
    SB_LUT4 sub_11_add_2_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[22] ), 
            .I2(n76[22]), .I3(n37094), .O(n61[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_16 (.CI(n38696), .I0(n1798[13]), .I1(GND_net), 
            .CO(n38697));
    SB_LUT4 add_3300_2_lut (.I0(GND_net), .I1(n32_adj_3711), .I2(n125), 
            .I3(GND_net), .O(n13112[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3300_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_15_lut (.I0(GND_net), .I1(n1798[12]), .I2(GND_net), 
            .I3(n38695), .O(n1797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_17_lut (.I0(GND_net), .I1(n8234[14]), .I2(GND_net), 
            .I3(n38359), .O(n8211[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3300_2 (.CI(GND_net), .I0(n32_adj_3711), .I1(n125), .CO(n37296));
    SB_CARRY add_3093_17 (.CI(n38359), .I0(n8234[14]), .I1(GND_net), .CO(n38360));
    SB_LUT4 add_3322_22_lut (.I0(GND_net), .I1(n14038[19]), .I2(GND_net), 
            .I3(n37295), .O(n13597[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_24 (.CI(n37094), .I0(\PID_CONTROLLER.err_prev[22] ), 
            .I1(n76[22]), .CO(n37095));
    SB_LUT4 sub_11_add_2_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[21] ), 
            .I2(n76[21]), .I3(n37093), .O(n61[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_21_lut (.I0(GND_net), .I1(n14038[18]), .I2(GND_net), 
            .I3(n37294), .O(n13597[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_23 (.CI(n37093), .I0(\PID_CONTROLLER.err_prev[21] ), 
            .I1(n76[21]), .CO(n37094));
    SB_LUT4 sub_11_add_2_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[20] ), 
            .I2(n76[20]), .I3(n37092), .O(n61[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_15 (.CI(n38695), .I0(n1798[12]), .I1(GND_net), 
            .CO(n38696));
    SB_LUT4 add_3093_16_lut (.I0(GND_net), .I1(n8234[13]), .I2(GND_net), 
            .I3(n38358), .O(n8211[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_21 (.CI(n37294), .I0(n14038[18]), .I1(GND_net), 
            .CO(n37295));
    SB_CARRY sub_11_add_2_22 (.CI(n37092), .I0(\PID_CONTROLLER.err_prev[20] ), 
            .I1(n76[20]), .CO(n37093));
    SB_LUT4 sub_11_add_2_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[19] ), 
            .I2(n76[19]), .I3(n37091), .O(n61[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_20_lut (.I0(GND_net), .I1(n14038[17]), .I2(GND_net), 
            .I3(n37293), .O(n13597[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_21 (.CI(n37091), .I0(\PID_CONTROLLER.err_prev[19] ), 
            .I1(n76[19]), .CO(n37092));
    SB_LUT4 sub_11_add_2_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[18] ), 
            .I2(n76[18]), .I3(n37090), .O(n61[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_16 (.CI(n38358), .I0(n8234[13]), .I1(GND_net), .CO(n38359));
    SB_LUT4 add_3093_15_lut (.I0(GND_net), .I1(n8234[12]), .I2(GND_net), 
            .I3(n38357), .O(n8211[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3329_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n37491));
    SB_CARRY add_3322_20 (.CI(n37293), .I0(n14038[17]), .I1(GND_net), 
            .CO(n37294));
    SB_CARRY sub_11_add_2_20 (.CI(n37090), .I0(\PID_CONTROLLER.err_prev[18] ), 
            .I1(n76[18]), .CO(n37091));
    SB_LUT4 sub_11_add_2_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[17] ), 
            .I2(n76[17]), .I3(n37089), .O(n61[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_15 (.CI(n38357), .I0(n8234[12]), .I1(GND_net), .CO(n38358));
    SB_LUT4 add_3170_28_lut (.I0(GND_net), .I1(n10674[25]), .I2(GND_net), 
            .I3(n37490), .O(n9932[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_19_lut (.I0(GND_net), .I1(n14038[16]), .I2(GND_net), 
            .I3(n37292), .O(n13597[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_19 (.CI(n37089), .I0(\PID_CONTROLLER.err_prev[17] ), 
            .I1(n76[17]), .CO(n37090));
    SB_LUT4 sub_11_add_2_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[16] ), 
            .I2(n76[16]), .I3(n37088), .O(n61[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_14_lut (.I0(GND_net), .I1(n1798[11]), .I2(GND_net), 
            .I3(n38694), .O(n1797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_14_lut (.I0(GND_net), .I1(n8234[11]), .I2(GND_net), 
            .I3(n38356), .O(n8211[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_14 (.CI(n38356), .I0(n8234[11]), .I1(GND_net), .CO(n38357));
    SB_CARRY mult_14_add_1212_14 (.CI(n38694), .I0(n1798[11]), .I1(GND_net), 
            .CO(n38695));
    SB_LUT4 add_3093_13_lut (.I0(GND_net), .I1(n8234[10]), .I2(GND_net), 
            .I3(n38355), .O(n8211[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_27_lut (.I0(GND_net), .I1(n10674[24]), .I2(GND_net), 
            .I3(n37489), .O(n9932[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_19 (.CI(n37292), .I0(n14038[16]), .I1(GND_net), 
            .CO(n37293));
    SB_LUT4 add_3322_18_lut (.I0(GND_net), .I1(n14038[15]), .I2(GND_net), 
            .I3(n37291), .O(n13597[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_18 (.CI(n37088), .I0(\PID_CONTROLLER.err_prev[16] ), 
            .I1(n76[16]), .CO(n37089));
    SB_LUT4 sub_11_add_2_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[15] ), 
            .I2(n76[15]), .I3(n37087), .O(n61[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_17 (.CI(n37087), .I0(\PID_CONTROLLER.err_prev[15] ), 
            .I1(n76[15]), .CO(n37088));
    SB_LUT4 sub_11_add_2_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[14] ), 
            .I2(n76[14]), .I3(n37086), .O(n61[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_18 (.CI(n37291), .I0(n14038[15]), .I1(GND_net), 
            .CO(n37292));
    SB_CARRY sub_11_add_2_16 (.CI(n37086), .I0(\PID_CONTROLLER.err_prev[14] ), 
            .I1(n76[14]), .CO(n37087));
    SB_CARRY add_3093_13 (.CI(n38355), .I0(n8234[10]), .I1(GND_net), .CO(n38356));
    SB_LUT4 sub_11_add_2_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[13] ), 
            .I2(n76[13]), .I3(n37085), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_12_lut (.I0(GND_net), .I1(n8234[9]), .I2(GND_net), 
            .I3(n38354), .O(n8211[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_27 (.CI(n37489), .I0(n10674[24]), .I1(GND_net), 
            .CO(n37490));
    SB_LUT4 add_3322_17_lut (.I0(GND_net), .I1(n14038[14]), .I2(GND_net), 
            .I3(n37290), .O(n13597[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_12 (.CI(n38354), .I0(n8234[9]), .I1(GND_net), .CO(n38355));
    SB_LUT4 mult_14_add_1212_13_lut (.I0(GND_net), .I1(n1798[10]), .I2(GND_net), 
            .I3(n38693), .O(n1797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_15 (.CI(n37085), .I0(\PID_CONTROLLER.err_prev[13] ), 
            .I1(n76[13]), .CO(n37086));
    SB_LUT4 add_3093_11_lut (.I0(GND_net), .I1(n8234[8]), .I2(GND_net), 
            .I3(n38353), .O(n8211[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_13 (.CI(n38693), .I0(n1798[10]), .I1(GND_net), 
            .CO(n38694));
    SB_LUT4 sub_11_add_2_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[12] ), 
            .I2(n76[12]), .I3(n37084), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_11 (.CI(n38353), .I0(n8234[8]), .I1(GND_net), .CO(n38354));
    SB_LUT4 add_3093_10_lut (.I0(GND_net), .I1(n8234[7]), .I2(GND_net), 
            .I3(n38352), .O(n8211[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_12_lut (.I0(GND_net), .I1(n1798[9]), .I2(GND_net), 
            .I3(n38692), .O(n1797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_10 (.CI(n38352), .I0(n8234[7]), .I1(GND_net), .CO(n38353));
    SB_LUT4 add_3093_9_lut (.I0(GND_net), .I1(n8234[6]), .I2(GND_net), 
            .I3(n38351), .O(n8211[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_9 (.CI(n38351), .I0(n8234[6]), .I1(GND_net), .CO(n38352));
    SB_LUT4 add_3093_8_lut (.I0(GND_net), .I1(n8234[5]), .I2(n710), .I3(n38350), 
            .O(n8211[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_12 (.CI(n38692), .I0(n1798[9]), .I1(GND_net), 
            .CO(n38693));
    SB_CARRY add_3093_8 (.CI(n38350), .I0(n8234[5]), .I1(n710), .CO(n38351));
    SB_LUT4 mult_14_add_1212_11_lut (.I0(GND_net), .I1(n1798[8]), .I2(GND_net), 
            .I3(n38691), .O(n1797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_10_lut (.I0(GND_net), .I1(n1804[22]), .I2(n1711), 
            .I3(n38893), .O(n7068[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_26_lut (.I0(GND_net), .I1(n10674[23]), .I2(GND_net), 
            .I3(n37488), .O(n9932[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_17 (.CI(n37290), .I0(n14038[14]), .I1(GND_net), 
            .CO(n37291));
    SB_CARRY sub_11_add_2_14 (.CI(n37084), .I0(\PID_CONTROLLER.err_prev[12] ), 
            .I1(n76[12]), .CO(n37085));
    SB_LUT4 add_3093_7_lut (.I0(GND_net), .I1(n8234[4]), .I2(n613), .I3(n38349), 
            .O(n8211[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_9_lut (.I0(GND_net), .I1(n1803[22]), .I2(n1707), 
            .I3(n38892), .O(n7068[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_7 (.CI(n38349), .I0(n8234[4]), .I1(n613), .CO(n38350));
    SB_LUT4 add_3322_16_lut (.I0(GND_net), .I1(n14038[13]), .I2(GND_net), 
            .I3(n37289), .O(n13597[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_6_lut (.I0(GND_net), .I1(n8234[3]), .I2(n516), .I3(n38348), 
            .O(n8211[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3052_9 (.CI(n38892), .I0(n1803[22]), .I1(n1707), .CO(n38893));
    SB_CARRY add_3322_16 (.CI(n37289), .I0(n14038[13]), .I1(GND_net), 
            .CO(n37290));
    SB_LUT4 add_3052_8_lut (.I0(GND_net), .I1(n1802[22]), .I2(n1703), 
            .I3(n38891), .O(n7068[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[11] ), 
            .I2(n76[11]), .I3(n37083), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_13 (.CI(n37083), .I0(\PID_CONTROLLER.err_prev[11] ), 
            .I1(n76[11]), .CO(n37084));
    SB_CARRY mult_14_add_1212_11 (.CI(n38691), .I0(n1798[8]), .I1(GND_net), 
            .CO(n38692));
    SB_LUT4 add_3322_15_lut (.I0(GND_net), .I1(n14038[12]), .I2(GND_net), 
            .I3(n37288), .O(n13597[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_6 (.CI(n38348), .I0(n8234[3]), .I1(n516), .CO(n38349));
    SB_CARRY add_3052_8 (.CI(n38891), .I0(n1802[22]), .I1(n1703), .CO(n38892));
    SB_LUT4 mult_14_add_1212_10_lut (.I0(GND_net), .I1(n1798[7]), .I2(GND_net), 
            .I3(n38690), .O(n1797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_15 (.CI(n37288), .I0(n14038[12]), .I1(GND_net), 
            .CO(n37289));
    SB_LUT4 sub_11_add_2_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[10] ), 
            .I2(n76[10]), .I3(n37082), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_10 (.CI(n38690), .I0(n1798[7]), .I1(GND_net), 
            .CO(n38691));
    SB_CARRY sub_11_add_2_12 (.CI(n37082), .I0(\PID_CONTROLLER.err_prev[10] ), 
            .I1(n76[10]), .CO(n37083));
    SB_LUT4 add_3322_14_lut (.I0(GND_net), .I1(n14038[11]), .I2(GND_net), 
            .I3(n37287), .O(n13597[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[9] ), 
            .I2(n76[9]), .I3(n37081), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_11 (.CI(n37081), .I0(\PID_CONTROLLER.err_prev[9] ), 
            .I1(n76[9]), .CO(n37082));
    SB_CARRY add_3322_14 (.CI(n37287), .I0(n14038[11]), .I1(GND_net), 
            .CO(n37288));
    SB_LUT4 add_3322_13_lut (.I0(GND_net), .I1(n14038[10]), .I2(GND_net), 
            .I3(n37286), .O(n13597[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_26 (.CI(n37488), .I0(n10674[23]), .I1(GND_net), 
            .CO(n37489));
    SB_LUT4 add_3170_25_lut (.I0(GND_net), .I1(n10674[22]), .I2(GND_net), 
            .I3(n37487), .O(n9932[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_13 (.CI(n37286), .I0(n14038[10]), .I1(GND_net), 
            .CO(n37287));
    SB_LUT4 add_3322_12_lut (.I0(GND_net), .I1(n14038[9]), .I2(GND_net), 
            .I3(n37285), .O(n13597[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_12 (.CI(n37285), .I0(n14038[9]), .I1(GND_net), .CO(n37286));
    SB_LUT4 mult_14_add_1212_9_lut (.I0(GND_net), .I1(n1798[6]), .I2(GND_net), 
            .I3(n38689), .O(n1797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[8] ), 
            .I2(n76[8]), .I3(n37080), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_5_lut (.I0(GND_net), .I1(n8234[2]), .I2(n419_adj_3731), 
            .I3(n38347), .O(n8211[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_9 (.CI(n38689), .I0(n1798[6]), .I1(GND_net), 
            .CO(n38690));
    SB_LUT4 add_3322_11_lut (.I0(GND_net), .I1(n14038[8]), .I2(GND_net), 
            .I3(n37284), .O(n13597[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_10 (.CI(n37080), .I0(\PID_CONTROLLER.err_prev[8] ), 
            .I1(n76[8]), .CO(n37081));
    SB_LUT4 sub_11_add_2_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[7] ), 
            .I2(n76[7]), .I3(n37079), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_9 (.CI(n37079), .I0(\PID_CONTROLLER.err_prev[7] ), 
            .I1(n76[7]), .CO(n37080));
    SB_CARRY add_3093_5 (.CI(n38347), .I0(n8234[2]), .I1(n419_adj_3731), 
            .CO(n38348));
    SB_LUT4 add_3093_4_lut (.I0(GND_net), .I1(n8234[1]), .I2(n322), .I3(n38346), 
            .O(n8211[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_25 (.CI(n37487), .I0(n10674[22]), .I1(GND_net), 
            .CO(n37488));
    SB_CARRY add_3093_4 (.CI(n38346), .I0(n8234[1]), .I1(n322), .CO(n38347));
    SB_CARRY add_3322_11 (.CI(n37284), .I0(n14038[8]), .I1(GND_net), .CO(n37285));
    SB_LUT4 add_3093_3_lut (.I0(GND_net), .I1(n8234[0]), .I2(n225_adj_3733), 
            .I3(n38345), .O(n8211[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[6] ), 
            .I2(n76[6]), .I3(n37078), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_10_lut (.I0(GND_net), .I1(n14038[7]), .I2(GND_net), 
            .I3(n37283), .O(n13597[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_8 (.CI(n37078), .I0(\PID_CONTROLLER.err_prev[6] ), 
            .I1(n76[6]), .CO(n37079));
    SB_LUT4 sub_11_add_2_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[5] ), 
            .I2(n76[5]), .I3(n37077), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_17_inv_0_i32_1_lut (.I0(\deadband[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n64[31]));   // verilog/motorControl.v(37[41:50])
    defparam unary_minus_17_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_11_add_2_7 (.CI(n37077), .I0(\PID_CONTROLLER.err_prev[5] ), 
            .I1(n76[5]), .CO(n37078));
    SB_LUT4 sub_11_add_2_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[4] ), 
            .I2(n76[4]), .I3(n37076), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i105_2_lut (.I0(\Kd[1] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n155_adj_3530));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i105_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_11_add_2_6 (.CI(n37076), .I0(\PID_CONTROLLER.err_prev[4] ), 
            .I1(n76[4]), .CO(n37077));
    SB_LUT4 mult_12_i42_2_lut (.I0(\Kd[0] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_3529));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3322_10 (.CI(n37283), .I0(n14038[7]), .I1(GND_net), .CO(n37284));
    SB_LUT4 sub_11_add_2_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[3] ), 
            .I2(n76[3]), .I3(n37075), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_5 (.CI(n37075), .I0(\PID_CONTROLLER.err_prev[3] ), 
            .I1(n76[3]), .CO(n37076));
    SB_LUT4 add_3052_7_lut (.I0(GND_net), .I1(n1801[22]), .I2(n1699), 
            .I3(n38890), .O(n7068[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_8_lut (.I0(GND_net), .I1(n1798[5]), .I2(n515), 
            .I3(n38688), .O(n1797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3093_3 (.CI(n38345), .I0(n8234[0]), .I1(n225_adj_3733), 
            .CO(n38346));
    SB_LUT4 add_3322_9_lut (.I0(GND_net), .I1(n14038[6]), .I2(GND_net), 
            .I3(n37282), .O(n13597[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_11_add_2_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[2] ), 
            .I2(n76[2]), .I3(n37074), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_9 (.CI(n37282), .I0(n14038[6]), .I1(GND_net), .CO(n37283));
    SB_CARRY sub_11_add_2_4 (.CI(n37074), .I0(\PID_CONTROLLER.err_prev[2] ), 
            .I1(n76[2]), .CO(n37075));
    SB_LUT4 sub_11_add_2_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[1] ), 
            .I2(n76[1]), .I3(n37073), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3093_2_lut (.I0(GND_net), .I1(n35_adj_3741), .I2(n128_adj_3742), 
            .I3(GND_net), .O(n8211[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3093_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3322_8_lut (.I0(GND_net), .I1(n14038[5]), .I2(n710_adj_3743), 
            .I3(n37281), .O(n13597[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_3 (.CI(n37073), .I0(\PID_CONTROLLER.err_prev[1] ), 
            .I1(n76[1]), .CO(n37074));
    SB_CARRY add_3322_8 (.CI(n37281), .I0(n14038[5]), .I1(n710_adj_3743), 
            .CO(n37282));
    SB_LUT4 sub_11_add_2_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.err_prev[0] ), 
            .I2(n76[0]), .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_11_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_8 (.CI(n38688), .I0(n1798[5]), .I1(n515), 
            .CO(n38689));
    SB_CARRY add_3093_2 (.CI(GND_net), .I0(n35_adj_3741), .I1(n128_adj_3742), 
            .CO(n38345));
    SB_LUT4 add_3322_7_lut (.I0(GND_net), .I1(n14038[4]), .I2(n613_adj_3745), 
            .I3(n37280), .O(n13597[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_11_add_2_2 (.CI(VCC_net), .I0(\PID_CONTROLLER.err_prev[0] ), 
            .I1(n76[0]), .CO(n37073));
    SB_LUT4 unary_minus_70_add_3_25_lut (.I0(n852[14]), .I1(GND_net), .I2(PHASES_5__N_3046), 
            .I3(n37072), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3322_7 (.CI(n37280), .I0(n14038[4]), .I1(n613_adj_3745), 
            .CO(n37281));
    SB_LUT4 unary_minus_70_add_3_24_lut (.I0(n852[18]), .I1(GND_net), .I2(n79[22]), 
            .I3(n37071), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_24_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_3322_6_lut (.I0(GND_net), .I1(n14038[3]), .I2(n516_adj_3749), 
            .I3(n37279), .O(n13597[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_6 (.CI(n37279), .I0(n14038[3]), .I1(n516_adj_3749), 
            .CO(n37280));
    SB_LUT4 add_3322_5_lut (.I0(GND_net), .I1(n14038[2]), .I2(n419_adj_3750), 
            .I3(n37278), .O(n13597[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_23_lut (.I0(GND_net), .I1(n8211[20]), .I2(GND_net), 
            .I3(n38344), .O(n8187[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_24 (.CI(n37071), .I0(GND_net), .I1(n79[22]), 
            .CO(n37072));
    SB_CARRY add_3052_7 (.CI(n38890), .I0(n1801[22]), .I1(n1699), .CO(n38891));
    SB_DFF \PID_CONTROLLER.err_prev__i2  (.Q(\PID_CONTROLLER.err_prev[1] ), 
           .C(clk32MHz), .D(n23900));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 mult_14_add_1212_7_lut (.I0(GND_net), .I1(n1798[4]), .I2(n442), 
            .I3(n38687), .O(n1797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i3  (.Q(\PID_CONTROLLER.err_prev[2] ), 
           .C(clk32MHz), .D(n23899));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3322_5 (.CI(n37278), .I0(n14038[2]), .I1(n419_adj_3750), 
            .CO(n37279));
    SB_DFF \PID_CONTROLLER.err_prev__i4  (.Q(\PID_CONTROLLER.err_prev[3] ), 
           .C(clk32MHz), .D(n23898));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3322_4_lut (.I0(GND_net), .I1(n14038[1]), .I2(n322_adj_3752), 
            .I3(n37277), .O(n13597[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i5  (.Q(\PID_CONTROLLER.err_prev[4] ), 
           .C(clk32MHz), .D(n23897));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i6  (.Q(\PID_CONTROLLER.err_prev[5] ), 
           .C(clk32MHz), .D(n23896));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3052_6_lut (.I0(GND_net), .I1(n1800[22]), .I2(n1695), 
            .I3(n38889), .O(n7068[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i7  (.Q(\PID_CONTROLLER.err_prev[6] ), 
           .C(clk32MHz), .D(n23895));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3092_22_lut (.I0(GND_net), .I1(n8211[19]), .I2(GND_net), 
            .I3(n38343), .O(n8187[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_22_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i8  (.Q(\PID_CONTROLLER.err_prev[7] ), 
           .C(clk32MHz), .D(n23894));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY mult_14_add_1212_7 (.CI(n38687), .I0(n1798[4]), .I1(n442), 
            .CO(n38688));
    SB_DFF \PID_CONTROLLER.err_prev__i9  (.Q(\PID_CONTROLLER.err_prev[8] ), 
           .C(clk32MHz), .D(n23893));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i10  (.Q(\PID_CONTROLLER.err_prev[9] ), 
           .C(clk32MHz), .D(n23892));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3092_22 (.CI(n38343), .I0(n8211[19]), .I1(GND_net), .CO(n38344));
    SB_DFF \PID_CONTROLLER.err_prev__i11  (.Q(\PID_CONTROLLER.err_prev[10] ), 
           .C(clk32MHz), .D(n23891));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i12  (.Q(\PID_CONTROLLER.err_prev[11] ), 
           .C(clk32MHz), .D(n23890));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i13  (.Q(\PID_CONTROLLER.err_prev[12] ), 
           .C(clk32MHz), .D(n23889));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 unary_minus_70_add_3_23_lut (.I0(n852[10]), .I1(GND_net), .I2(n79[21]), 
            .I3(n37070), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_23_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_3092_21_lut (.I0(GND_net), .I1(n8211[18]), .I2(GND_net), 
            .I3(n38342), .O(n8187[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i14  (.Q(\PID_CONTROLLER.err_prev[13] ), 
           .C(clk32MHz), .D(n23888));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3322_4 (.CI(n37277), .I0(n14038[1]), .I1(n322_adj_3752), 
            .CO(n37278));
    SB_DFF \PID_CONTROLLER.err_prev__i15  (.Q(\PID_CONTROLLER.err_prev[14] ), 
           .C(clk32MHz), .D(n23887));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3322_3_lut (.I0(GND_net), .I1(n14038[0]), .I2(n225_adj_3755), 
            .I3(n37276), .O(n13597[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3322_3 (.CI(n37276), .I0(n14038[0]), .I1(n225_adj_3755), 
            .CO(n37277));
    SB_DFF \PID_CONTROLLER.err_prev__i16  (.Q(\PID_CONTROLLER.err_prev[15] ), 
           .C(clk32MHz), .D(n23886));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i17  (.Q(\PID_CONTROLLER.err_prev[16] ), 
           .C(clk32MHz), .D(n23885));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i18  (.Q(\PID_CONTROLLER.err_prev[17] ), 
           .C(clk32MHz), .D(n23884));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 add_3322_2_lut (.I0(GND_net), .I1(n35_adj_3756), .I2(n128_adj_3757), 
            .I3(GND_net), .O(n13597[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3322_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i19  (.Q(\PID_CONTROLLER.err_prev[18] ), 
           .C(clk32MHz), .D(n23883));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY unary_minus_70_add_3_23 (.CI(n37070), .I0(GND_net), .I1(n79[21]), 
            .CO(n37071));
    SB_CARRY add_3052_6 (.CI(n38889), .I0(n1800[22]), .I1(n1695), .CO(n38890));
    SB_DFF \PID_CONTROLLER.err_prev__i20  (.Q(\PID_CONTROLLER.err_prev[19] ), 
           .C(clk32MHz), .D(n23882));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i21  (.Q(\PID_CONTROLLER.err_prev[20] ), 
           .C(clk32MHz), .D(n23881));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 mult_14_add_1212_6_lut (.I0(GND_net), .I1(n1798[3]), .I2(n369), 
            .I3(n38686), .O(n1797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_prev__i22  (.Q(\PID_CONTROLLER.err_prev[21] ), 
           .C(clk32MHz), .D(n23880));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_prev__i23  (.Q(\PID_CONTROLLER.err_prev[22] ), 
           .C(clk32MHz), .D(n23879));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY mult_14_add_1212_6 (.CI(n38686), .I0(n1798[3]), .I1(n369), 
            .CO(n38687));
    SB_DFF \PID_CONTROLLER.err_prev__i24  (.Q(\PID_CONTROLLER.err_prev[23] ), 
           .C(clk32MHz), .D(n23878));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 unary_minus_70_add_3_22_lut (.I0(n852[16]), .I1(GND_net), .I2(n79[20]), 
            .I3(n37069), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3322_2 (.CI(GND_net), .I0(n35_adj_3756), .I1(n128_adj_3757), 
            .CO(n37276));
    SB_CARRY add_3092_21 (.CI(n38342), .I0(n8211[18]), .I1(GND_net), .CO(n38343));
    SB_CARRY unary_minus_70_add_3_22 (.CI(n37069), .I0(GND_net), .I1(n79[20]), 
            .CO(n37070));
    SB_DFF \PID_CONTROLLER.err_prev__i25  (.Q(\PID_CONTROLLER.err_prev[31] ), 
           .C(clk32MHz), .D(n23877));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 unary_minus_70_add_3_21_lut (.I0(n852[11]), .I1(GND_net), .I2(n79[19]), 
            .I3(n37068), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_21_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mult_14_add_1212_5_lut (.I0(GND_net), .I1(n1798[2]), .I2(n296_adj_3764), 
            .I3(n38685), .O(n1797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_20_lut (.I0(GND_net), .I1(n8211[17]), .I2(GND_net), 
            .I3(n38341), .O(n8187[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_21 (.CI(n37068), .I0(GND_net), .I1(n79[19]), 
            .CO(n37069));
    SB_CARRY add_3092_20 (.CI(n38341), .I0(n8211[17]), .I1(GND_net), .CO(n38342));
    SB_LUT4 add_3052_5_lut (.I0(GND_net), .I1(n1799[22]), .I2(n1691), 
            .I3(n38888), .O(n7068[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1212_5 (.CI(n38685), .I0(n1798[2]), .I1(n296_adj_3764), 
            .CO(n38686));
    SB_LUT4 add_3492_11_lut (.I0(GND_net), .I1(n16508[8]), .I2(GND_net), 
            .I3(n37275), .O(n16423[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n79[18]), 
            .I3(n37067), .O(n852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_10_lut (.I0(GND_net), .I1(n16508[7]), .I2(GND_net), 
            .I3(n37274), .O(n16423[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_19_lut (.I0(GND_net), .I1(n8211[16]), .I2(GND_net), 
            .I3(n38340), .O(n8187[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_10 (.CI(n37274), .I0(n16508[7]), .I1(GND_net), .CO(n37275));
    SB_CARRY unary_minus_70_add_3_20 (.CI(n37067), .I0(GND_net), .I1(n79[18]), 
            .CO(n37068));
    SB_CARRY add_3092_19 (.CI(n38340), .I0(n8211[16]), .I1(GND_net), .CO(n38341));
    SB_LUT4 add_3492_9_lut (.I0(GND_net), .I1(n16508[6]), .I2(GND_net), 
            .I3(n37273), .O(n16423[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_19_lut (.I0(n852[15]), .I1(GND_net), .I2(n79[17]), 
            .I3(n37066), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_19_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_3092_18_lut (.I0(GND_net), .I1(n8211[15]), .I2(GND_net), 
            .I3(n38339), .O(n8187[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_19 (.CI(n37066), .I0(GND_net), .I1(n79[17]), 
            .CO(n37067));
    SB_CARRY add_3492_9 (.CI(n37273), .I0(n16508[6]), .I1(GND_net), .CO(n37274));
    SB_LUT4 unary_minus_70_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n79[16]), 
            .I3(n37065), .O(n852[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3092_18 (.CI(n38339), .I0(n8211[15]), .I1(GND_net), .CO(n38340));
    SB_CARRY unary_minus_70_add_3_18 (.CI(n37065), .I0(GND_net), .I1(n79[16]), 
            .CO(n37066));
    SB_LUT4 add_3492_8_lut (.I0(GND_net), .I1(n16508[5]), .I2(n743_adj_3769), 
            .I3(n37272), .O(n16423[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n79[15]), 
            .I3(n37064), .O(n852[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_4_lut (.I0(GND_net), .I1(n1798[1]), .I2(n223_adj_3772), 
            .I3(n38684), .O(n1797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_17_lut (.I0(GND_net), .I1(n8211[14]), .I2(GND_net), 
            .I3(n38338), .O(n8187[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_17_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.result_i1  (.Q(\PID_CONTROLLER.result [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [1]));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3492_8 (.CI(n37272), .I0(n16508[5]), .I1(n743_adj_3769), 
            .CO(n37273));
    SB_CARRY unary_minus_70_add_3_17 (.CI(n37064), .I0(GND_net), .I1(n79[15]), 
            .CO(n37065));
    SB_LUT4 unary_minus_70_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n79[14]), 
            .I3(n37063), .O(n852[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_7_lut (.I0(GND_net), .I1(n16508[4]), .I2(n646_adj_3774), 
            .I3(n37271), .O(n16423[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_16 (.CI(n37063), .I0(GND_net), .I1(n79[14]), 
            .CO(n37064));
    SB_LUT4 mult_12_i170_2_lut (.I0(\Kd[2] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n252_adj_3527));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i170_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_add_3_15_lut (.I0(n48782), .I1(GND_net), .I2(n79[13]), 
            .I3(n37062), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_3092_17 (.CI(n38338), .I0(n8211[14]), .I1(GND_net), .CO(n38339));
    SB_CARRY add_3492_7 (.CI(n37271), .I0(n16508[4]), .I1(n646_adj_3774), 
            .CO(n37272));
    SB_CARRY mult_14_add_1212_4 (.CI(n38684), .I0(n1798[1]), .I1(n223_adj_3772), 
            .CO(n38685));
    SB_CARRY unary_minus_70_add_3_15 (.CI(n37062), .I0(GND_net), .I1(n79[13]), 
            .CO(n37063));
    SB_LUT4 add_3092_16_lut (.I0(GND_net), .I1(n8211[13]), .I2(GND_net), 
            .I3(n38337), .O(n8187[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_24_lut (.I0(GND_net), .I1(n10674[21]), .I2(GND_net), 
            .I3(n37486), .O(n9932[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_6_lut (.I0(GND_net), .I1(n16508[3]), .I2(n549_adj_3777), 
            .I3(n37270), .O(n16423[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_6 (.CI(n37270), .I0(n16508[3]), .I1(n549_adj_3777), 
            .CO(n37271));
    SB_LUT4 mult_14_add_1212_3_lut (.I0(GND_net), .I1(n1798[0]), .I2(n150_adj_3779), 
            .I3(n38683), .O(n1797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_14_lut (.I0(n852[9]), .I1(GND_net), .I2(n79[12]), 
            .I3(n37061), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_14_lut.LUT_INIT = 16'hebbe;
    SB_DFF \PID_CONTROLLER.result_i2  (.Q(\PID_CONTROLLER.result [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [2]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i3  (.Q(\PID_CONTROLLER.result [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [3]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i4  (.Q(\PID_CONTROLLER.result [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [4]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i5  (.Q(\PID_CONTROLLER.result[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [5]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i6  (.Q(\PID_CONTROLLER.result[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [6]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i7  (.Q(\PID_CONTROLLER.result[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [7]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i8  (.Q(\PID_CONTROLLER.result [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [8]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i9  (.Q(\PID_CONTROLLER.result [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [9]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i10  (.Q(\PID_CONTROLLER.result [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [10]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i11  (.Q(\PID_CONTROLLER.result [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [11]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i12  (.Q(\PID_CONTROLLER.result [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [12]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i13  (.Q(\PID_CONTROLLER.result [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [13]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i14  (.Q(\PID_CONTROLLER.result [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [14]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i15  (.Q(\PID_CONTROLLER.result [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [15]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i16  (.Q(\PID_CONTROLLER.result [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [16]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i17  (.Q(\PID_CONTROLLER.result [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [17]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i18  (.Q(\PID_CONTROLLER.result [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [18]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i19  (.Q(\PID_CONTROLLER.result [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [19]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i20  (.Q(\PID_CONTROLLER.result [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [20]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i21  (.Q(\PID_CONTROLLER.result [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [21]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i22  (.Q(\PID_CONTROLLER.result [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [22]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i23  (.Q(\PID_CONTROLLER.result [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [23]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i24  (.Q(\PID_CONTROLLER.result [24]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [24]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i25  (.Q(\PID_CONTROLLER.result [25]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [25]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i26  (.Q(\PID_CONTROLLER.result [26]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [26]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i27  (.Q(\PID_CONTROLLER.result [27]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [27]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i28  (.Q(\PID_CONTROLLER.result [28]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [28]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i29  (.Q(\PID_CONTROLLER.result [29]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [29]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i30  (.Q(\PID_CONTROLLER.result [30]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [30]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.result_i31  (.Q(\PID_CONTROLLER.result [31]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.result_31__N_2994 [31]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err[1] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [1]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFFE PHASES_i3 (.Q(PIN_8_c_2), .C(clk32MHz), .E(n10_adj_3782), 
            .D(PHASES_5__N_2779[2]));   // verilog/motorControl.v(57[10] 100[6])
    SB_DFFE PHASES_i4 (.Q(PIN_9_c_3), .C(clk32MHz), .E(n10_adj_3783), 
            .D(PHASES_5__N_2779[3]));   // verilog/motorControl.v(57[10] 100[6])
    SB_DFFE PHASES_i5 (.Q(PIN_10_c_4), .C(clk32MHz), .E(n43196), .D(PHASES_5__N_2779[4]));   // verilog/motorControl.v(57[10] 100[6])
    SB_DFFE PHASES_i6 (.Q(PIN_11_c_5), .C(clk32MHz), .E(n43194), .D(PHASES_5__N_2779[5]));   // verilog/motorControl.v(57[10] 100[6])
    SB_CARRY add_3092_16 (.CI(n38337), .I0(n8211[13]), .I1(GND_net), .CO(n38338));
    SB_CARRY add_3170_24 (.CI(n37486), .I0(n10674[21]), .I1(GND_net), 
            .CO(n37487));
    SB_LUT4 add_3492_5_lut (.I0(GND_net), .I1(n16508[2]), .I2(n452_adj_3784), 
            .I3(n37269), .O(n16423[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_14 (.CI(n37061), .I0(GND_net), .I1(n79[12]), 
            .CO(n37062));
    SB_LUT4 unary_minus_70_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n79[11]), 
            .I3(n37060), .O(n852[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3052_5 (.CI(n38888), .I0(n1799[22]), .I1(n1691), .CO(n38889));
    SB_CARRY add_3492_5 (.CI(n37269), .I0(n16508[2]), .I1(n452_adj_3784), 
            .CO(n37270));
    SB_CARRY mult_14_add_1212_3 (.CI(n38683), .I0(n1798[0]), .I1(n150_adj_3779), 
            .CO(n38684));
    SB_CARRY unary_minus_70_add_3_13 (.CI(n37060), .I0(GND_net), .I1(n79[11]), 
            .CO(n37061));
    SB_LUT4 add_3092_15_lut (.I0(GND_net), .I1(n8211[12]), .I2(GND_net), 
            .I3(n38336), .O(n8187[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3092_15 (.CI(n38336), .I0(n8211[12]), .I1(GND_net), .CO(n38337));
    SB_LUT4 unary_minus_70_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n79[10]), 
            .I3(n37059), .O(n852[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1212_2_lut (.I0(GND_net), .I1(n8_adj_3787), .I2(n77), 
            .I3(GND_net), .O(n1797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1212_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_14_lut (.I0(GND_net), .I1(n8211[11]), .I2(GND_net), 
            .I3(n38335), .O(n8187[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_4_lut (.I0(GND_net), .I1(n1798[22]), .I2(n1687), 
            .I3(n38887), .O(n7068[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_23_lut (.I0(GND_net), .I1(n10674[20]), .I2(GND_net), 
            .I3(n37485), .O(n9932[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3492_4_lut (.I0(GND_net), .I1(n16508[1]), .I2(n355_adj_3788), 
            .I3(n37268), .O(n16423[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_12 (.CI(n37059), .I0(GND_net), .I1(n79[10]), 
            .CO(n37060));
    SB_CARRY mult_14_add_1212_2 (.CI(GND_net), .I0(n8_adj_3787), .I1(n77), 
            .CO(n38683));
    SB_CARRY add_3092_14 (.CI(n38335), .I0(n8211[11]), .I1(GND_net), .CO(n38336));
    SB_LUT4 unary_minus_70_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n79[9]), 
            .I3(n37058), .O(n852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_13_lut (.I0(GND_net), .I1(n8211[10]), .I2(GND_net), 
            .I3(n38334), .O(n8187[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_23 (.CI(n37485), .I0(n10674[20]), .I1(GND_net), 
            .CO(n37486));
    SB_CARRY add_3492_4 (.CI(n37268), .I0(n16508[1]), .I1(n355_adj_3788), 
            .CO(n37269));
    SB_CARRY unary_minus_70_add_3_11 (.CI(n37058), .I0(GND_net), .I1(n79[9]), 
            .CO(n37059));
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err[2] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [2]));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 unary_minus_70_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n79[8]), 
            .I3(n37057), .O(n868)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err[3] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [3]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err[4] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [4]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err[5] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [5]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err[6] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [6]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err[7] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [7]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err[8] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [8]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err[9] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [9]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err[10] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [10]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err[11] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [11]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err[12] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [12]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err[13] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [13]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err[14] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [14]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err[15] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [15]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err[16] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [16]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err[17] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [17]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err[18] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [18]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err[19] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [19]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err[20] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [20]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err[21] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [21]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err[22] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [22]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i24  (.Q(\PID_CONTROLLER.err[23] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [23]));   // verilog/motorControl.v(31[14] 52[8])
    SB_DFF \PID_CONTROLLER.err_i25  (.Q(\PID_CONTROLLER.err[31] ), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_31__N_2816 [24]));   // verilog/motorControl.v(31[14] 52[8])
    SB_CARRY add_3052_4 (.CI(n38887), .I0(n1798[22]), .I1(n1687), .CO(n38888));
    SB_LUT4 mult_14_add_1211_24_lut (.I0(GND_net), .I1(n1797[21]), .I2(GND_net), 
            .I3(n38681), .O(n1796[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3092_13 (.CI(n38334), .I0(n8211[10]), .I1(GND_net), .CO(n38335));
    SB_LUT4 add_3492_3_lut (.I0(GND_net), .I1(n16508[0]), .I2(n258_adj_3791), 
            .I3(n37267), .O(n16423[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_3 (.CI(n37267), .I0(n16508[0]), .I1(n258_adj_3791), 
            .CO(n37268));
    SB_LUT4 add_3092_12_lut (.I0(GND_net), .I1(n8211[9]), .I2(GND_net), 
            .I3(n38333), .O(n8187[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3092_12 (.CI(n38333), .I0(n8211[9]), .I1(GND_net), .CO(n38334));
    SB_CARRY mult_14_add_1211_24 (.CI(n38681), .I0(n1797[21]), .I1(GND_net), 
            .CO(n1683));
    SB_LUT4 add_3492_2_lut (.I0(GND_net), .I1(n68_adj_3792), .I2(n161_adj_3793), 
            .I3(GND_net), .O(n16423[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3492_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3492_2 (.CI(GND_net), .I0(n68_adj_3792), .I1(n161_adj_3793), 
            .CO(n37267));
    SB_LUT4 add_3092_11_lut (.I0(GND_net), .I1(n8211[8]), .I2(GND_net), 
            .I3(n38332), .O(n8187[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_23_lut (.I0(GND_net), .I1(n1797[20]), .I2(GND_net), 
            .I3(n38680), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_23 (.CI(n38680), .I0(n1797[20]), .I1(GND_net), 
            .CO(n38681));
    SB_CARRY add_3092_11 (.CI(n38332), .I0(n8211[8]), .I1(GND_net), .CO(n38333));
    SB_LUT4 add_3343_21_lut (.I0(GND_net), .I1(n14437[18]), .I2(GND_net), 
            .I3(n37266), .O(n14038[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_10 (.CI(n37057), .I0(GND_net), .I1(n79[8]), 
            .CO(n37058));
    SB_LUT4 add_3343_20_lut (.I0(GND_net), .I1(n14437[17]), .I2(GND_net), 
            .I3(n37265), .O(n14038[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n79[7]), 
            .I3(n37056), .O(n869)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_10_lut (.I0(GND_net), .I1(n8211[7]), .I2(GND_net), 
            .I3(n38331), .O(n8187[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3092_10 (.CI(n38331), .I0(n8211[7]), .I1(GND_net), .CO(n38332));
    SB_LUT4 mult_14_add_1211_22_lut (.I0(GND_net), .I1(n1797[19]), .I2(GND_net), 
            .I3(n38679), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_22 (.CI(n38679), .I0(n1797[19]), .I1(GND_net), 
            .CO(n38680));
    SB_CARRY add_3343_20 (.CI(n37265), .I0(n14437[17]), .I1(GND_net), 
            .CO(n37266));
    SB_CARRY unary_minus_70_add_3_9 (.CI(n37056), .I0(GND_net), .I1(n79[7]), 
            .CO(n37057));
    SB_LUT4 add_3343_19_lut (.I0(GND_net), .I1(n14437[16]), .I2(GND_net), 
            .I3(n37264), .O(n14038[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n79[6]), 
            .I3(n37055), .O(n870)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3052_3_lut (.I0(GND_net), .I1(n1797[22]), .I2(n1683), 
            .I3(n38886), .O(n7068[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_22_lut (.I0(GND_net), .I1(n10674[19]), .I2(GND_net), 
            .I3(n37484), .O(n9932[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_21_lut (.I0(GND_net), .I1(n1797[18]), .I2(GND_net), 
            .I3(n38678), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_9_lut (.I0(GND_net), .I1(n8211[6]), .I2(GND_net), 
            .I3(n38330), .O(n8187[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_19 (.CI(n37264), .I0(n14437[16]), .I1(GND_net), 
            .CO(n37265));
    SB_LUT4 add_3343_18_lut (.I0(GND_net), .I1(n14437[15]), .I2(GND_net), 
            .I3(n37263), .O(n14038[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_18 (.CI(n37263), .I0(n14437[15]), .I1(GND_net), 
            .CO(n37264));
    SB_CARRY unary_minus_70_add_3_8 (.CI(n37055), .I0(GND_net), .I1(n79[6]), 
            .CO(n37056));
    SB_CARRY add_3092_9 (.CI(n38330), .I0(n8211[6]), .I1(GND_net), .CO(n38331));
    SB_CARRY add_3170_22 (.CI(n37484), .I0(n10674[19]), .I1(GND_net), 
            .CO(n37485));
    SB_LUT4 add_3343_17_lut (.I0(GND_net), .I1(n14437[14]), .I2(GND_net), 
            .I3(n37262), .O(n14038[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n79[5]), 
            .I3(n37054), .O(n871)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_7 (.CI(n37054), .I0(GND_net), .I1(n79[5]), 
            .CO(n37055));
    SB_CARRY add_3343_17 (.CI(n37262), .I0(n14437[14]), .I1(GND_net), 
            .CO(n37263));
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3526));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3092_8_lut (.I0(GND_net), .I1(n8211[5]), .I2(n707_adj_3797), 
            .I3(n38329), .O(n8187[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_16_lut (.I0(GND_net), .I1(n14437[13]), .I2(GND_net), 
            .I3(n37261), .O(n14038[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_16 (.CI(n37261), .I0(n14437[13]), .I1(GND_net), 
            .CO(n37262));
    SB_CARRY mult_14_add_1211_21 (.CI(n38678), .I0(n1797[18]), .I1(GND_net), 
            .CO(n38679));
    SB_CARRY add_3092_8 (.CI(n38329), .I0(n8211[5]), .I1(n707_adj_3797), 
            .CO(n38330));
    SB_CARRY add_3052_3 (.CI(n38886), .I0(n1797[22]), .I1(n1683), .CO(n38887));
    SB_DFFE PHASES_i1 (.Q(PIN_6_c_0), .C(clk32MHz), .E(n12_adj_3798), 
            .D(PHASES_5__N_2779[0]));   // verilog/motorControl.v(57[10] 100[6])
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3525));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_DFF Kd_delay_counter_1046__i1 (.Q(Kd_delay_counter[1]), .C(clk32MHz), 
           .D(n69[1]));   // verilog/motorControl.v(48[27:47])
    SB_LUT4 mult_10_i136_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n201_adj_3524));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i235_2_lut (.I0(\Kd[3] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n349_adj_3523));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i235_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i300_2_lut (.I0(\Kd[4] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n446_adj_3522));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_add_1211_20_lut (.I0(GND_net), .I1(n1797[17]), .I2(GND_net), 
            .I3(n38677), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_7_lut (.I0(GND_net), .I1(n8211[4]), .I2(n610_adj_3799), 
            .I3(n38328), .O(n8187[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_15_lut (.I0(GND_net), .I1(n14437[12]), .I2(GND_net), 
            .I3(n37260), .O(n14038[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_15 (.CI(n37260), .I0(n14437[12]), .I1(GND_net), 
            .CO(n37261));
    SB_LUT4 mult_14_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i365_2_lut (.I0(\Kd[5] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n543_adj_3520));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i201_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n298_adj_3519));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i201_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3092_7 (.CI(n38328), .I0(n8211[4]), .I1(n610_adj_3799), 
            .CO(n38329));
    SB_LUT4 add_3343_14_lut (.I0(GND_net), .I1(n14437[11]), .I2(GND_net), 
            .I3(n37259), .O(n14038[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n79[4]), 
            .I3(n37053), .O(n872)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_6_lut (.I0(GND_net), .I1(n8211[3]), .I2(n513_adj_3801), 
            .I3(n38327), .O(n8187[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_14 (.CI(n37259), .I0(n14437[11]), .I1(GND_net), 
            .CO(n37260));
    SB_CARRY unary_minus_70_add_3_6 (.CI(n37053), .I0(GND_net), .I1(n79[4]), 
            .CO(n37054));
    SB_CARRY add_3092_6 (.CI(n38327), .I0(n8211[3]), .I1(n513_adj_3801), 
            .CO(n38328));
    SB_LUT4 add_3343_13_lut (.I0(GND_net), .I1(n14437[10]), .I2(GND_net), 
            .I3(n37258), .O(n14038[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_70_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n79[3]), 
            .I3(n37052), .O(n873)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_5_lut (.I0(GND_net), .I1(n8211[2]), .I2(n416_adj_3803), 
            .I3(n38326), .O(n8187[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i430_2_lut (.I0(\Kd[6] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n640_adj_3518));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i430_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3343_13 (.CI(n37258), .I0(n14437[10]), .I1(GND_net), 
            .CO(n37259));
    SB_CARRY unary_minus_70_add_3_5 (.CI(n37052), .I0(GND_net), .I1(n79[3]), 
            .CO(n37053));
    SB_LUT4 add_3052_2_lut (.I0(GND_net), .I1(n1796[22]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n7068[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3052_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_20 (.CI(n38677), .I0(n1797[17]), .I1(GND_net), 
            .CO(n38678));
    SB_LUT4 mult_12_i495_2_lut (.I0(\Kd[7] ), .I1(n61[19]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_3517));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i495_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n79[2]), 
            .I3(n37051), .O(n874)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_19_lut (.I0(GND_net), .I1(n1797[16]), .I2(GND_net), 
            .I3(n38676), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3092_5 (.CI(n38326), .I0(n8211[2]), .I1(n416_adj_3803), 
            .CO(n38327));
    SB_LUT4 add_3092_4_lut (.I0(GND_net), .I1(n8211[1]), .I2(n319_adj_3805), 
            .I3(n38325), .O(n8187[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3343_12_lut (.I0(GND_net), .I1(n14437[9]), .I2(GND_net), 
            .I3(n37257), .O(n14038[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_12 (.CI(n37257), .I0(n14437[9]), .I1(GND_net), .CO(n37258));
    SB_CARRY add_3092_4 (.CI(n38325), .I0(n8211[1]), .I1(n319_adj_3805), 
            .CO(n38326));
    SB_LUT4 add_3092_3_lut (.I0(GND_net), .I1(n8211[0]), .I2(n222_adj_3806), 
            .I3(n38324), .O(n8187[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i266_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n395_adj_3516));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i266_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3343_11_lut (.I0(GND_net), .I1(n14437[8]), .I2(GND_net), 
            .I3(n37256), .O(n14038[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3170_21_lut (.I0(GND_net), .I1(n10674[18]), .I2(GND_net), 
            .I3(n37483), .O(n9932[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_11 (.CI(n37256), .I0(n14437[8]), .I1(GND_net), .CO(n37257));
    SB_DFF Kd_delay_counter_1046__i2 (.Q(Kd_delay_counter[2]), .C(clk32MHz), 
           .D(n69[2]));   // verilog/motorControl.v(48[27:47])
    SB_CARRY mult_14_add_1211_19 (.CI(n38676), .I0(n1797[16]), .I1(GND_net), 
            .CO(n38677));
    SB_CARRY add_3092_3 (.CI(n38324), .I0(n8211[0]), .I1(n222_adj_3806), 
            .CO(n38325));
    SB_LUT4 mult_10_i331_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n492_adj_3515));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n589_adj_3514));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_DFF Kd_delay_counter_1046__i3 (.Q(Kd_delay_counter[3]), .C(clk32MHz), 
           .D(n69[3]));   // verilog/motorControl.v(48[27:47])
    SB_DFF Kd_delay_counter_1046__i4 (.Q(Kd_delay_counter[4]), .C(clk32MHz), 
           .D(n69[4]));   // verilog/motorControl.v(48[27:47])
    SB_DFF Kd_delay_counter_1046__i5 (.Q(Kd_delay_counter[5]), .C(clk32MHz), 
           .D(n69[5]));   // verilog/motorControl.v(48[27:47])
    SB_DFF Kd_delay_counter_1046__i6 (.Q(Kd_delay_counter[6]), .C(clk32MHz), 
           .D(n69[6]));   // verilog/motorControl.v(48[27:47])
    SB_DFF pwm_count_1047__i1 (.Q(pwm_count[1]), .C(clk32MHz), .D(n73[1]));   // verilog/motorControl.v(99[18:29])
    SB_LUT4 mult_14_add_1211_18_lut (.I0(GND_net), .I1(n1797[15]), .I2(GND_net), 
            .I3(n38675), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3092_2_lut (.I0(GND_net), .I1(n32_adj_3807), .I2(n125_adj_3808), 
            .I3(GND_net), .O(n8187[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3092_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_21 (.CI(n37483), .I0(n10674[18]), .I1(GND_net), 
            .CO(n37484));
    SB_LUT4 add_3343_10_lut (.I0(GND_net), .I1(n14437[7]), .I2(GND_net), 
            .I3(n37255), .O(n14038[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_4 (.CI(n37051), .I0(GND_net), .I1(n79[2]), 
            .CO(n37052));
    SB_LUT4 unary_minus_70_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n79[1]), 
            .I3(n37050), .O(n875)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3092_2 (.CI(GND_net), .I0(n32_adj_3807), .I1(n125_adj_3808), 
            .CO(n38324));
    SB_LUT4 add_3170_20_lut (.I0(GND_net), .I1(n10674[17]), .I2(GND_net), 
            .I3(n37482), .O(n9932[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_10 (.CI(n37255), .I0(n14437[7]), .I1(GND_net), .CO(n37256));
    SB_CARRY unary_minus_70_add_3_3 (.CI(n37050), .I0(GND_net), .I1(n79[1]), 
            .CO(n37051));
    SB_LUT4 unary_minus_70_add_3_2_lut (.I0(n28495), .I1(GND_net), .I2(n79[0]), 
            .I3(VCC_net), .O(n47156)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_70_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3343_9_lut (.I0(GND_net), .I1(n14437[6]), .I2(GND_net), 
            .I3(n37254), .O(n14038[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_9 (.CI(n37254), .I0(n14437[6]), .I1(GND_net), .CO(n37255));
    SB_LUT4 add_3091_24_lut (.I0(GND_net), .I1(n8187[21]), .I2(GND_net), 
            .I3(n38323), .O(n8162[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_8_lut (.I0(GND_net), .I1(n14437[5]), .I2(n713_adj_3811), 
            .I3(n37253), .O(n14038[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_8 (.CI(n37253), .I0(n14437[5]), .I1(n713_adj_3811), 
            .CO(n37254));
    SB_CARRY add_3052_2 (.CI(GND_net), .I0(n1796[22]), .I1(\PID_CONTROLLER.integral [9]), 
            .CO(n38886));
    SB_DFF pwm_count_1047__i2 (.Q(pwm_count[2]), .C(clk32MHz), .D(n73[2]));   // verilog/motorControl.v(99[18:29])
    SB_LUT4 add_3343_7_lut (.I0(GND_net), .I1(n14437[4]), .I2(n616_adj_3812), 
            .I3(n37252), .O(n14038[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_7 (.CI(n37252), .I0(n14437[4]), .I1(n616_adj_3812), 
            .CO(n37253));
    SB_LUT4 add_3109_22_lut (.I0(GND_net), .I1(n9330[19]), .I2(GND_net), 
            .I3(n38885), .O(n8475[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_70_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n79[0]), 
            .CO(n37050));
    SB_CARRY mult_14_add_1211_18 (.CI(n38675), .I0(n1797[15]), .I1(GND_net), 
            .CO(n38676));
    SB_LUT4 add_3091_23_lut (.I0(GND_net), .I1(n8187[20]), .I2(GND_net), 
            .I3(n38322), .O(n8162[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_23 (.CI(n38322), .I0(n8187[20]), .I1(GND_net), .CO(n38323));
    SB_LUT4 mult_14_add_1211_17_lut (.I0(GND_net), .I1(n1797[14]), .I2(GND_net), 
            .I3(n38674), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_22_lut (.I0(GND_net), .I1(n8187[19]), .I2(GND_net), 
            .I3(n38321), .O(n8162[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_20 (.CI(n37482), .I0(n10674[17]), .I1(GND_net), 
            .CO(n37483));
    SB_LUT4 add_3343_6_lut (.I0(GND_net), .I1(n14437[3]), .I2(n519_adj_3813), 
            .I3(n37251), .O(n14038[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_3814), 
            .I3(n37049), .O(n63[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_count_1047__i3 (.Q(pwm_count[3]), .C(clk32MHz), .D(n73[3]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1047__i4 (.Q(pwm_count[4]), .C(clk32MHz), .D(n73[4]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1047__i5 (.Q(pwm_count[5]), .C(clk32MHz), .D(n73[5]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1047__i6 (.Q(pwm_count[6]), .C(clk32MHz), .D(n73[6]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1047__i7 (.Q(pwm_count[7]), .C(clk32MHz), .D(n73[7]));   // verilog/motorControl.v(99[18:29])
    SB_DFF pwm_count_1047__i8 (.Q(pwm_count[8]), .C(clk32MHz), .D(n73[8]));   // verilog/motorControl.v(99[18:29])
    SB_DFFE \PID_CONTROLLER.integral_1048__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[1]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[2]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[3]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[4]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[5]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[6]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[7]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[8]));   // verilog/motorControl.v(34[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1048__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(n55_adj_3646), .D(n70[9]));   // verilog/motorControl.v(34[21:33])
    SB_CARRY mult_14_add_1211_17 (.CI(n38674), .I0(n1797[14]), .I1(GND_net), 
            .CO(n38675));
    SB_CARRY add_3091_22 (.CI(n38321), .I0(n8187[19]), .I1(GND_net), .CO(n38322));
    SB_CARRY add_3343_6 (.CI(n37251), .I0(n14437[3]), .I1(n519_adj_3813), 
            .CO(n37252));
    SB_LUT4 add_3091_21_lut (.I0(GND_net), .I1(n8187[18]), .I2(GND_net), 
            .I3(n38320), .O(n8162[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_5_lut (.I0(GND_net), .I1(n14437[2]), .I2(n422_adj_3815), 
            .I3(n37250), .O(n14038[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_21 (.CI(n38320), .I0(n8187[18]), .I1(GND_net), .CO(n38321));
    SB_LUT4 unary_minus_21_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_3814), 
            .I3(n37048), .O(n63[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_11 (.CI(n37048), .I0(GND_net), .I1(n6_adj_3814), 
            .CO(n37049));
    SB_DFF \PID_CONTROLLER.err_prev__i1  (.Q(\PID_CONTROLLER.err_prev[0] ), 
           .C(clk32MHz), .D(n23743));   // verilog/motorControl.v(31[14] 52[8])
    SB_LUT4 mult_14_add_1211_16_lut (.I0(GND_net), .I1(n1797[13]), .I2(GND_net), 
            .I3(n38673), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n82[8]), 
            .I3(n37047), .O(n63[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3343_5 (.CI(n37250), .I0(n14437[2]), .I1(n422_adj_3815), 
            .CO(n37251));
    SB_LUT4 add_3343_4_lut (.I0(GND_net), .I1(n14437[1]), .I2(n325_adj_3817), 
            .I3(n37249), .O(n14038[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_16 (.CI(n38673), .I0(n1797[13]), .I1(GND_net), 
            .CO(n38674));
    SB_CARRY add_3343_4 (.CI(n37249), .I0(n14437[1]), .I1(n325_adj_3817), 
            .CO(n37250));
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n686_adj_3513));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3109_21_lut (.I0(GND_net), .I1(n9330[18]), .I2(GND_net), 
            .I3(n38884), .O(n8475[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_15_lut (.I0(GND_net), .I1(n1797[12]), .I2(GND_net), 
            .I3(n38672), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_15 (.CI(n38672), .I0(n1797[12]), .I1(GND_net), 
            .CO(n38673));
    SB_CARRY add_3109_21 (.CI(n38884), .I0(n9330[18]), .I1(GND_net), .CO(n38885));
    SB_LUT4 add_3091_20_lut (.I0(GND_net), .I1(n8187[17]), .I2(GND_net), 
            .I3(n38319), .O(n8162[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_20 (.CI(n38319), .I0(n8187[17]), .I1(GND_net), .CO(n38320));
    SB_LUT4 mult_14_add_1211_14_lut (.I0(GND_net), .I1(n1797[11]), .I2(GND_net), 
            .I3(n38671), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_19_lut (.I0(GND_net), .I1(n8187[16]), .I2(GND_net), 
            .I3(n38318), .O(n8162[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_19 (.CI(n38318), .I0(n8187[16]), .I1(GND_net), .CO(n38319));
    SB_CARRY mult_14_add_1211_14 (.CI(n38671), .I0(n1797[11]), .I1(GND_net), 
            .CO(n38672));
    SB_LUT4 add_3109_20_lut (.I0(GND_net), .I1(n9330[17]), .I2(GND_net), 
            .I3(n38883), .O(n8475[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_18_lut (.I0(GND_net), .I1(n8187[15]), .I2(GND_net), 
            .I3(n38317), .O(n8162[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_18 (.CI(n38317), .I0(n8187[15]), .I1(GND_net), .CO(n38318));
    SB_LUT4 mult_14_add_1211_13_lut (.I0(GND_net), .I1(n1797[10]), .I2(GND_net), 
            .I3(n38670), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_17_lut (.I0(GND_net), .I1(n8187[14]), .I2(GND_net), 
            .I3(n38316), .O(n8162[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_17 (.CI(n38316), .I0(n8187[14]), .I1(GND_net), .CO(n38317));
    SB_CARRY mult_14_add_1211_13 (.CI(n38670), .I0(n1797[10]), .I1(GND_net), 
            .CO(n38671));
    SB_CARRY add_3109_20 (.CI(n38883), .I0(n9330[17]), .I1(GND_net), .CO(n38884));
    SB_LUT4 add_3091_16_lut (.I0(GND_net), .I1(n8187[13]), .I2(GND_net), 
            .I3(n38315), .O(n8162[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_16 (.CI(n38315), .I0(n8187[13]), .I1(GND_net), .CO(n38316));
    SB_LUT4 mult_14_add_1211_12_lut (.I0(GND_net), .I1(n1797[9]), .I2(GND_net), 
            .I3(n38669), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_15_lut (.I0(GND_net), .I1(n8187[12]), .I2(GND_net), 
            .I3(n38314), .O(n8162[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_15 (.CI(n38314), .I0(n8187[12]), .I1(GND_net), .CO(n38315));
    SB_CARRY mult_14_add_1211_12 (.CI(n38669), .I0(n1797[9]), .I1(GND_net), 
            .CO(n38670));
    SB_LUT4 add_3109_19_lut (.I0(GND_net), .I1(n9330[16]), .I2(GND_net), 
            .I3(n38882), .O(n8475[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_14_lut (.I0(GND_net), .I1(n8187[11]), .I2(GND_net), 
            .I3(n38313), .O(n8162[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_14 (.CI(n38313), .I0(n8187[11]), .I1(GND_net), .CO(n38314));
    SB_LUT4 mult_14_add_1211_11_lut (.I0(GND_net), .I1(n1797[8]), .I2(GND_net), 
            .I3(n38668), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_13_lut (.I0(GND_net), .I1(n8187[10]), .I2(GND_net), 
            .I3(n38312), .O(n8162[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_13 (.CI(n38312), .I0(n8187[10]), .I1(GND_net), .CO(n38313));
    SB_CARRY mult_14_add_1211_11 (.CI(n38668), .I0(n1797[8]), .I1(GND_net), 
            .CO(n38669));
    SB_CARRY add_3109_19 (.CI(n38882), .I0(n9330[16]), .I1(GND_net), .CO(n38883));
    SB_LUT4 add_3091_12_lut (.I0(GND_net), .I1(n8187[9]), .I2(GND_net), 
            .I3(n38311), .O(n8162[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_12 (.CI(n38311), .I0(n8187[9]), .I1(GND_net), .CO(n38312));
    SB_LUT4 mult_14_add_1211_10_lut (.I0(GND_net), .I1(n1797[7]), .I2(GND_net), 
            .I3(n38667), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_11_lut (.I0(GND_net), .I1(n8187[8]), .I2(GND_net), 
            .I3(n38310), .O(n8162[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_11 (.CI(n38310), .I0(n8187[8]), .I1(GND_net), .CO(n38311));
    SB_CARRY mult_14_add_1211_10 (.CI(n38667), .I0(n1797[7]), .I1(GND_net), 
            .CO(n38668));
    SB_LUT4 add_3109_18_lut (.I0(GND_net), .I1(n9330[15]), .I2(GND_net), 
            .I3(n38881), .O(n8475[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_10_lut (.I0(GND_net), .I1(n8187[7]), .I2(GND_net), 
            .I3(n38309), .O(n8162[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_10 (.CI(n38309), .I0(n8187[7]), .I1(GND_net), .CO(n38310));
    SB_LUT4 mult_14_add_1211_9_lut (.I0(GND_net), .I1(n1797[6]), .I2(GND_net), 
            .I3(n38666), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_9_lut (.I0(GND_net), .I1(n8187[6]), .I2(GND_net), 
            .I3(n38308), .O(n8162[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_9 (.CI(n38308), .I0(n8187[6]), .I1(GND_net), .CO(n38309));
    SB_CARRY mult_14_add_1211_9 (.CI(n38666), .I0(n1797[6]), .I1(GND_net), 
            .CO(n38667));
    SB_CARRY add_3109_18 (.CI(n38881), .I0(n9330[15]), .I1(GND_net), .CO(n38882));
    SB_LUT4 add_3091_8_lut (.I0(GND_net), .I1(n8187[5]), .I2(n704_adj_3818), 
            .I3(n38307), .O(n8162[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_8 (.CI(n38307), .I0(n8187[5]), .I1(n704_adj_3818), 
            .CO(n38308));
    SB_LUT4 mult_14_add_1211_8_lut (.I0(GND_net), .I1(n1797[5]), .I2(n512), 
            .I3(n38665), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_7_lut (.I0(GND_net), .I1(n8187[4]), .I2(n607_adj_3819), 
            .I3(n38306), .O(n8162[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_7 (.CI(n38306), .I0(n8187[4]), .I1(n607_adj_3819), 
            .CO(n38307));
    SB_CARRY mult_14_add_1211_8 (.CI(n38665), .I0(n1797[5]), .I1(n512), 
            .CO(n38666));
    SB_LUT4 add_3109_17_lut (.I0(GND_net), .I1(n9330[14]), .I2(GND_net), 
            .I3(n38880), .O(n8475[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_6_lut (.I0(GND_net), .I1(n8187[3]), .I2(n510_adj_3820), 
            .I3(n38305), .O(n8162[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_6 (.CI(n38305), .I0(n8187[3]), .I1(n510_adj_3820), 
            .CO(n38306));
    SB_LUT4 mult_14_add_1211_7_lut (.I0(GND_net), .I1(n1797[4]), .I2(n439), 
            .I3(n38664), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_5_lut (.I0(GND_net), .I1(n8187[2]), .I2(n413_adj_3821), 
            .I3(n38304), .O(n8162[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_5 (.CI(n38304), .I0(n8187[2]), .I1(n413_adj_3821), 
            .CO(n38305));
    SB_CARRY mult_14_add_1211_7 (.CI(n38664), .I0(n1797[4]), .I1(n439), 
            .CO(n38665));
    SB_CARRY add_3109_17 (.CI(n38880), .I0(n9330[14]), .I1(GND_net), .CO(n38881));
    SB_LUT4 add_3091_4_lut (.I0(GND_net), .I1(n8187[1]), .I2(n316_adj_3822), 
            .I3(n38303), .O(n8162[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_4 (.CI(n38303), .I0(n8187[1]), .I1(n316_adj_3822), 
            .CO(n38304));
    SB_LUT4 mult_14_add_1211_6_lut (.I0(GND_net), .I1(n1797[3]), .I2(n366), 
            .I3(n38663), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_3_lut (.I0(GND_net), .I1(n8187[0]), .I2(n219_adj_3823), 
            .I3(n38302), .O(n8162[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_3 (.CI(n38302), .I0(n8187[0]), .I1(n219_adj_3823), 
            .CO(n38303));
    SB_CARRY mult_14_add_1211_6 (.CI(n38663), .I0(n1797[3]), .I1(n366), 
            .CO(n38664));
    SB_LUT4 add_3109_16_lut (.I0(GND_net), .I1(n9330[13]), .I2(GND_net), 
            .I3(n38879), .O(n8475[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3091_2_lut (.I0(GND_net), .I1(n29_adj_3824), .I2(n122_adj_3825), 
            .I3(GND_net), .O(n8162[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3091_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3091_2 (.CI(GND_net), .I0(n29_adj_3824), .I1(n122_adj_3825), 
            .CO(n38302));
    SB_LUT4 mult_14_add_1211_5_lut (.I0(GND_net), .I1(n1797[2]), .I2(n293), 
            .I3(n38662), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_25_lut (.I0(GND_net), .I1(n8162[22]), .I2(GND_net), 
            .I3(n38301), .O(n8136[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_24_lut (.I0(GND_net), .I1(n8162[21]), .I2(GND_net), 
            .I3(n38300), .O(n8136[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_5 (.CI(n38662), .I0(n1797[2]), .I1(n293), 
            .CO(n38663));
    SB_CARRY add_3109_16 (.CI(n38879), .I0(n9330[13]), .I1(GND_net), .CO(n38880));
    SB_CARRY add_3090_24 (.CI(n38300), .I0(n8162[21]), .I1(GND_net), .CO(n38301));
    SB_LUT4 add_3090_23_lut (.I0(GND_net), .I1(n8162[20]), .I2(GND_net), 
            .I3(n38299), .O(n8136[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_4_lut (.I0(GND_net), .I1(n1797[1]), .I2(n220_adj_3826), 
            .I3(n38661), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_23 (.CI(n38299), .I0(n8162[20]), .I1(GND_net), .CO(n38300));
    SB_LUT4 add_3090_22_lut (.I0(GND_net), .I1(n8162[19]), .I2(GND_net), 
            .I3(n38298), .O(n8136[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_4 (.CI(n38661), .I0(n1797[1]), .I1(n220_adj_3826), 
            .CO(n38662));
    SB_LUT4 add_3109_15_lut (.I0(GND_net), .I1(n9330[12]), .I2(GND_net), 
            .I3(n38878), .O(n8475[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_22 (.CI(n38298), .I0(n8162[19]), .I1(GND_net), .CO(n38299));
    SB_LUT4 add_3090_21_lut (.I0(GND_net), .I1(n8162[18]), .I2(GND_net), 
            .I3(n38297), .O(n8136[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_3_lut (.I0(GND_net), .I1(n1797[0]), .I2(n147_adj_3827), 
            .I3(n38660), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_21 (.CI(n38297), .I0(n8162[18]), .I1(GND_net), .CO(n38298));
    SB_LUT4 add_3090_20_lut (.I0(GND_net), .I1(n8162[17]), .I2(GND_net), 
            .I3(n38296), .O(n8136[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_3 (.CI(n38660), .I0(n1797[0]), .I1(n147_adj_3827), 
            .CO(n38661));
    SB_CARRY add_3109_15 (.CI(n38878), .I0(n9330[12]), .I1(GND_net), .CO(n38879));
    SB_CARRY unary_minus_21_add_3_10 (.CI(n37047), .I0(GND_net), .I1(n82[8]), 
            .CO(n37048));
    SB_LUT4 unary_minus_21_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n82[7]), 
            .I3(n37046), .O(n413)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_3_lut (.I0(GND_net), .I1(n14437[0]), .I2(n228_adj_3829), 
            .I3(n37248), .O(n14038[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_20 (.CI(n38296), .I0(n8162[17]), .I1(GND_net), .CO(n38297));
    SB_CARRY unary_minus_21_add_3_9 (.CI(n37046), .I0(GND_net), .I1(n82[7]), 
            .CO(n37047));
    SB_CARRY add_3343_3 (.CI(n37248), .I0(n14437[0]), .I1(n228_adj_3829), 
            .CO(n37249));
    SB_LUT4 unary_minus_21_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n82[6]), 
            .I3(n37045), .O(n414)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3343_2_lut (.I0(GND_net), .I1(n38_adj_3831), .I2(n131_adj_3832), 
            .I3(GND_net), .O(n14038[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3343_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_19_lut (.I0(GND_net), .I1(n8162[16]), .I2(GND_net), 
            .I3(n38295), .O(n8136[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1211_2_lut (.I0(GND_net), .I1(n5_adj_3833), .I2(n74_adj_3834), 
            .I3(GND_net), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1211_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_8 (.CI(n37045), .I0(GND_net), .I1(n82[6]), 
            .CO(n37046));
    SB_CARRY add_3343_2 (.CI(GND_net), .I0(n38_adj_3831), .I1(n131_adj_3832), 
            .CO(n37248));
    SB_CARRY add_3090_19 (.CI(n38295), .I0(n8162[16]), .I1(GND_net), .CO(n38296));
    SB_LUT4 add_3363_20_lut (.I0(GND_net), .I1(n14796[17]), .I2(GND_net), 
            .I3(n37247), .O(n14437[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3363_19_lut (.I0(GND_net), .I1(n14796[16]), .I2(GND_net), 
            .I3(n37246), .O(n14437[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_18_lut (.I0(GND_net), .I1(n8162[15]), .I2(GND_net), 
            .I3(n38294), .O(n8136[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1211_2 (.CI(GND_net), .I0(n5_adj_3833), .I1(n74_adj_3834), 
            .CO(n38660));
    SB_LUT4 add_3109_14_lut (.I0(GND_net), .I1(n9330[11]), .I2(GND_net), 
            .I3(n38877), .O(n8475[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n82[5]), 
            .I3(n37044), .O(n415)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_7 (.CI(n37044), .I0(GND_net), .I1(n82[5]), 
            .CO(n37045));
    SB_CARRY add_3363_19 (.CI(n37246), .I0(n14796[16]), .I1(GND_net), 
            .CO(n37247));
    SB_LUT4 unary_minus_21_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n82[4]), 
            .I3(n37043), .O(n63[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_6 (.CI(n37043), .I0(GND_net), .I1(n82[4]), 
            .CO(n37044));
    SB_LUT4 add_3363_18_lut (.I0(GND_net), .I1(n14796[15]), .I2(GND_net), 
            .I3(n37245), .O(n14437[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_18 (.CI(n38294), .I0(n8162[15]), .I1(GND_net), .CO(n38295));
    SB_LUT4 unary_minus_21_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n82[3]), 
            .I3(n37042), .O(n63[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_18 (.CI(n37245), .I0(n14796[15]), .I1(GND_net), 
            .CO(n37246));
    SB_CARRY unary_minus_21_add_3_5 (.CI(n37042), .I0(GND_net), .I1(n82[3]), 
            .CO(n37043));
    SB_LUT4 add_3363_17_lut (.I0(GND_net), .I1(n14796[14]), .I2(GND_net), 
            .I3(n37244), .O(n14437[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_17_lut (.I0(GND_net), .I1(n8162[14]), .I2(GND_net), 
            .I3(n38293), .O(n8136[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_18_lut (.I0(GND_net), .I1(n15402[15]), .I2(GND_net), 
            .I3(n38659), .O(n15117[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_21_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n82[2]), 
            .I3(n37041), .O(n63[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_17 (.CI(n37244), .I0(n14796[14]), .I1(GND_net), 
            .CO(n37245));
    SB_CARRY unary_minus_21_add_3_4 (.CI(n37041), .I0(GND_net), .I1(n82[2]), 
            .CO(n37042));
    SB_LUT4 add_3363_16_lut (.I0(GND_net), .I1(n14796[13]), .I2(GND_net), 
            .I3(n37243), .O(n14437[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_17 (.CI(n38293), .I0(n8162[14]), .I1(GND_net), .CO(n38294));
    SB_CARRY add_3363_16 (.CI(n37243), .I0(n14796[13]), .I1(GND_net), 
            .CO(n37244));
    SB_LUT4 add_3363_15_lut (.I0(GND_net), .I1(n14796[12]), .I2(GND_net), 
            .I3(n37242), .O(n14437[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_16_lut (.I0(GND_net), .I1(n8162[13]), .I2(GND_net), 
            .I3(n38292), .O(n8136[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_17_lut (.I0(GND_net), .I1(n15402[14]), .I2(GND_net), 
            .I3(n38658), .O(n15117[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_14 (.CI(n38877), .I0(n9330[11]), .I1(GND_net), .CO(n38878));
    SB_LUT4 add_3170_19_lut (.I0(GND_net), .I1(n10674[16]), .I2(GND_net), 
            .I3(n37481), .O(n9932[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_17 (.CI(n38658), .I0(n15402[14]), .I1(GND_net), 
            .CO(n38659));
    SB_LUT4 add_3400_16_lut (.I0(GND_net), .I1(n15402[13]), .I2(GND_net), 
            .I3(n38657), .O(n15117[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_13_lut (.I0(GND_net), .I1(n9330[10]), .I2(GND_net), 
            .I3(n38876), .O(n8475[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_16 (.CI(n38657), .I0(n15402[13]), .I1(GND_net), 
            .CO(n38658));
    SB_LUT4 add_3400_15_lut (.I0(GND_net), .I1(n15402[12]), .I2(GND_net), 
            .I3(n38656), .O(n15117[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_13 (.CI(n38876), .I0(n9330[10]), .I1(GND_net), .CO(n38877));
    SB_LUT4 unary_minus_21_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n82[1]), 
            .I3(n37040), .O(n63[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_3 (.CI(n37040), .I0(GND_net), .I1(n82[1]), 
            .CO(n37041));
    SB_CARRY add_3363_15 (.CI(n37242), .I0(n14796[12]), .I1(GND_net), 
            .CO(n37243));
    SB_LUT4 unary_minus_21_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n82[0]), 
            .I3(VCC_net), .O(n63[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_21_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_21_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n82[0]), 
            .CO(n37040));
    SB_LUT4 add_3363_14_lut (.I0(GND_net), .I1(n14796[11]), .I2(GND_net), 
            .I3(n37241), .O(n14437[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_16 (.CI(n38292), .I0(n8162[13]), .I1(GND_net), .CO(n38293));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n57[23]), 
            .I3(n37039), .O(n67[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3363_14 (.CI(n37241), .I0(n14796[11]), .I1(GND_net), 
            .CO(n37242));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[22]), .I3(n37038), .O(n45_adj_3843)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3363_13_lut (.I0(GND_net), .I1(n14796[10]), .I2(GND_net), 
            .I3(n37240), .O(n14437[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_15_lut (.I0(GND_net), .I1(n8162[12]), .I2(GND_net), 
            .I3(n38291), .O(n8136[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_15 (.CI(n38656), .I0(n15402[12]), .I1(GND_net), 
            .CO(n38657));
    SB_CARRY unary_minus_5_add_3_24 (.CI(n37038), .I0(GND_net), .I1(n57[22]), 
            .CO(n37039));
    SB_CARRY add_3363_13 (.CI(n37240), .I0(n14796[10]), .I1(GND_net), 
            .CO(n37241));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[21]), .I3(n37037), .O(n43_adj_3845)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3363_12_lut (.I0(GND_net), .I1(n14796[9]), .I2(GND_net), 
            .I3(n37239), .O(n14437[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_15 (.CI(n38291), .I0(n8162[12]), .I1(GND_net), .CO(n38292));
    SB_CARRY add_3363_12 (.CI(n37239), .I0(n14796[9]), .I1(GND_net), .CO(n37240));
    SB_LUT4 add_3363_11_lut (.I0(GND_net), .I1(n14796[8]), .I2(GND_net), 
            .I3(n37238), .O(n14437[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_14_lut (.I0(GND_net), .I1(n8162[11]), .I2(GND_net), 
            .I3(n38290), .O(n8136[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_14_lut (.I0(GND_net), .I1(n15402[11]), .I2(GND_net), 
            .I3(n38655), .O(n15117[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_12_lut (.I0(GND_net), .I1(n9330[9]), .I2(GND_net), 
            .I3(n38875), .O(n8475[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n37037), .I0(GND_net), .I1(n57[21]), 
            .CO(n37038));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[20]), .I3(n37036), .O(n41_adj_3847)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3363_11 (.CI(n37238), .I0(n14796[8]), .I1(GND_net), .CO(n37239));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n37036), .I0(GND_net), .I1(n57[20]), 
            .CO(n37037));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[19]), .I3(n37035), .O(n39_adj_3849)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3363_10_lut (.I0(GND_net), .I1(n14796[7]), .I2(GND_net), 
            .I3(n37237), .O(n14437[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_14 (.CI(n38290), .I0(n8162[11]), .I1(GND_net), .CO(n38291));
    SB_CARRY unary_minus_5_add_3_21 (.CI(n37035), .I0(GND_net), .I1(n57[19]), 
            .CO(n37036));
    SB_CARRY add_3363_10 (.CI(n37237), .I0(n14796[7]), .I1(GND_net), .CO(n37238));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[18]), .I3(n37034), .O(n37_adj_3851)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3363_9_lut (.I0(GND_net), .I1(n14796[6]), .I2(GND_net), 
            .I3(n37236), .O(n14437[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_13_lut (.I0(GND_net), .I1(n8162[10]), .I2(GND_net), 
            .I3(n38289), .O(n8136[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_14 (.CI(n38655), .I0(n15402[11]), .I1(GND_net), 
            .CO(n38656));
    SB_CARRY unary_minus_5_add_3_20 (.CI(n37034), .I0(GND_net), .I1(n57[18]), 
            .CO(n37035));
    SB_CARRY add_3363_9 (.CI(n37236), .I0(n14796[6]), .I1(GND_net), .CO(n37237));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n57[17]), .I3(n37033), .O(n35_adj_3853)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3363_8_lut (.I0(GND_net), .I1(n14796[5]), .I2(n716_adj_3854), 
            .I3(n37235), .O(n14437[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_13 (.CI(n38289), .I0(n8162[10]), .I1(GND_net), .CO(n38290));
    SB_CARRY add_3363_8 (.CI(n37235), .I0(n14796[5]), .I1(n716_adj_3854), 
            .CO(n37236));
    SB_LUT4 add_3363_7_lut (.I0(GND_net), .I1(n14796[4]), .I2(n619), .I3(n37234), 
            .O(n14437[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3363_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_12_lut (.I0(GND_net), .I1(n8162[9]), .I2(GND_net), 
            .I3(n38288), .O(n8136[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_13_lut (.I0(GND_net), .I1(n15402[10]), .I2(GND_net), 
            .I3(n38654), .O(n15117[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_12 (.CI(n38875), .I0(n9330[9]), .I1(GND_net), .CO(n38876));
    SB_CARRY add_3400_13 (.CI(n38654), .I0(n15402[10]), .I1(GND_net), 
            .CO(n38655));
    SB_LUT4 add_3400_12_lut (.I0(GND_net), .I1(n15402[9]), .I2(GND_net), 
            .I3(n38653), .O(n15117[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_11_lut (.I0(GND_net), .I1(n9330[8]), .I2(GND_net), 
            .I3(n38874), .O(n8475[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_12 (.CI(n38653), .I0(n15402[9]), .I1(GND_net), .CO(n38654));
    SB_LUT4 add_3400_11_lut (.I0(GND_net), .I1(n15402[8]), .I2(GND_net), 
            .I3(n38652), .O(n15117[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_11 (.CI(n38874), .I0(n9330[8]), .I1(GND_net), .CO(n38875));
    SB_CARRY add_3170_19 (.CI(n37481), .I0(n10674[16]), .I1(GND_net), 
            .CO(n37482));
    SB_LUT4 add_3170_18_lut (.I0(GND_net), .I1(n10674[15]), .I2(GND_net), 
            .I3(n37480), .O(n9932[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_12 (.CI(n38288), .I0(n8162[9]), .I1(GND_net), .CO(n38289));
    SB_CARRY add_3170_18 (.CI(n37480), .I0(n10674[15]), .I1(GND_net), 
            .CO(n37481));
    SB_LUT4 add_3170_17_lut (.I0(GND_net), .I1(n10674[14]), .I2(GND_net), 
            .I3(n37479), .O(n9932[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_11_lut (.I0(GND_net), .I1(n8162[8]), .I2(GND_net), 
            .I3(n38287), .O(n8136[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_11 (.CI(n38652), .I0(n15402[8]), .I1(GND_net), .CO(n38653));
    SB_CARRY add_3170_17 (.CI(n37479), .I0(n10674[14]), .I1(GND_net), 
            .CO(n37480));
    SB_LUT4 add_3170_16_lut (.I0(GND_net), .I1(n10674[13]), .I2(GND_net), 
            .I3(n37478), .O(n9932[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_11 (.CI(n38287), .I0(n8162[8]), .I1(GND_net), .CO(n38288));
    SB_CARRY add_3170_16 (.CI(n37478), .I0(n10674[13]), .I1(GND_net), 
            .CO(n37479));
    SB_LUT4 add_3170_15_lut (.I0(GND_net), .I1(n10674[12]), .I2(GND_net), 
            .I3(n37477), .O(n9932[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_10_lut (.I0(GND_net), .I1(n8162[7]), .I2(GND_net), 
            .I3(n38286), .O(n8136[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_10_lut (.I0(GND_net), .I1(n15402[7]), .I2(GND_net), 
            .I3(n38651), .O(n15117[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_10_lut (.I0(GND_net), .I1(n9330[7]), .I2(GND_net), 
            .I3(n38873), .O(n8475[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_15 (.CI(n37477), .I0(n10674[12]), .I1(GND_net), 
            .CO(n37478));
    SB_LUT4 add_3170_14_lut (.I0(GND_net), .I1(n10674[11]), .I2(GND_net), 
            .I3(n37476), .O(n9932[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_10 (.CI(n38286), .I0(n8162[7]), .I1(GND_net), .CO(n38287));
    SB_CARRY add_3170_14 (.CI(n37476), .I0(n10674[11]), .I1(GND_net), 
            .CO(n37477));
    SB_LUT4 add_3170_13_lut (.I0(GND_net), .I1(n10674[10]), .I2(GND_net), 
            .I3(n37475), .O(n9932[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_9_lut (.I0(GND_net), .I1(n8162[6]), .I2(GND_net), 
            .I3(n38285), .O(n8136[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_10 (.CI(n38651), .I0(n15402[7]), .I1(GND_net), .CO(n38652));
    SB_CARRY add_3170_13 (.CI(n37475), .I0(n10674[10]), .I1(GND_net), 
            .CO(n37476));
    SB_LUT4 add_3170_12_lut (.I0(GND_net), .I1(n10674[9]), .I2(GND_net), 
            .I3(n37474), .O(n9932[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_9 (.CI(n38285), .I0(n8162[6]), .I1(GND_net), .CO(n38286));
    SB_CARRY add_3170_12 (.CI(n37474), .I0(n10674[9]), .I1(GND_net), .CO(n37475));
    SB_LUT4 add_3170_11_lut (.I0(GND_net), .I1(n10674[8]), .I2(GND_net), 
            .I3(n37473), .O(n9932[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_8_lut (.I0(GND_net), .I1(n8162[5]), .I2(n701_adj_3855), 
            .I3(n38284), .O(n8136[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_9_lut (.I0(GND_net), .I1(n15402[6]), .I2(GND_net), 
            .I3(n38650), .O(n15117[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_10 (.CI(n38873), .I0(n9330[7]), .I1(GND_net), .CO(n38874));
    SB_CARRY add_3170_11 (.CI(n37473), .I0(n10674[8]), .I1(GND_net), .CO(n37474));
    SB_LUT4 add_3170_10_lut (.I0(GND_net), .I1(n10674[7]), .I2(GND_net), 
            .I3(n37472), .O(n9932[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_10 (.CI(n37472), .I0(n10674[7]), .I1(GND_net), .CO(n37473));
    SB_LUT4 add_3170_9_lut (.I0(GND_net), .I1(n10674[6]), .I2(GND_net), 
            .I3(n37471), .O(n9932[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_9 (.CI(n38650), .I0(n15402[6]), .I1(GND_net), .CO(n38651));
    SB_CARRY add_3170_9 (.CI(n37471), .I0(n10674[6]), .I1(GND_net), .CO(n37472));
    SB_LUT4 add_3170_8_lut (.I0(GND_net), .I1(n10674[5]), .I2(n692_adj_3856), 
            .I3(n37470), .O(n9932[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_8 (.CI(n37470), .I0(n10674[5]), .I1(n692_adj_3856), 
            .CO(n37471));
    SB_LUT4 add_3170_7_lut (.I0(GND_net), .I1(n10674[4]), .I2(n595_adj_3857), 
            .I3(n37469), .O(n9932[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_8_lut (.I0(GND_net), .I1(n15402[5]), .I2(n722_adj_3858), 
            .I3(n38649), .O(n15117[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_9_lut (.I0(GND_net), .I1(n9330[6]), .I2(GND_net), 
            .I3(n38872), .O(n8475[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_7 (.CI(n37469), .I0(n10674[4]), .I1(n595_adj_3857), 
            .CO(n37470));
    SB_LUT4 add_3170_6_lut (.I0(GND_net), .I1(n10674[3]), .I2(n498_adj_3859), 
            .I3(n37468), .O(n9932[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_6 (.CI(n37468), .I0(n10674[3]), .I1(n498_adj_3859), 
            .CO(n37469));
    SB_LUT4 add_3170_5_lut (.I0(GND_net), .I1(n10674[2]), .I2(n401_adj_3860), 
            .I3(n37467), .O(n9932[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_8 (.CI(n38649), .I0(n15402[5]), .I1(n722_adj_3858), 
            .CO(n38650));
    SB_CARRY add_3170_5 (.CI(n37467), .I0(n10674[2]), .I1(n401_adj_3860), 
            .CO(n37468));
    SB_LUT4 add_3170_4_lut (.I0(GND_net), .I1(n10674[1]), .I2(n304_adj_3861), 
            .I3(n37466), .O(n9932[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3170_4 (.CI(n37466), .I0(n10674[1]), .I1(n304_adj_3861), 
            .CO(n37467));
    SB_LUT4 add_3170_3_lut (.I0(GND_net), .I1(n10674[0]), .I2(n207_adj_3862), 
            .I3(n37465), .O(n9932[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_7_lut (.I0(GND_net), .I1(n15402[4]), .I2(n625_adj_3863), 
            .I3(n38648), .O(n15117[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_9 (.CI(n38872), .I0(n9330[6]), .I1(GND_net), .CO(n38873));
    SB_CARRY add_3170_3 (.CI(n37465), .I0(n10674[0]), .I1(n207_adj_3862), 
            .CO(n37466));
    SB_LUT4 add_3170_2_lut (.I0(GND_net), .I1(n17_adj_3864), .I2(n110_adj_3865), 
            .I3(GND_net), .O(n9932[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3170_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_8 (.CI(n38284), .I0(n8162[5]), .I1(n701_adj_3855), 
            .CO(n38285));
    SB_CARRY add_3170_2 (.CI(GND_net), .I0(n17_adj_3864), .I1(n110_adj_3865), 
            .CO(n37465));
    SB_LUT4 add_3350_13_lut (.I0(GND_net), .I1(n14563[10]), .I2(GND_net), 
            .I3(n37464), .O(n14171[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_7_lut (.I0(GND_net), .I1(n8162[4]), .I2(n604_adj_3866), 
            .I3(n38283), .O(n8136[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_7 (.CI(n38648), .I0(n15402[4]), .I1(n625_adj_3863), 
            .CO(n38649));
    SB_LUT4 add_3350_12_lut (.I0(GND_net), .I1(n14563[9]), .I2(GND_net), 
            .I3(n37463), .O(n14171[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_12 (.CI(n37463), .I0(n14563[9]), .I1(GND_net), .CO(n37464));
    SB_CARRY add_3090_7 (.CI(n38283), .I0(n8162[4]), .I1(n604_adj_3866), 
            .CO(n38284));
    SB_LUT4 add_3350_11_lut (.I0(GND_net), .I1(n14563[8]), .I2(GND_net), 
            .I3(n37462), .O(n14171[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_11 (.CI(n37462), .I0(n14563[8]), .I1(GND_net), .CO(n37463));
    SB_LUT4 add_3090_6_lut (.I0(GND_net), .I1(n8162[3]), .I2(n507_adj_3867), 
            .I3(n38282), .O(n8136[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_6_lut (.I0(GND_net), .I1(n15402[3]), .I2(n528_adj_3868), 
            .I3(n38647), .O(n15117[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_8_lut (.I0(GND_net), .I1(n9330[5]), .I2(n545), .I3(n38871), 
            .O(n8475[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3350_10_lut (.I0(GND_net), .I1(n14563[7]), .I2(GND_net), 
            .I3(n37461), .O(n14171[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_10 (.CI(n37461), .I0(n14563[7]), .I1(GND_net), .CO(n37462));
    SB_CARRY add_3090_6 (.CI(n38282), .I0(n8162[3]), .I1(n507_adj_3867), 
            .CO(n38283));
    SB_LUT4 add_3350_9_lut (.I0(GND_net), .I1(n14563[6]), .I2(GND_net), 
            .I3(n37460), .O(n14171[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_9 (.CI(n37460), .I0(n14563[6]), .I1(GND_net), .CO(n37461));
    SB_LUT4 add_3090_5_lut (.I0(GND_net), .I1(n8162[2]), .I2(n410_adj_3869), 
            .I3(n38281), .O(n8136[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_6 (.CI(n38647), .I0(n15402[3]), .I1(n528_adj_3868), 
            .CO(n38648));
    SB_LUT4 add_3350_8_lut (.I0(GND_net), .I1(n14563[5]), .I2(n545), .I3(n37459), 
            .O(n14171[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_8 (.CI(n37459), .I0(n14563[5]), .I1(n545), .CO(n37460));
    SB_CARRY add_3090_5 (.CI(n38281), .I0(n8162[2]), .I1(n410_adj_3869), 
            .CO(n38282));
    SB_LUT4 add_3350_7_lut (.I0(GND_net), .I1(n14563[4]), .I2(n472), .I3(n37458), 
            .O(n14171[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3090_4_lut (.I0(GND_net), .I1(n8162[1]), .I2(n313_adj_3870), 
            .I3(n38280), .O(n8136[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_5_lut (.I0(GND_net), .I1(n15402[2]), .I2(n431_adj_3871), 
            .I3(n38646), .O(n15117[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_8 (.CI(n38871), .I0(n9330[5]), .I1(n545), .CO(n38872));
    SB_CARRY add_3350_7 (.CI(n37458), .I0(n14563[4]), .I1(n472), .CO(n37459));
    SB_LUT4 add_3350_6_lut (.I0(GND_net), .I1(n14563[3]), .I2(n399), .I3(n37457), 
            .O(n14171[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_6 (.CI(n37457), .I0(n14563[3]), .I1(n399), .CO(n37458));
    SB_LUT4 add_3350_5_lut (.I0(GND_net), .I1(n14563[2]), .I2(n326), .I3(n37456), 
            .O(n14171[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_5 (.CI(n38646), .I0(n15402[2]), .I1(n431_adj_3871), 
            .CO(n38647));
    SB_CARRY add_3350_5 (.CI(n37456), .I0(n14563[2]), .I1(n326), .CO(n37457));
    SB_LUT4 add_3350_4_lut (.I0(GND_net), .I1(n14563[1]), .I2(n253), .I3(n37455), 
            .O(n14171[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_4 (.CI(n37455), .I0(n14563[1]), .I1(n253), .CO(n37456));
    SB_LUT4 add_3350_3_lut (.I0(GND_net), .I1(n14563[0]), .I2(n180), .I3(n37454), 
            .O(n14171[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_4_lut (.I0(GND_net), .I1(n15402[1]), .I2(n334_adj_3872), 
            .I3(n38645), .O(n15117[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_7_lut (.I0(GND_net), .I1(n9330[4]), .I2(n472), .I3(n38870), 
            .O(n8475[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_3 (.CI(n37454), .I0(n14563[0]), .I1(n180), .CO(n37455));
    SB_LUT4 add_3350_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n14171[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3350_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3350_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n37454));
    SB_LUT4 add_3198_27_lut (.I0(GND_net), .I1(n11361[24]), .I2(GND_net), 
            .I3(n37453), .O(n10674[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_4 (.CI(n38645), .I0(n15402[1]), .I1(n334_adj_3872), 
            .CO(n38646));
    SB_LUT4 add_3198_26_lut (.I0(GND_net), .I1(n11361[23]), .I2(GND_net), 
            .I3(n37452), .O(n10674[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_26 (.CI(n37452), .I0(n11361[23]), .I1(GND_net), 
            .CO(n37453));
    SB_LUT4 add_3198_25_lut (.I0(GND_net), .I1(n11361[22]), .I2(GND_net), 
            .I3(n37451), .O(n10674[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3198_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3198_25 (.CI(n37451), .I0(n11361[22]), .I1(GND_net), 
            .CO(n37452));
    SB_LUT4 add_3400_3_lut (.I0(GND_net), .I1(n15402[0]), .I2(n237_adj_3873), 
            .I3(n38644), .O(n15117[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_7 (.CI(n38870), .I0(n9330[4]), .I1(n472), .CO(n38871));
    SB_CARRY add_3090_4 (.CI(n38280), .I0(n8162[1]), .I1(n313_adj_3870), 
            .CO(n38281));
    SB_LUT4 add_3090_3_lut (.I0(GND_net), .I1(n8162[0]), .I2(n216_adj_3874), 
            .I3(n38279), .O(n8136[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_3 (.CI(n38644), .I0(n15402[0]), .I1(n237_adj_3873), 
            .CO(n38645));
    SB_CARRY add_3090_3 (.CI(n38279), .I0(n8162[0]), .I1(n216_adj_3874), 
            .CO(n38280));
    SB_LUT4 add_3090_2_lut (.I0(GND_net), .I1(n26_adj_3875), .I2(n119_adj_3876), 
            .I3(GND_net), .O(n8136[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3090_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3400_2_lut (.I0(GND_net), .I1(n47_adj_3877), .I2(n140_adj_3878), 
            .I3(GND_net), .O(n15117[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3400_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3109_6_lut (.I0(GND_net), .I1(n9330[3]), .I2(n399), .I3(n38869), 
            .O(n8475[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3090_2 (.CI(GND_net), .I0(n26_adj_3875), .I1(n119_adj_3876), 
            .CO(n38279));
    SB_LUT4 add_3089_26_lut (.I0(GND_net), .I1(n8136[23]), .I2(GND_net), 
            .I3(n38278), .O(n8109[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3400_2 (.CI(GND_net), .I0(n47_adj_3877), .I1(n140_adj_3878), 
            .CO(n38644));
    SB_LUT4 add_3089_25_lut (.I0(GND_net), .I1(n8136[22]), .I2(GND_net), 
            .I3(n38277), .O(n8109[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_25 (.CI(n38277), .I0(n8136[22]), .I1(GND_net), .CO(n38278));
    SB_LUT4 add_3509_9_lut (.I0(GND_net), .I1(n16623[6]), .I2(GND_net), 
            .I3(n38643), .O(n16574[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_6 (.CI(n38869), .I0(n9330[3]), .I1(n399), .CO(n38870));
    SB_LUT4 add_3509_8_lut (.I0(GND_net), .I1(n16623[5]), .I2(n749_adj_3879), 
            .I3(n38642), .O(n16574[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_8 (.CI(n38642), .I0(n16623[5]), .I1(n749_adj_3879), 
            .CO(n38643));
    SB_LUT4 add_3109_5_lut (.I0(GND_net), .I1(n9330[2]), .I2(n326), .I3(n38868), 
            .O(n8475[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3509_7_lut (.I0(GND_net), .I1(n16623[4]), .I2(n652_adj_3880), 
            .I3(n38641), .O(n16574[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_7 (.CI(n38641), .I0(n16623[4]), .I1(n652_adj_3880), 
            .CO(n38642));
    SB_CARRY add_3109_5 (.CI(n38868), .I0(n9330[2]), .I1(n326), .CO(n38869));
    SB_LUT4 add_3089_24_lut (.I0(GND_net), .I1(n8136[21]), .I2(GND_net), 
            .I3(n38276), .O(n8109[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_24 (.CI(n38276), .I0(n8136[21]), .I1(GND_net), .CO(n38277));
    SB_LUT4 add_3509_6_lut (.I0(GND_net), .I1(n16623[3]), .I2(n555_adj_3881), 
            .I3(n38640), .O(n16574[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_23_lut (.I0(GND_net), .I1(n8136[20]), .I2(GND_net), 
            .I3(n38275), .O(n8109[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_23 (.CI(n38275), .I0(n8136[20]), .I1(GND_net), .CO(n38276));
    SB_CARRY add_3509_6 (.CI(n38640), .I0(n16623[3]), .I1(n555_adj_3881), 
            .CO(n38641));
    SB_LUT4 add_3109_4_lut (.I0(GND_net), .I1(n9330[1]), .I2(n253), .I3(n38867), 
            .O(n8475[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_22_lut (.I0(GND_net), .I1(n8136[19]), .I2(GND_net), 
            .I3(n38274), .O(n8109[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_22 (.CI(n38274), .I0(n8136[19]), .I1(GND_net), .CO(n38275));
    SB_LUT4 add_3509_5_lut (.I0(GND_net), .I1(n16623[2]), .I2(n458_adj_3882), 
            .I3(n38639), .O(n16574[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_21_lut (.I0(GND_net), .I1(n8136[18]), .I2(GND_net), 
            .I3(n38273), .O(n8109[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_21 (.CI(n38273), .I0(n8136[18]), .I1(GND_net), .CO(n38274));
    SB_CARRY add_3509_5 (.CI(n38639), .I0(n16623[2]), .I1(n458_adj_3882), 
            .CO(n38640));
    SB_CARRY add_3109_4 (.CI(n38867), .I0(n9330[1]), .I1(n253), .CO(n38868));
    SB_LUT4 add_3509_4_lut (.I0(GND_net), .I1(n16623[1]), .I2(n361_adj_3883), 
            .I3(n38638), .O(n16574[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_4 (.CI(n38638), .I0(n16623[1]), .I1(n361_adj_3883), 
            .CO(n38639));
    SB_LUT4 add_3109_3_lut (.I0(GND_net), .I1(n9330[0]), .I2(n180), .I3(n38866), 
            .O(n8475[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3509_3_lut (.I0(GND_net), .I1(n16623[0]), .I2(n264_adj_3884), 
            .I3(n38637), .O(n16574[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3509_3 (.CI(n38637), .I0(n16623[0]), .I1(n264_adj_3884), 
            .CO(n38638));
    SB_CARRY add_3109_3 (.CI(n38866), .I0(n9330[0]), .I1(n180), .CO(n38867));
    SB_LUT4 add_3089_20_lut (.I0(GND_net), .I1(n8136[17]), .I2(GND_net), 
            .I3(n38272), .O(n8109[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_20 (.CI(n38272), .I0(n8136[17]), .I1(GND_net), .CO(n38273));
    SB_LUT4 add_3509_2_lut (.I0(GND_net), .I1(n86), .I2(n167_adj_3885), 
            .I3(GND_net), .O(n16574[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3509_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_19_lut (.I0(GND_net), .I1(n8136[16]), .I2(GND_net), 
            .I3(n38271), .O(n8109[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_19 (.CI(n38271), .I0(n8136[16]), .I1(GND_net), .CO(n38272));
    SB_CARRY add_3509_2 (.CI(GND_net), .I0(n86), .I1(n167_adj_3885), .CO(n38637));
    SB_LUT4 add_3109_2_lut (.I0(GND_net), .I1(n35), .I2(n107_adj_3418), 
            .I3(GND_net), .O(n8475[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3109_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_18_lut (.I0(GND_net), .I1(n8136[15]), .I2(GND_net), 
            .I3(n38270), .O(n8109[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_18 (.CI(n38270), .I0(n8136[15]), .I1(GND_net), .CO(n38271));
    SB_LUT4 add_3417_17_lut (.I0(GND_net), .I1(n15643[14]), .I2(GND_net), 
            .I3(n38636), .O(n15402[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_17_lut (.I0(GND_net), .I1(n8136[14]), .I2(GND_net), 
            .I3(n38269), .O(n8109[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_17 (.CI(n38269), .I0(n8136[14]), .I1(GND_net), .CO(n38270));
    SB_LUT4 add_3417_16_lut (.I0(GND_net), .I1(n15643[13]), .I2(GND_net), 
            .I3(n38635), .O(n15402[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3109_2 (.CI(GND_net), .I0(n35), .I1(n107_adj_3418), .CO(n38866));
    SB_LUT4 add_3089_16_lut (.I0(GND_net), .I1(n8136[13]), .I2(GND_net), 
            .I3(n38268), .O(n8109[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_16 (.CI(n38268), .I0(n8136[13]), .I1(GND_net), .CO(n38269));
    SB_CARRY add_3417_16 (.CI(n38635), .I0(n15643[13]), .I1(GND_net), 
            .CO(n38636));
    SB_LUT4 add_3089_15_lut (.I0(GND_net), .I1(n8136[12]), .I2(GND_net), 
            .I3(n38267), .O(n8109[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_15 (.CI(n38267), .I0(n8136[12]), .I1(GND_net), .CO(n38268));
    SB_LUT4 add_3417_15_lut (.I0(GND_net), .I1(n15643[12]), .I2(GND_net), 
            .I3(n38634), .O(n15402[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_24_lut (.I0(GND_net), .I1(n8451[21]), .I2(GND_net), 
            .I3(n38865), .O(n1804[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_14_lut (.I0(GND_net), .I1(n8136[11]), .I2(GND_net), 
            .I3(n38266), .O(n8109[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_14 (.CI(n38266), .I0(n8136[11]), .I1(GND_net), .CO(n38267));
    SB_CARRY add_3417_15 (.CI(n38634), .I0(n15643[12]), .I1(GND_net), 
            .CO(n38635));
    SB_LUT4 add_3089_13_lut (.I0(GND_net), .I1(n8136[10]), .I2(GND_net), 
            .I3(n38265), .O(n8109[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_13 (.CI(n38265), .I0(n8136[10]), .I1(GND_net), .CO(n38266));
    SB_LUT4 add_3417_14_lut (.I0(GND_net), .I1(n15643[11]), .I2(GND_net), 
            .I3(n38633), .O(n15402[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_23_lut (.I0(GND_net), .I1(n8451[20]), .I2(GND_net), 
            .I3(n38864), .O(n1804[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_12_lut (.I0(GND_net), .I1(n8136[9]), .I2(GND_net), 
            .I3(n38264), .O(n8109[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_12 (.CI(n38264), .I0(n8136[9]), .I1(GND_net), .CO(n38265));
    SB_CARRY add_3417_14 (.CI(n38633), .I0(n15643[11]), .I1(GND_net), 
            .CO(n38634));
    SB_LUT4 add_3089_11_lut (.I0(GND_net), .I1(n8136[8]), .I2(GND_net), 
            .I3(n38263), .O(n8109[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_11 (.CI(n38263), .I0(n8136[8]), .I1(GND_net), .CO(n38264));
    SB_LUT4 add_3417_13_lut (.I0(GND_net), .I1(n15643[10]), .I2(GND_net), 
            .I3(n38632), .O(n15402[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_23 (.CI(n38864), .I0(n8451[20]), .I1(GND_net), 
            .CO(n38865));
    SB_LUT4 add_3089_10_lut (.I0(GND_net), .I1(n8136[7]), .I2(GND_net), 
            .I3(n38262), .O(n8109[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_10 (.CI(n38262), .I0(n8136[7]), .I1(GND_net), .CO(n38263));
    SB_CARRY add_3417_13 (.CI(n38632), .I0(n15643[10]), .I1(GND_net), 
            .CO(n38633));
    SB_LUT4 add_3089_9_lut (.I0(GND_net), .I1(n8136[6]), .I2(GND_net), 
            .I3(n38261), .O(n8109[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_9 (.CI(n38261), .I0(n8136[6]), .I1(GND_net), .CO(n38262));
    SB_LUT4 add_3417_12_lut (.I0(GND_net), .I1(n15643[9]), .I2(GND_net), 
            .I3(n38631), .O(n15402[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_22_lut (.I0(GND_net), .I1(n8451[19]), .I2(GND_net), 
            .I3(n38863), .O(n1804[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3089_8_lut (.I0(GND_net), .I1(n8136[5]), .I2(n698_adj_3886), 
            .I3(n38260), .O(n8109[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_8 (.CI(n38260), .I0(n8136[5]), .I1(n698_adj_3886), 
            .CO(n38261));
    SB_CARRY add_3417_12 (.CI(n38631), .I0(n15643[9]), .I1(GND_net), .CO(n38632));
    SB_LUT4 add_3089_7_lut (.I0(GND_net), .I1(n8136[4]), .I2(n601_adj_3887), 
            .I3(n38259), .O(n8109[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_7 (.CI(n38259), .I0(n8136[4]), .I1(n601_adj_3887), 
            .CO(n38260));
    SB_LUT4 add_3417_11_lut (.I0(GND_net), .I1(n15643[8]), .I2(GND_net), 
            .I3(n38630), .O(n15402[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_22 (.CI(n38863), .I0(n8451[19]), .I1(GND_net), 
            .CO(n38864));
    SB_LUT4 add_3089_6_lut (.I0(GND_net), .I1(n8136[3]), .I2(n504_adj_3888), 
            .I3(n38258), .O(n8109[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_6 (.CI(n38258), .I0(n8136[3]), .I1(n504_adj_3888), 
            .CO(n38259));
    SB_CARRY add_3417_11 (.CI(n38630), .I0(n15643[8]), .I1(GND_net), .CO(n38631));
    SB_LUT4 add_3089_5_lut (.I0(GND_net), .I1(n8136[2]), .I2(n407_adj_3889), 
            .I3(n38257), .O(n8109[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_10_lut (.I0(GND_net), .I1(n15643[7]), .I2(GND_net), 
            .I3(n38629), .O(n15402[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_21_lut (.I0(GND_net), .I1(n8451[18]), .I2(GND_net), 
            .I3(n38862), .O(n1804[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_10 (.CI(n38629), .I0(n15643[7]), .I1(GND_net), .CO(n38630));
    SB_LUT4 add_3417_9_lut (.I0(GND_net), .I1(n15643[6]), .I2(GND_net), 
            .I3(n38628), .O(n15402[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_21 (.CI(n38862), .I0(n8451[18]), .I1(GND_net), 
            .CO(n38863));
    SB_CARRY add_3417_9 (.CI(n38628), .I0(n15643[6]), .I1(GND_net), .CO(n38629));
    SB_LUT4 add_3417_8_lut (.I0(GND_net), .I1(n15643[5]), .I2(n725_adj_3890), 
            .I3(n38627), .O(n15402[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_20_lut (.I0(GND_net), .I1(n8451[17]), .I2(GND_net), 
            .I3(n38861), .O(n1804[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_8 (.CI(n38627), .I0(n15643[5]), .I1(n725_adj_3890), 
            .CO(n38628));
    SB_LUT4 add_3417_7_lut (.I0(GND_net), .I1(n15643[4]), .I2(n628_adj_3891), 
            .I3(n38626), .O(n15402[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_20 (.CI(n38861), .I0(n8451[17]), .I1(GND_net), 
            .CO(n38862));
    SB_CARRY add_3417_7 (.CI(n38626), .I0(n15643[4]), .I1(n628_adj_3891), 
            .CO(n38627));
    SB_LUT4 add_3417_6_lut (.I0(GND_net), .I1(n15643[3]), .I2(n531_adj_3892), 
            .I3(n38625), .O(n15402[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_19_lut (.I0(GND_net), .I1(n8451[16]), .I2(GND_net), 
            .I3(n38860), .O(n1804[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3089_5 (.CI(n38257), .I0(n8136[2]), .I1(n407_adj_3889), 
            .CO(n38258));
    SB_LUT4 add_3089_4_lut (.I0(GND_net), .I1(n8136[1]), .I2(n310_adj_3893), 
            .I3(n38256), .O(n8109[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_6 (.CI(n38625), .I0(n15643[3]), .I1(n531_adj_3892), 
            .CO(n38626));
    SB_CARRY add_3089_4 (.CI(n38256), .I0(n8136[1]), .I1(n310_adj_3893), 
            .CO(n38257));
    SB_LUT4 add_3089_3_lut (.I0(GND_net), .I1(n8136[0]), .I2(n213_adj_3894), 
            .I3(n38255), .O(n8109[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_5_lut (.I0(GND_net), .I1(n15643[2]), .I2(n434_adj_3895), 
            .I3(n38624), .O(n15402[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_19 (.CI(n38860), .I0(n8451[16]), .I1(GND_net), 
            .CO(n38861));
    SB_CARRY add_3089_3 (.CI(n38255), .I0(n8136[0]), .I1(n213_adj_3894), 
            .CO(n38256));
    SB_LUT4 add_3089_2_lut (.I0(GND_net), .I1(n23_adj_3896), .I2(n116_adj_3897), 
            .I3(GND_net), .O(n8109[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3089_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3417_5 (.CI(n38624), .I0(n15643[2]), .I1(n434_adj_3895), 
            .CO(n38625));
    SB_CARRY add_3089_2 (.CI(GND_net), .I0(n23_adj_3896), .I1(n116_adj_3897), 
            .CO(n38255));
    SB_LUT4 add_3088_27_lut (.I0(GND_net), .I1(n8109[24]), .I2(GND_net), 
            .I3(n38254), .O(n8081[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3417_4_lut (.I0(GND_net), .I1(n15643[1]), .I2(n337_adj_3898), 
            .I3(n38623), .O(n15402[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_18_lut (.I0(GND_net), .I1(n8451[15]), .I2(GND_net), 
            .I3(n38859), .O(n1804[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_26_lut (.I0(GND_net), .I1(n8109[23]), .I2(GND_net), 
            .I3(n38253), .O(n8081[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_26 (.CI(n38253), .I0(n8109[23]), .I1(GND_net), .CO(n38254));
    SB_CARRY add_3417_4 (.CI(n38623), .I0(n15643[1]), .I1(n337_adj_3898), 
            .CO(n38624));
    SB_LUT4 add_3088_25_lut (.I0(GND_net), .I1(n8109[22]), .I2(GND_net), 
            .I3(n38252), .O(n8081[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_25 (.CI(n38252), .I0(n8109[22]), .I1(GND_net), .CO(n38253));
    SB_LUT4 add_3417_3_lut (.I0(GND_net), .I1(n15643[0]), .I2(n240_adj_3899), 
            .I3(n38622), .O(n15402[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_18 (.CI(n38859), .I0(n8451[15]), .I1(GND_net), 
            .CO(n38860));
    SB_LUT4 add_3088_24_lut (.I0(GND_net), .I1(n8109[21]), .I2(GND_net), 
            .I3(n38251), .O(n8081[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_24 (.CI(n38251), .I0(n8109[21]), .I1(GND_net), .CO(n38252));
    SB_CARRY add_3417_3 (.CI(n38622), .I0(n15643[0]), .I1(n240_adj_3899), 
            .CO(n38623));
    SB_LUT4 add_3088_23_lut (.I0(GND_net), .I1(n8109[20]), .I2(GND_net), 
            .I3(n38250), .O(n8081[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_23 (.CI(n38250), .I0(n8109[20]), .I1(GND_net), .CO(n38251));
    SB_LUT4 add_3417_2_lut (.I0(GND_net), .I1(n50_adj_3900), .I2(n143_adj_3901), 
            .I3(GND_net), .O(n15402[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3417_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_17_lut (.I0(GND_net), .I1(n8451[14]), .I2(GND_net), 
            .I3(n38858), .O(n1804[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_22_lut (.I0(GND_net), .I1(n8109[19]), .I2(GND_net), 
            .I3(n38249), .O(n8081[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_22 (.CI(n38249), .I0(n8109[19]), .I1(GND_net), .CO(n38250));
    SB_CARRY add_3417_2 (.CI(GND_net), .I0(n50_adj_3900), .I1(n143_adj_3901), 
            .CO(n38622));
    SB_LUT4 add_3088_21_lut (.I0(GND_net), .I1(n8109[18]), .I2(GND_net), 
            .I3(n38248), .O(n8081[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_21 (.CI(n38248), .I0(n8109[18]), .I1(GND_net), .CO(n38249));
    SB_LUT4 add_3517_7_lut (.I0(GND_net), .I1(n44573), .I2(n658), .I3(n38621), 
            .O(n16632[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_17 (.CI(n38858), .I0(n8451[14]), .I1(GND_net), 
            .CO(n38859));
    SB_LUT4 add_3088_20_lut (.I0(GND_net), .I1(n8109[17]), .I2(GND_net), 
            .I3(n38247), .O(n8081[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_20 (.CI(n38247), .I0(n8109[17]), .I1(GND_net), .CO(n38248));
    SB_LUT4 add_3517_6_lut (.I0(GND_net), .I1(n16640[3]), .I2(n558), .I3(n38620), 
            .O(n16632[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_19_lut (.I0(GND_net), .I1(n8109[16]), .I2(GND_net), 
            .I3(n38246), .O(n8081[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_19 (.CI(n38246), .I0(n8109[16]), .I1(GND_net), .CO(n38247));
    SB_CARRY add_3517_6 (.CI(n38620), .I0(n16640[3]), .I1(n558), .CO(n38621));
    SB_LUT4 mult_14_add_1219_16_lut (.I0(GND_net), .I1(n8451[13]), .I2(GND_net), 
            .I3(n38857), .O(n1804[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_18_lut (.I0(GND_net), .I1(n8109[15]), .I2(GND_net), 
            .I3(n38245), .O(n8081[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_18 (.CI(n38245), .I0(n8109[15]), .I1(GND_net), .CO(n38246));
    SB_LUT4 add_3517_5_lut (.I0(GND_net), .I1(n16647[2]), .I2(n464_adj_3377), 
            .I3(n38619), .O(n16632[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_17_lut (.I0(GND_net), .I1(n8109[14]), .I2(GND_net), 
            .I3(n38244), .O(n8081[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_17 (.CI(n38244), .I0(n8109[14]), .I1(GND_net), .CO(n38245));
    SB_CARRY add_3517_5 (.CI(n38619), .I0(n16647[2]), .I1(n464_adj_3377), 
            .CO(n38620));
    SB_CARRY mult_14_add_1219_16 (.CI(n38857), .I0(n8451[13]), .I1(GND_net), 
            .CO(n38858));
    SB_LUT4 add_3088_16_lut (.I0(GND_net), .I1(n8109[13]), .I2(GND_net), 
            .I3(n38243), .O(n8081[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_16 (.CI(n38243), .I0(n8109[13]), .I1(GND_net), .CO(n38244));
    SB_LUT4 add_3517_4_lut (.I0(GND_net), .I1(n16653[1]), .I2(n370), .I3(n38618), 
            .O(n16632[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_15_lut (.I0(GND_net), .I1(n8109[12]), .I2(GND_net), 
            .I3(n38242), .O(n8081[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_15 (.CI(n38242), .I0(n8109[12]), .I1(GND_net), .CO(n38243));
    SB_CARRY add_3517_4 (.CI(n38618), .I0(n16653[1]), .I1(n370), .CO(n38619));
    SB_LUT4 mult_14_add_1219_15_lut (.I0(GND_net), .I1(n8451[12]), .I2(GND_net), 
            .I3(n38856), .O(n1804[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_14_lut (.I0(GND_net), .I1(n8109[11]), .I2(GND_net), 
            .I3(n38241), .O(n8081[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_14 (.CI(n38241), .I0(n8109[11]), .I1(GND_net), .CO(n38242));
    SB_LUT4 add_3517_3_lut (.I0(GND_net), .I1(n16640[0]), .I2(n276), .I3(n38617), 
            .O(n16632[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_13_lut (.I0(GND_net), .I1(n8109[10]), .I2(GND_net), 
            .I3(n38240), .O(n8081[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_13 (.CI(n38240), .I0(n8109[10]), .I1(GND_net), .CO(n38241));
    SB_CARRY add_3517_3 (.CI(n38617), .I0(n16640[0]), .I1(n276), .CO(n38618));
    SB_CARRY mult_14_add_1219_15 (.CI(n38856), .I0(n8451[12]), .I1(GND_net), 
            .CO(n38857));
    SB_LUT4 add_3088_12_lut (.I0(GND_net), .I1(n8109[9]), .I2(GND_net), 
            .I3(n38239), .O(n8081[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_12 (.CI(n38239), .I0(n8109[9]), .I1(GND_net), .CO(n38240));
    SB_LUT4 add_3517_2_lut (.I0(GND_net), .I1(n86), .I2(n182), .I3(GND_net), 
            .O(n16632[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3517_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_11_lut (.I0(GND_net), .I1(n8109[8]), .I2(GND_net), 
            .I3(n38238), .O(n8081[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_11 (.CI(n38238), .I0(n8109[8]), .I1(GND_net), .CO(n38239));
    SB_CARRY add_3517_2 (.CI(GND_net), .I0(n86), .I1(n182), .CO(n38617));
    SB_LUT4 mult_14_add_1219_14_lut (.I0(GND_net), .I1(n8451[11]), .I2(GND_net), 
            .I3(n38855), .O(n1804[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_10_lut (.I0(GND_net), .I1(n8109[7]), .I2(GND_net), 
            .I3(n38237), .O(n8081[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_10 (.CI(n38237), .I0(n8109[7]), .I1(GND_net), .CO(n38238));
    SB_LUT4 add_3432_16_lut (.I0(GND_net), .I1(n15853[13]), .I2(GND_net), 
            .I3(n38616), .O(n15643[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3088_9_lut (.I0(GND_net), .I1(n8109[6]), .I2(GND_net), 
            .I3(n38236), .O(n8081[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_9 (.CI(n38236), .I0(n8109[6]), .I1(GND_net), .CO(n38237));
    SB_LUT4 add_3432_15_lut (.I0(GND_net), .I1(n15853[12]), .I2(GND_net), 
            .I3(n38615), .O(n15643[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_14_add_1219_14 (.CI(n38855), .I0(n8451[11]), .I1(GND_net), 
            .CO(n38856));
    SB_LUT4 add_3088_8_lut (.I0(GND_net), .I1(n8109[5]), .I2(n695_adj_3902), 
            .I3(n38235), .O(n8081[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_8 (.CI(n38235), .I0(n8109[5]), .I1(n695_adj_3902), 
            .CO(n38236));
    SB_CARRY add_3432_15 (.CI(n38615), .I0(n15853[12]), .I1(GND_net), 
            .CO(n38616));
    SB_LUT4 add_3088_7_lut (.I0(GND_net), .I1(n8109[4]), .I2(n598_adj_3903), 
            .I3(n38234), .O(n8081[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3088_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3088_7 (.CI(n38234), .I0(n8109[4]), .I1(n598_adj_3903), 
            .CO(n38235));
    SB_LUT4 add_3432_14_lut (.I0(GND_net), .I1(n15853[11]), .I2(GND_net), 
            .I3(n38614), .O(n15643[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3432_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_14_add_1219_13_lut (.I0(GND_net), .I1(n8451[10]), .I2(GND_net), 
            .I3(n38854), .O(n1804[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_14_add_1219_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_12_i107_2_lut (.I0(\Kd[1] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n158));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i44_2_lut (.I0(\Kd[0] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n65));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i172_2_lut (.I0(\Kd[2] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n255));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i237_2_lut (.I0(\Kd[3] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n352));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i302_2_lut (.I0(\Kd[4] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n449));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i367_2_lut (.I0(\Kd[5] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n546));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i432_2_lut (.I0(\Kd[6] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n643));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i497_2_lut (.I0(\Kd[7] ), .I1(n61[20]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i109_2_lut (.I0(\Kd[1] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n161));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i46_2_lut (.I0(\Kd[0] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n68));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[0]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i174_2_lut (.I0(\Kd[2] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n258));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i239_2_lut (.I0(\Kd[3] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n355));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i304_2_lut (.I0(\Kd[4] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n452));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i369_2_lut (.I0(\Kd[5] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n549));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i434_2_lut (.I0(\Kd[6] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n646));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i499_2_lut (.I0(\Kd[7] ), .I1(n61[21]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i111_2_lut (.I0(\Kd[1] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n164_adj_3507));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i111_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i48_2_lut (.I0(\Kd[0] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n71_adj_3506));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i48_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[1]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i176_2_lut (.I0(\Kd[2] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n261_adj_3504));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i176_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[2]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[3]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i241_2_lut (.I0(\Kd[3] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n358_adj_3499));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i241_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[4]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[5]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i306_2_lut (.I0(\Kd[4] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n455_adj_3494));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[6]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i371_2_lut (.I0(\Kd[5] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n552_adj_3491));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3490));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[7]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i436_2_lut (.I0(\Kd[6] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n649_adj_3487));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i436_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_3486));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3485));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i442_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[6] ), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3484));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i505_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i505_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i142_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n210_adj_3483));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i501_2_lut (.I0(\Kd[7] ), .I1(n61[22]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_3482));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i501_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i207_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n307_adj_3481));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i272_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n404_adj_3480));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_3479));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i99_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n146));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i99_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[17] ), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i337_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n501_adj_3477));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i113_2_lut (.I0(\Kd[1] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n167));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i50_2_lut (.I0(\Kd[0] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i50_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n598));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i178_2_lut (.I0(\Kd[2] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n264));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n695));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i243_2_lut (.I0(\Kd[3] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n361));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[8]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i308_2_lut (.I0(\Kd[4] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n458_c));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i373_2_lut (.I0(\Kd[5] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n555));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3471));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i438_2_lut (.I0(\Kd[6] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n652));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i199_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n295));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i199_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i503_2_lut (.I0(\Kd[7] ), .I1(n61[23]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i264_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n392));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i264_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i402_2_lut (.I0(\Kd[6] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n598_adj_3903));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i467_2_lut (.I0(\Kd[7] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n695_adj_3902));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1418 (.I0(n36452), .I1(n16647[2]), .I2(n464_adj_3377), 
            .I3(n6_adj_3904), .O(n9_adj_3905));   // verilog/motorControl.v(36[17:23])
    defparam i3_4_lut_adj_1418.LUT_INIT = 16'h566a;
    SB_LUT4 i1_3_lut_4_lut (.I0(n16647[2]), .I1(\Kp[4] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n6_adj_3904), .O(n16640[3]));   // verilog/motorControl.v(36[17:23])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h956a;
    SB_LUT4 i5_4_lut (.I0(n9_adj_3905), .I1(n7_adj_3906), .I2(n558), .I3(n43578), 
            .O(n44573));   // verilog/motorControl.v(36[17:23])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i97_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n143_adj_3901));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i97_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3900));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i162_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n240_adj_3899));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i162_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i227_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n337_adj_3898));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i227_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i164_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n243));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i79_2_lut (.I0(\Kd[1] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_3897));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i229_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n340));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i16_2_lut (.I0(\Kd[0] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3896));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i292_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n434_adj_3895));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i292_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i144_2_lut (.I0(\Kd[2] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n213_adj_3894));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i209_2_lut (.I0(\Kd[3] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n310_adj_3893));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i209_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n531_adj_3892));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n628_adj_3891));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i294_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n437));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i294_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_c));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i487_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n725_adj_3890));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i487_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i274_2_lut (.I0(\Kd[4] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n407_adj_3889));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i274_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i339_2_lut (.I0(\Kd[5] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n504_adj_3888));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i339_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i329_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n489));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i329_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i404_2_lut (.I0(\Kd[6] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n601_adj_3887));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i469_2_lut (.I0(\Kd[7] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n698_adj_3886));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i113_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n167_adj_3885));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i178_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n264_adj_3884));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i178_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n534));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n631));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i243_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n361_adj_3883));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i243_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n458_adj_3882));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n555_adj_3881));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i438_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n652_adj_3880));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i438_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i503_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[23] ), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_3879));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i77_2_lut (.I0(\Kd[1] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i95_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n140_adj_3878));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i95_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[15] ), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3877));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i14_2_lut (.I0(\Kd[0] ), .I1(n61[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_c));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i489_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[16] ), 
            .I2(GND_net), .I3(GND_net), .O(n728));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i489_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i81_2_lut (.I0(\Kd[1] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_3876));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[15]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i18_2_lut (.I0(\Kd[0] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_3875));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i146_2_lut (.I0(\Kd[2] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n216_adj_3874));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i160_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n237_adj_3873));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i160_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i225_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n334_adj_3872));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i225_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i290_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n431_adj_3871));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i290_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i211_2_lut (.I0(\Kd[3] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n313_adj_3870));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i276_2_lut (.I0(\Kd[4] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n410_adj_3869));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i276_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n528_adj_3868));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i341_2_lut (.I0(\Kd[5] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n507_adj_3867));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i341_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i406_2_lut (.I0(\Kd[6] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n604_adj_3866));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3865));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i142_2_lut (.I0(\Kd[2] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n210));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[5] ), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3864));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n625_adj_3863));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n586));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i140_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n207_adj_3862));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i205_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n304_adj_3861));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i205_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i270_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n401_adj_3860));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i270_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i115_2_lut (.I0(\Kd[1] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n170));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i115_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i335_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n498_adj_3859));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i335_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i485_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[14] ), 
            .I2(GND_net), .I3(GND_net), .O(n722_adj_3858));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n595_adj_3857));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n692_adj_3856));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i471_2_lut (.I0(\Kd[7] ), .I1(n61[7]), .I2(GND_net), 
            .I3(GND_net), .O(n701_adj_3855));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n683_adj_3468));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i207_2_lut (.I0(\Kd[3] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n307));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i481_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n716_adj_3854));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[18]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i286_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n425));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[19]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[20]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[21]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[22]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[23]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i1_1_lut (.I0(\PWMLimit[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[0]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i2_1_lut (.I0(\PWMLimit[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[1]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i180_2_lut (.I0(\Kd[2] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n267));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i180_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[16]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n57[17]));   // verilog/motorControl.v(33[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i3_1_lut (.I0(\PWMLimit[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[2]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i4_1_lut (.I0(\PWMLimit[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[3]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i81_2_lut (.I0(n880), .I1(hall3), .I2(GND_net), .I3(GND_net), 
            .O(n892));   // verilog/motorControl.v(81[10:35])
    defparam i81_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n522));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_21_inv_0_i5_1_lut (.I0(\PWMLimit[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[4]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_21_inv_0_i6_1_lut (.I0(\PWMLimit[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[5]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n619));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3834));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6294_2_lut_3_lut (.I0(n911), .I1(hall3), .I2(n19566), .I3(GND_net), 
            .O(n19600));   // verilog/motorControl.v(90[10:34])
    defparam i6294_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i2_3_lut_4_lut (.I0(n911), .I1(hall3), .I2(n934), .I3(n19566), 
            .O(n22310));   // verilog/motorControl.v(90[10:34])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfff8;
    SB_LUT4 mult_12_i272_2_lut (.I0(\Kd[4] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n404));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i272_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3833));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_3832));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[12] ), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3831));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23299_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(n61[25]), 
            .I3(GND_net), .O(n10114[0]));   // verilog/motorControl.v(36[26:45])
    defparam i23299_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i6479_2_lut (.I0(hall3), .I1(hall1), .I2(GND_net), .I3(GND_net), 
            .O(n19608));   // verilog/motorControl.v(93[7] 95[10])
    defparam i6479_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 unary_minus_21_inv_0_i7_1_lut (.I0(\PWMLimit[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[6]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i154_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n228_adj_3829));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut (.I0(hall2), .I1(n19608), .I2(GND_net), .I3(GND_net), 
            .O(n934));   // verilog/motorControl.v(93[10:35])
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 unary_minus_21_inv_0_i8_1_lut (.I0(\PWMLimit[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[7]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_3827));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_3826));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i83_2_lut (.I0(\Kd[1] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_3825));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i73_3_lut (.I0(pwm[23]), .I1(n29), .I2(n30), .I3(GND_net), 
            .O(n878));   // verilog/motorControl.v(77[19:44])
    defparam i73_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 mult_12_i20_2_lut (.I0(\Kd[0] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3824));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i148_2_lut (.I0(\Kd[2] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n219_adj_3823));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i213_2_lut (.I0(\Kd[3] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n316_adj_3822));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i278_2_lut (.I0(\Kd[4] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n413_adj_3821));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i88_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n911));   // verilog/motorControl.v(87[10:25])
    defparam i88_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i343_2_lut (.I0(\Kd[5] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n510_adj_3820));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i408_2_lut (.I0(\Kd[6] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n607_adj_3819));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i473_2_lut (.I0(\Kd[7] ), .I1(n61[8]), .I2(GND_net), 
            .I3(GND_net), .O(n704_adj_3818));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23242_2_lut_3_lut (.I0(\Kd[0] ), .I1(\Kd[1] ), .I2(\Kd[2] ), 
            .I3(GND_net), .O(n36747));   // verilog/motorControl.v(36[26:45])
    defparam i23242_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6010_2_lut (.I0(hall3), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n19292));   // verilog/motorControl.v(87[7] 89[10])
    defparam i6010_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_10_i219_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n325_adj_3817));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_1419 (.I0(hall1), .I1(n19292), .I2(GND_net), 
            .I3(GND_net), .O(n902_adj_3909));   // verilog/motorControl.v(84[10:34])
    defparam i2_2_lut_adj_1419.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1420 (.I0(n370_adj_3463), .I1(n4_adj_3910), 
            .I2(n36747), .I3(n61[25]), .O(n7_adj_3911));   // verilog/motorControl.v(36[26:45])
    defparam i1_3_lut_4_lut_adj_1420.LUT_INIT = 16'h6966;
    SB_LUT4 unary_minus_21_inv_0_i9_1_lut (.I0(\PWMLimit[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n82[8]));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i284_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n422_adj_3815));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i9_4_lut (.I0(pwm[16]), .I1(pwm[9]), .I2(pwm[10]), .I3(n48778), 
            .O(n24_adj_3912));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1421 (.I0(pwm[22]), .I1(pwm[17]), .I2(pwm[19]), 
            .I3(pwm[12]), .O(n26_adj_3913));
    defparam i11_4_lut_adj_1421.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1422 (.I0(pwm[21]), .I1(pwm[14]), .I2(pwm[11]), 
            .I3(pwm[13]), .O(n25_adj_3914));
    defparam i10_4_lut_adj_1422.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1423 (.I0(pwm[15]), .I1(n24_adj_3912), .I2(pwm[18]), 
            .I3(pwm[20]), .O(n27_adj_3915));
    defparam i12_4_lut_adj_1423.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1424 (.I0(pwm[23]), .I1(n27_adj_3915), .I2(n25_adj_3914), 
            .I3(n26_adj_3913), .O(n17_adj_3916));   // verilog/motorControl.v(58[9:32])
    defparam i1_4_lut_adj_1424.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_21_inv_0_i32_1_lut (.I0(\PWMLimit[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3814));   // verilog/motorControl.v(40[28:37])
    defparam unary_minus_21_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n519_adj_3813));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n616_adj_3812));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i75_2_lut (.I0(hall1), .I1(hall2), .I2(GND_net), .I3(GND_net), 
            .O(n880));   // verilog/motorControl.v(78[10:25])
    defparam i75_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mult_10_i479_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n713_adj_3811));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1425 (.I0(n880), .I1(n17_adj_3916), .I2(n20352), 
            .I3(n902_adj_3909), .O(n44847));
    defparam i3_4_lut_adj_1425.LUT_INIT = 16'hfffb;
    SB_LUT4 i15093_1_lut (.I0(pwm_count[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n28495));   // verilog/motorControl.v(99[18:29])
    defparam i15093_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i1_1_lut (.I0(pwm[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[0]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i2_1_lut (.I0(pwm[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[1]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1426 (.I0(n19292), .I1(n44847), .I2(n6_adj_3917), 
            .I3(n17_adj_3916), .O(n23569));
    defparam i1_4_lut_adj_1426.LUT_INIT = 16'hccc8;
    SB_LUT4 mult_12_i85_2_lut (.I0(\Kd[1] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_3808));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i22_2_lut (.I0(\Kd[0] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_3807));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 PHASES_5__I_0_i2_4_lut (.I0(n20352), .I1(PHASES_5__N_3039[1]), 
            .I2(n17_adj_3916), .I3(n902_adj_3909), .O(PHASES_5__N_2779[1]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i2_4_lut.LUT_INIT = 16'h5c0c;
    SB_LUT4 mult_12_i150_2_lut (.I0(\Kd[2] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n222_adj_3806));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i215_2_lut (.I0(\Kd[3] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n319_adj_3805));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i3_1_lut (.I0(pwm[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[2]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i280_2_lut (.I0(\Kd[4] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n416_adj_3803));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i4_1_lut (.I0(pwm[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[3]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i345_2_lut (.I0(\Kd[5] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n513_adj_3801));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i117_2_lut (.I0(\Kd[1] ), .I1(n61[25]), .I2(GND_net), 
            .I3(GND_net), .O(n182_adj_3466));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i117_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i182_2_lut (.I0(\Kd[2] ), .I1(n61[25]), .I2(GND_net), 
            .I3(GND_net), .O(n276_adj_3464));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i182_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i5_1_lut (.I0(pwm[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[4]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i410_2_lut (.I0(\Kd[6] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n610_adj_3799));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i245_2_lut (.I0(\Kd[3] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n364));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i245_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i310_2_lut (.I0(\Kd[4] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n461_adj_3461));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i52_2_lut (.I0(\Kd[0] ), .I1(n61[25]), .I2(GND_net), 
            .I3(GND_net), .O(n86_adj_3465));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i52_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut (.I0(n47234), .I1(n44840), .I2(n17_adj_3916), .I3(n6_adj_3917), 
            .O(n12_adj_3798));
    defparam i20_4_lut.LUT_INIT = 16'hfc5c;
    SB_LUT4 i31838_2_lut (.I0(PHASES_5__N_3039[1]), .I1(n878), .I2(GND_net), 
            .I3(GND_net), .O(n47079));   // verilog/motorControl.v(77[14] 98[8])
    defparam i31838_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 PHASES_5__I_0_i1_4_lut (.I0(n47079), .I1(n16801), .I2(n17_adj_3916), 
            .I3(n902_adj_3909), .O(PHASES_5__N_2779[0]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i1_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i2_4_lut_adj_1427 (.I0(\Kd[2] ), .I1(\Kd[0] ), .I2(n61[25]), 
            .I3(\Kd[1] ), .O(n4_adj_3910));   // verilog/motorControl.v(36[26:45])
    defparam i2_4_lut_adj_1427.LUT_INIT = 16'ha080;
    SB_LUT4 mult_12_i247_2_lut (.I0(\Kd[3] ), .I1(n61[25]), .I2(GND_net), 
            .I3(GND_net), .O(n370_adj_3463));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23301_3_lut (.I0(n61[25]), .I1(n36732), .I2(n36747), .I3(GND_net), 
            .O(n11529[1]));   // verilog/motorControl.v(36[26:45])
    defparam i23301_3_lut.LUT_INIT = 16'h6c6c;
    SB_LUT4 mult_12_i475_2_lut (.I0(\Kd[7] ), .I1(n61[9]), .I2(GND_net), 
            .I3(GND_net), .O(n707_adj_3797));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i312_2_lut (.I0(\Kd[4] ), .I1(n61[25]), .I2(GND_net), 
            .I3(GND_net), .O(n464_adj_3462));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i379_2_lut (.I0(\Kd[5] ), .I1(n61[25]), .I2(GND_net), 
            .I3(GND_net), .O(n564));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i379_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i442_2_lut (.I0(\Kd[6] ), .I1(n61[25]), .I2(GND_net), 
            .I3(GND_net), .O(n658_adj_3459));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i442_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i6_1_lut (.I0(pwm[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[5]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut_adj_1428 (.I0(n36732), .I1(n7_adj_3911), .I2(n8_adj_3918), 
            .I3(n8_adj_3919), .O(n44998));   // verilog/motorControl.v(36[26:45])
    defparam i5_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 mult_12_i375_2_lut (.I0(\Kd[5] ), .I1(n61[24]), .I2(GND_net), 
            .I3(GND_net), .O(n558_adj_3456));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i7_1_lut (.I0(pwm[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[6]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i8_1_lut (.I0(pwm[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[7]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i109_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n161_adj_3793));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i109_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i46_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[22] ), 
            .I2(GND_net), .I3(GND_net), .O(n68_adj_3792));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i46_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i174_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n258_adj_3791));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i174_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i9_1_lut (.I0(pwm[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[8]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i10_1_lut (.I0(pwm[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n79[9]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i239_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n355_adj_3788));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i239_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3787));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i11_1_lut (.I0(pwm[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[10]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i12_1_lut (.I0(pwm[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[11]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n452_adj_3784));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34453_4_lut (.I0(n47229), .I1(n44015), .I2(n19600), .I3(n17_adj_3916), 
            .O(n43194));
    defparam i34453_4_lut.LUT_INIT = 16'hddfc;
    SB_LUT4 PHASES_5__I_0_i6_4_lut (.I0(PHASES_5__N_3039[4]), .I1(n22310), 
            .I2(n17_adj_3916), .I3(n878), .O(PHASES_5__N_2779[5]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i6_4_lut.LUT_INIT = 16'ha303;
    SB_LUT4 i1_4_lut_adj_1429 (.I0(n892), .I1(n934), .I2(n911), .I3(n902_adj_3909), 
            .O(PHASES_5__N_3039[4]));
    defparam i1_4_lut_adj_1429.LUT_INIT = 16'h3032;
    SB_LUT4 i28542_3_lut (.I0(n911), .I1(hall3), .I2(hall1), .I3(GND_net), 
            .O(n44039));
    defparam i28542_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i32425_2_lut (.I0(n19600), .I1(n878), .I2(GND_net), .I3(GND_net), 
            .O(n47230));
    defparam i32425_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i34455_4_lut (.I0(n47230), .I1(n44015), .I2(n44039), .I3(n17_adj_3916), 
            .O(n43196));
    defparam i34455_4_lut.LUT_INIT = 16'hddfc;
    SB_LUT4 PHASES_5__I_0_i5_4_lut (.I0(n878), .I1(PHASES_5__N_3039[4]), 
            .I2(n17_adj_3916), .I3(n22310), .O(PHASES_5__N_2779[4]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i5_4_lut.LUT_INIT = 16'h0cac;
    SB_LUT4 i18_4_lut_adj_1430 (.I0(n44079), .I1(n44081), .I2(n17_adj_3916), 
            .I3(n878), .O(n10_adj_3783));
    defparam i18_4_lut_adj_1430.LUT_INIT = 16'hacfc;
    SB_LUT4 PHASES_5__I_0_i4_4_lut (.I0(n47192), .I1(n19608), .I2(n17_adj_3916), 
            .I3(n19292), .O(PHASES_5__N_2779[3]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i4_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i6580_3_lut (.I0(hall3), .I1(hall1), .I2(hall2), .I3(GND_net), 
            .O(n19566));   // verilog/motorControl.v(68[7] 70[10])
    defparam i6580_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i28519_3_lut (.I0(n934), .I1(n880), .I2(hall3), .I3(GND_net), 
            .O(n44015));
    defparam i28519_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i28582_2_lut (.I0(n19600), .I1(n44015), .I2(GND_net), .I3(GND_net), 
            .O(n44079));
    defparam i28582_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1431 (.I0(n19615), .I1(n44079), .I2(n17_adj_3916), 
            .I3(n44011), .O(n10_adj_3782));
    defparam i18_4_lut_adj_1431.LUT_INIT = 16'hfcac;
    SB_LUT4 PHASES_5__I_0_i3_4_lut (.I0(n19615), .I1(PHASES_5__N_3039[2]), 
            .I2(n17_adj_3916), .I3(n19292), .O(PHASES_5__N_2779[2]));   // verilog/motorControl.v(77[14] 98[8])
    defparam PHASES_5__I_0_i3_4_lut.LUT_INIT = 16'h5c0c;
    SB_LUT4 unary_minus_70_inv_0_i13_1_lut (.I0(pwm[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[12]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_3779));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n549_adj_3777));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i14_1_lut (.I0(pwm[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[13]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i434_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n646_adj_3774));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i434_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i15_1_lut (.I0(pwm[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[14]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_3772));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i16_1_lut (.I0(pwm[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[15]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i499_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_3769));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i499_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i17_1_lut (.I0(pwm[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[16]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i18_1_lut (.I0(pwm[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[17]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i19_1_lut (.I0(pwm[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[18]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_3764));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i20_1_lut (.I0(pwm[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[19]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_70_inv_0_i21_1_lut (.I0(pwm[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[20]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i1_3_lut (.I0(\PID_CONTROLLER.result [0]), .I1(n63[0]), 
            .I2(n421), .I3(GND_net), .O(n471));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i87_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n128_adj_3757));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[11] ), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3756));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i2_3_lut (.I0(\PID_CONTROLLER.result [1]), .I1(n63[1]), 
            .I2(n421), .I3(GND_net), .O(n470));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i3_3_lut (.I0(\PID_CONTROLLER.result [2]), .I1(n63[2]), 
            .I2(n421), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i152_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n225_adj_3755));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_70_inv_0_i22_1_lut (.I0(pwm[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[21]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_24_i4_3_lut (.I0(\PID_CONTROLLER.result [3]), .I1(n63[3]), 
            .I2(n421), .I3(GND_net), .O(n468));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i5_3_lut (.I0(\PID_CONTROLLER.result [4]), .I1(n63[4]), 
            .I2(n421), .I3(GND_net), .O(n467));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1432 (.I0(pwm_23__N_2948), .I1(n1), .I2(\PWMLimit[5] ), 
            .I3(n387), .O(n24366));   // verilog/motorControl.v(37[10:51])
    defparam i1_4_lut_adj_1432.LUT_INIT = 16'ha088;
    SB_LUT4 i1_4_lut_adj_1433 (.I0(pwm_23__N_2948), .I1(n28052), .I2(\PWMLimit[6] ), 
            .I3(n387), .O(n24367));   // verilog/motorControl.v(37[10:51])
    defparam i1_4_lut_adj_1433.LUT_INIT = 16'ha088;
    SB_LUT4 mult_10_i217_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n322_adj_3752));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1434 (.I0(pwm_23__N_2948), .I1(n1_adj_16), .I2(\PWMLimit[7] ), 
            .I3(n387), .O(n24368));   // verilog/motorControl.v(37[10:51])
    defparam i1_4_lut_adj_1434.LUT_INIT = 16'ha088;
    SB_LUT4 mux_24_i9_3_lut (.I0(\PID_CONTROLLER.result [8]), .I1(n63[8]), 
            .I2(n421), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_14_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1435 (.I0(Kd_delay_counter[5]), .I1(Kd_delay_counter[3]), 
            .I2(Kd_delay_counter[6]), .I3(Kd_delay_counter[4]), .O(n12_adj_3922));   // verilog/motorControl.v(49[10:29])
    defparam i5_4_lut_adj_1435.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1436 (.I0(Kd_delay_counter[1]), .I1(n12_adj_3922), 
            .I2(Kd_delay_counter[2]), .I3(Kd_delay_counter[0]), .O(n44626));   // verilog/motorControl.v(49[10:29])
    defparam i6_4_lut_adj_1436.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_24_i10_3_lut (.I0(\PID_CONTROLLER.result [9]), .I1(n63[9]), 
            .I2(n421), .I3(GND_net), .O(n462));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i11_3_lut (.I0(\PID_CONTROLLER.result [10]), .I1(n63[10]), 
            .I2(n421), .I3(GND_net), .O(n461));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i282_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n419_adj_3750));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i12_3_lut (.I0(\PID_CONTROLLER.result [11]), .I1(n63[10]), 
            .I2(n421), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n516_adj_3749));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_24_i13_3_lut (.I0(\PID_CONTROLLER.result [12]), .I1(n63[10]), 
            .I2(n421), .I3(GND_net), .O(n459));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_70_inv_0_i23_1_lut (.I0(pwm[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n79[22]));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_24_i14_3_lut (.I0(\PID_CONTROLLER.result [13]), .I1(n63[10]), 
            .I2(n421), .I3(GND_net), .O(n458));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_70_inv_0_i24_1_lut (.I0(pwm[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(PHASES_5__N_3046));   // verilog/motorControl.v(77[38:44])
    defparam unary_minus_70_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_24_i15_3_lut (.I0(\PID_CONTROLLER.result [14]), .I1(n63[10]), 
            .I2(n421), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n613_adj_3745));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i1_1_lut (.I0(\PID_CONTROLLER.err[0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[0]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_24_i16_3_lut (.I0(\PID_CONTROLLER.result [15]), .I1(n63[10]), 
            .I2(n421), .I3(GND_net), .O(n456));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_24_i17_3_lut (.I0(\PID_CONTROLLER.result [16]), .I1(n63[10]), 
            .I2(n421), .I3(GND_net), .O(n455));   // verilog/motorControl.v(42[18] 44[12])
    defparam mux_24_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1437 (.I0(pwm_23__N_2948), .I1(n47227), .I2(\PWMLimit[9] ), 
            .I3(n387), .O(n42013));
    defparam i1_4_lut_adj_1437.LUT_INIT = 16'ha088;
    SB_LUT4 mult_10_i477_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n710_adj_3743));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i87_2_lut (.I0(\Kd[1] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n128_adj_3742));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i87_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i24_2_lut (.I0(\Kd[0] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3741));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i2_1_lut (.I0(\PID_CONTROLLER.err[1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[1]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i3_1_lut (.I0(\PID_CONTROLLER.err[2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[2]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_14_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i4_1_lut (.I0(\PID_CONTROLLER.err[3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[3]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i5_1_lut (.I0(\PID_CONTROLLER.err[4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[4]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i6_1_lut (.I0(\PID_CONTROLLER.err[5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[5]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i7_1_lut (.I0(\PID_CONTROLLER.err[6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[6]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i7_2_lut  (.I0(\deadband[3] ), 
            .I1(\PID_CONTROLLER.result [3]), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_3928));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i7_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 mult_12_i152_2_lut (.I0(\Kd[2] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n225_adj_3733));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i152_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i9_2_lut  (.I0(\deadband[4] ), 
            .I1(\PID_CONTROLLER.result [4]), .I2(GND_net), .I3(GND_net), 
            .O(n9_adj_3929));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i9_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i17_2_lut  (.I0(\deadband[8] ), 
            .I1(\PID_CONTROLLER.result [8]), .I2(GND_net), .I3(GND_net), 
            .O(n17_adj_3930));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i17_2_lut .LUT_INIT = 16'h6666;
    SB_LUT4 i32911_4_lut (.I0(\deadband[9] ), .I1(n17_adj_3930), .I2(\PID_CONTROLLER.result [9]), 
            .I3(n9_adj_3929), .O(n48413));
    defparam i32911_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_12_i217_2_lut (.I0(\Kd[3] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n322));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i217_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32907_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(n48413), .O(n48409));
    defparam i32907_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 sub_11_inv_0_i8_1_lut (.I0(\PID_CONTROLLER.err[7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[7]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i282_2_lut (.I0(\Kd[4] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n419_adj_3731));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i282_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i9_1_lut (.I0(\PID_CONTROLLER.err[8] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[8]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i10_1_lut (.I0(\PID_CONTROLLER.err[9] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[9]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32921_3_lut (.I0(n15_adj_17), .I1(n13_adj_18), .I2(n11_adj_19), 
            .I3(GND_net), .O(n48423));
    defparam i32921_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_11_inv_0_i11_1_lut (.I0(\PID_CONTROLLER.err[10] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[10]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32889_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [13]), 
            .I2(\PID_CONTROLLER.result [14]), .I3(n48423), .O(n48391));
    defparam i32889_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 sub_11_inv_0_i12_1_lut (.I0(\PID_CONTROLLER.err[11] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[11]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i347_2_lut (.I0(\Kd[5] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n516));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32873_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(\deadband[9] ), .I3(n15_adj_17), .O(n48375));
    defparam i32873_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 mult_12_i412_2_lut (.I0(\Kd[6] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n613));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i477_2_lut (.I0(\Kd[7] ), .I1(n61[10]), .I2(GND_net), 
            .I3(GND_net), .O(n710));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i477_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_11_inv_0_i13_1_lut (.I0(\PID_CONTROLLER.err[12] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[12]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i30_4_lut  (.I0(\PID_CONTROLLER.result[7] ), 
            .I1(\PID_CONTROLLER.result [17]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [16]), 
            .O(n30_adj_3934));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i30_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 sub_11_inv_0_i14_1_lut (.I0(\PID_CONTROLLER.err[13] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[13]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i15_1_lut (.I0(\PID_CONTROLLER.err[14] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[14]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i16_1_lut (.I0(\PID_CONTROLLER.err[15] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[15]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32929_4_lut (.I0(n9_adj_3929), .I1(n7_adj_3928), .I2(\deadband[2] ), 
            .I3(\PID_CONTROLLER.result [2]), .O(n48431));
    defparam i32929_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 i33163_4_lut (.I0(n15_adj_17), .I1(n13_adj_18), .I2(n11_adj_19), 
            .I3(n48431), .O(n48665));
    defparam i33163_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32915_4_lut (.I0(\deadband[9] ), .I1(n17_adj_3930), .I2(\PID_CONTROLLER.result [9]), 
            .I3(n48665), .O(n48417));
    defparam i32915_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i33401_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\PID_CONTROLLER.result [11]), .I3(n48417), .O(n48903));
    defparam i33401_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32306_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\PID_CONTROLLER.result [13]), .I3(n48903), .O(n47808));
    defparam i32306_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i33149_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [14]), 
            .I2(\PID_CONTROLLER.result [15]), .I3(n47808), .O(n48651));
    defparam i33149_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33561_4_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\PID_CONTROLLER.result [16]), 
            .I2(\deadband[9] ), .I3(n48651), .O(n49063));
    defparam i33561_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33705_4_lut (.I0(\PID_CONTROLLER.result [19]), .I1(\PID_CONTROLLER.result [18]), 
            .I2(\deadband[9] ), .I3(n49063), .O(n49207));
    defparam i33705_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33233_3_lut (.I0(n6_adj_3935), .I1(\PID_CONTROLLER.result [10]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n48735));   // verilog/motorControl.v(37[10:27])
    defparam i33233_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32845_4_lut (.I0(\PID_CONTROLLER.result [22]), .I1(\PID_CONTROLLER.result [21]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [9]), .O(n48347));
    defparam i32845_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i24_4_lut  (.I0(\PID_CONTROLLER.result [9]), 
            .I1(\PID_CONTROLLER.result [22]), .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [21]), 
            .O(n24_adj_3936));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i24_4_lut .LUT_INIT = 16'h8f0e;
    SB_LUT4 i32255_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\deadband[9] ), .I3(n48409), .O(n47757));
    defparam i32255_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i17_rep_193_2_lut (.I0(\PID_CONTROLLER.result [22]), .I1(\deadband[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n50294));   // verilog/TinyFPGA_B.v(76[22:30])
    defparam i17_rep_193_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33495_3_lut (.I0(n24_adj_3936), .I1(n8_adj_3937), .I2(n48347), 
            .I3(GND_net), .O(n48997));   // verilog/motorControl.v(37[10:27])
    defparam i33495_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32641_4_lut (.I0(n48735), .I1(\PID_CONTROLLER.result [12]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [11]), .O(n48143));   // verilog/motorControl.v(37[10:27])
    defparam i32641_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i4_4_lut  (.I0(\deadband[0] ), 
            .I1(\PID_CONTROLLER.result [1]), .I2(\deadband[1] ), .I3(\PID_CONTROLLER.result [0]), 
            .O(n4_adj_3938));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i4_4_lut .LUT_INIT = 16'h4d0c;
    SB_LUT4 i33229_3_lut (.I0(n4_adj_3938), .I1(\PID_CONTROLLER.result [13]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n48731));   // verilog/motorControl.v(37[10:27])
    defparam i33229_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32285_4_lut (.I0(\deadband[9] ), .I1(\PID_CONTROLLER.result [15]), 
            .I2(\PID_CONTROLLER.result [16]), .I3(n48391), .O(n47787));
    defparam i32285_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i19_rep_171_2_lut (.I0(\PID_CONTROLLER.result [17]), .I1(\deadband[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n50272));   // verilog/TinyFPGA_B.v(76[22:30])
    defparam i19_rep_171_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33603_3_lut (.I0(n30_adj_3934), .I1(n10_adj_3939), .I2(n48375), 
            .I3(GND_net), .O(n49105));   // verilog/motorControl.v(37[10:27])
    defparam i33603_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 sub_11_inv_0_i17_1_lut (.I0(\PID_CONTROLLER.err[16] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[16]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i18_1_lut (.I0(\PID_CONTROLLER.err[17] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[17]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i19_1_lut (.I0(\PID_CONTROLLER.err[18] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[18]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_11_inv_0_i20_1_lut (.I0(\PID_CONTROLLER.err[19] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[19]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32643_4_lut (.I0(n48731), .I1(\PID_CONTROLLER.result [15]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [14]), .O(n48145));   // verilog/motorControl.v(37[10:27])
    defparam i32643_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 sub_11_inv_0_i21_1_lut (.I0(\PID_CONTROLLER.err[20] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[20]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33725_4_lut (.I0(n48145), .I1(n49105), .I2(n50272), .I3(n47787), 
            .O(n49227));   // verilog/motorControl.v(37[10:27])
    defparam i33725_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 sub_11_inv_0_i22_1_lut (.I0(\PID_CONTROLLER.err[21] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[21]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33726_3_lut (.I0(n49227), .I1(\PID_CONTROLLER.result [18]), 
            .I2(\deadband[9] ), .I3(GND_net), .O(n49228));   // verilog/motorControl.v(37[10:27])
    defparam i33726_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[10] ), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3711));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32259_4_lut (.I0(\PID_CONTROLLER.result [21]), .I1(\PID_CONTROLLER.result [20]), 
            .I2(\deadband[9] ), .I3(n49207), .O(n47761));
    defparam i32259_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i33678_4_lut (.I0(n48143), .I1(n48997), .I2(n50294), .I3(n47757), 
            .O(n49180));   // verilog/motorControl.v(37[10:27])
    defparam i33678_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32649_4_lut (.I0(n49228), .I1(\PID_CONTROLLER.result [20]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [19]), .O(n48151));   // verilog/motorControl.v(37[10:27])
    defparam i32649_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 sub_11_inv_0_i23_1_lut (.I0(\PID_CONTROLLER.err[22] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[22]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33721_4_lut (.I0(n48151), .I1(n49180), .I2(n50294), .I3(n47761), 
            .O(n49223));   // verilog/motorControl.v(37[10:27])
    defparam i33721_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 sub_11_inv_0_i24_1_lut (.I0(\PID_CONTROLLER.err[23] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[23]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i150_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n222_adj_3706));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i33683_4_lut (.I0(n49223), .I1(\PID_CONTROLLER.result [24]), 
            .I2(\deadband[9] ), .I3(\PID_CONTROLLER.result [23]), .O(n50));   // verilog/motorControl.v(37[10:27])
    defparam i33683_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 sub_11_inv_0_i32_1_lut (.I0(\PID_CONTROLLER.err[31] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n76[26]));   // verilog/motorControl.v(36[31:45])
    defparam sub_11_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i215_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n319));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i215_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i280_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n416_adj_3704));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i280_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n513));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n610_adj_3703));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i89_2_lut (.I0(\Kd[1] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_3702));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i26_2_lut (.I0(\Kd[0] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_3701));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i154_2_lut (.I0(\Kd[2] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n228_adj_3700));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i154_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i475_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n707));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i219_2_lut (.I0(\Kd[3] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n325));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i219_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i284_2_lut (.I0(\Kd[4] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n422));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i284_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i349_2_lut (.I0(\Kd[5] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n519_adj_3699));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i414_2_lut (.I0(\Kd[6] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n616));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i479_2_lut (.I0(\Kd[7] ), .I1(n61[11]), .I2(GND_net), 
            .I3(GND_net), .O(n713));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i479_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3698));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i107_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n158_adj_3697));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i107_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i44_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[21] ), 
            .I2(GND_net), .I3(GND_net), .O(n65_adj_3696));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i44_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i172_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n255_adj_3695));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i172_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_3694));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i237_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n352_adj_3692));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i237_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_3691));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n449_adj_3689));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_3688));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n546_adj_3686));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i432_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n643_adj_3685));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i497_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[20] ), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_3684));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i497_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i91_2_lut (.I0(\Kd[1] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n134_adj_3682));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i91_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i28_2_lut (.I0(\Kd[0] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3681));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[0]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22993_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(GND_net), .O(n16640[0]));   // verilog/motorControl.v(36[17:23])
    defparam i22993_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i23193_2_lut_3_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\Kp[2] ), 
            .I3(GND_net), .O(n38898));   // verilog/motorControl.v(36[17:23])
    defparam i23193_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i32167_3_lut_3_lut (.I0(n63[10]), .I1(n421), .I2(\PID_CONTROLLER.result [17]), 
            .I3(GND_net), .O(n47225));   // verilog/motorControl.v(40[28:37])
    defparam i32167_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 i32404_3_lut_3_lut (.I0(n63[10]), .I1(n421), .I2(\PID_CONTROLLER.result [18]), 
            .I3(GND_net), .O(n47227));   // verilog/motorControl.v(40[28:37])
    defparam i32404_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[1]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[2]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[9] ), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3677));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[3]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32094_3_lut_3_lut (.I0(n63[10]), .I1(n421), .I2(\PID_CONTROLLER.result [19]), 
            .I3(GND_net), .O(n47180));   // verilog/motorControl.v(40[28:37])
    defparam i32094_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 mult_14_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[4]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i156_2_lut (.I0(\Kd[2] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n231_adj_3674));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i148_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n219_adj_3673));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[5]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i213_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n316_adj_3671));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i213_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[6]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i221_2_lut (.I0(\Kd[3] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n328_adj_3669));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i221_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32231_3_lut_3_lut (.I0(n63[10]), .I1(n421), .I2(\PID_CONTROLLER.result [20]), 
            .I3(GND_net), .O(n47182));   // verilog/motorControl.v(40[28:37])
    defparam i32231_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 i32229_3_lut_3_lut (.I0(n63[10]), .I1(n421), .I2(\PID_CONTROLLER.result [23]), 
            .I3(GND_net), .O(n47188));   // verilog/motorControl.v(40[28:37])
    defparam i32229_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 i32234_3_lut_3_lut (.I0(n63[10]), .I1(n421), .I2(\PID_CONTROLLER.result [22]), 
            .I3(GND_net), .O(n47186));   // verilog/motorControl.v(40[28:37])
    defparam i32234_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 LessThan_20_i6_3_lut_3_lut (.I0(\PWMLimit[3] ), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(38[12:27])
    defparam LessThan_20_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[7]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i278_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n413_adj_3666));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[8]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i286_2_lut (.I0(\Kd[4] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n425_adj_3664));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i286_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i343_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n510_adj_3663));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[9]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[10]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n607_adj_3660));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[11]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i473_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err[8] ), 
            .I2(GND_net), .I3(GND_net), .O(n704));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i473_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i351_2_lut (.I0(\Kd[5] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n522_adj_3658));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[12]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[13]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i416_2_lut (.I0(\Kd[6] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n619_adj_3655));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i481_2_lut (.I0(\Kd[7] ), .I1(n61[12]), .I2(GND_net), 
            .I3(GND_net), .O(n716));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i481_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[14]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[15]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[16]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[17]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[18]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[19]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[20]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[21]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31834_2_lut_3_lut_4_lut (.I0(n19600), .I1(hall2), .I2(n19608), 
            .I3(n878), .O(n47192));   // verilog/motorControl.v(77[14] 98[8])
    defparam i31834_2_lut_3_lut_4_lut.LUT_INIT = 16'h7500;
    SB_LUT4 LessThan_4_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3940));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i4_2_lut_adj_1438 (.I0(n19_adj_3381), .I1(n25), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_3941));   // verilog/motorControl.v(33[38:63])
    defparam i4_2_lut_adj_1438.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1439 (.I0(n33), .I1(n43_adj_3845), .I2(n27), 
            .I3(n35_adj_3853), .O(n24_adj_3942));   // verilog/motorControl.v(33[38:63])
    defparam i10_4_lut_adj_1439.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1440 (.I0(n41_adj_3847), .I1(n45_adj_3843), .I2(n31), 
            .I3(n23_c), .O(n22_adj_3943));   // verilog/motorControl.v(33[38:63])
    defparam i8_4_lut_adj_1440.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1441 (.I0(n29_c), .I1(n24_adj_3942), .I2(n18_adj_3941), 
            .I3(n37_adj_3851), .O(n26_adj_3944));   // verilog/motorControl.v(33[38:63])
    defparam i12_4_lut_adj_1441.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1442 (.I0(n21_c), .I1(n26_adj_3944), .I2(n22_adj_3943), 
            .I3(n39_adj_3849), .O(n45037));   // verilog/motorControl.v(33[38:63])
    defparam i13_4_lut_adj_1442.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_4_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), .I1(IntegralLimit[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3945));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(IntegralLimit[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_3946));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), .I1(IntegralLimit[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3947));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32963_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3947), 
            .I2(IntegralLimit[9]), .I3(n9_adj_3946), .O(n48465));
    defparam i32963_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32961_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[10]), 
            .I2(IntegralLimit[11]), .I3(n48465), .O(n48463));
    defparam i32961_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i32354_4_lut (.I0(n11_adj_3495), .I1(n9_adj_3497), .I2(n7_adj_3500), 
            .I3(n5_adj_3502), .O(n47856));
    defparam i32354_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_4_i13_rep_366_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n50467));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i13_rep_366_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32967_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n50467), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3945), .O(n48469));
    defparam i32967_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32955_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n48469), .O(n48457));
    defparam i32955_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i32368_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n47870));
    defparam i32368_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 LessThan_4_i35_rep_354_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n50455));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i35_rep_354_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_4_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3948));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_4_i30_4_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[16]), .O(n30_adj_3949));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i30_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_4_i5_2_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(IntegralLimit[2]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3950));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32971_4_lut (.I0(n9_adj_3946), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n5_adj_3950), .I3(IntegralLimit[3]), .O(n48473));
    defparam i32971_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i32969_4_lut (.I0(\PID_CONTROLLER.integral [6]), .I1(n11_adj_3945), 
            .I2(IntegralLimit[6]), .I3(n48473), .O(n48471));
    defparam i32969_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i32384_4_lut (.I0(n17_adj_3947), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n48471), .I3(IntegralLimit[7]), .O(n47886));
    defparam i32384_4_lut.LUT_INIT = 16'haeab;
    SB_LUT4 i33183_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[9]), 
            .I2(IntegralLimit[10]), .I3(n47886), .O(n48685));
    defparam i33183_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33575_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[11]), 
            .I2(IntegralLimit[12]), .I3(n48685), .O(n49077));
    defparam i33575_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i32957_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[13]), 
            .I2(IntegralLimit[14]), .I3(n49077), .O(n48459));
    defparam i32957_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i33407_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n48459), .O(n48909));
    defparam i33407_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33644_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[17]), 
            .I2(IntegralLimit[18]), .I3(n48909), .O(n49146));
    defparam i33644_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 i33743_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[19]), 
            .I2(IntegralLimit[20]), .I3(n49146), .O(n49245));
    defparam i33743_4_lut.LUT_INIT = 16'hff7e;
    SB_LUT4 LessThan_4_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3951));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32453_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(IntegralLimit[9]), .O(n47955));
    defparam i32453_4_lut.LUT_INIT = 16'h7ffe;
    SB_LUT4 LessThan_4_i24_4_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(IntegralLimit[21]), .O(n24_adj_3952));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i24_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33241_3_lut (.I0(n6_adj_3951), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48743));   // verilog/motorControl.v(33[10:34])
    defparam i33241_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32360_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[12]), 
            .I2(IntegralLimit[21]), .I3(n48463), .O(n47862));
    defparam i32360_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 LessThan_4_i45_rep_319_2_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n50420));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i45_rep_319_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i33259_3_lut (.I0(n24_adj_3952), .I1(n8_adj_3940), .I2(n47955), 
            .I3(GND_net), .O(n48761));   // verilog/motorControl.v(33[10:34])
    defparam i33259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32629_4_lut (.I0(n48743), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[11]), .O(n48131));   // verilog/motorControl.v(33[10:34])
    defparam i32629_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 LessThan_6_i4_4_lut (.I0(n67[0]), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3), .I3(\PID_CONTROLLER.integral [0]), .O(n4_adj_3953));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i4_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i33235_3_lut (.I0(n4_adj_3953), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n11_adj_3495), .I3(GND_net), .O(n48737));   // verilog/motorControl.v(33[38:63])
    defparam i33235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33236_3_lut (.I0(n48737), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n13_adj_3492), .I3(GND_net), .O(n48738));   // verilog/motorControl.v(33[38:63])
    defparam i33236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i8_3_lut (.I0(\PID_CONTROLLER.integral [4]), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n17_adj_3472), .I3(GND_net), .O(n8_adj_3954));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32348_2_lut (.I0(n17_adj_3472), .I1(n9_adj_3497), .I2(GND_net), 
            .I3(GND_net), .O(n47850));
    defparam i32348_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_6_i6_3_lut (.I0(\PID_CONTROLLER.integral [2]), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n7_adj_3500), .I3(GND_net), .O(n6_adj_3955));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_6_i16_3_lut (.I0(n8_adj_3954), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n45037), .I3(GND_net), .O(n16_adj_3956));   // verilog/motorControl.v(33[38:63])
    defparam LessThan_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32350_4_lut (.I0(n17_adj_3472), .I1(n15_adj_3488), .I2(n13_adj_3492), 
            .I3(n47856), .O(n47852));
    defparam i32350_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i33369_4_lut (.I0(n16_adj_3956), .I1(n6_adj_3955), .I2(n45037), 
            .I3(n47850), .O(n48871));   // verilog/motorControl.v(33[38:63])
    defparam i33369_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32639_3_lut (.I0(n48738), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n15_adj_3488), .I3(GND_net), .O(n48141));   // verilog/motorControl.v(33[38:63])
    defparam i32639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33625_4_lut (.I0(n48141), .I1(n48871), .I2(n45037), .I3(n47852), 
            .O(n49127));   // verilog/motorControl.v(33[38:63])
    defparam i33625_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 LessThan_4_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(IntegralLimit[1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), .O(n4_adj_3957));   // verilog/motorControl.v(33[10:34])
    defparam LessThan_4_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i33239_3_lut (.I0(n4_adj_3957), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n48741));   // verilog/motorControl.v(33[10:34])
    defparam i33239_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32370_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[15]), 
            .I2(IntegralLimit[16]), .I3(n48457), .O(n47872));
    defparam i32370_4_lut.LUT_INIT = 16'h5adb;
    SB_LUT4 i33601_4_lut (.I0(n30_adj_3949), .I1(n10_adj_3948), .I2(n50455), 
            .I3(n47870), .O(n49103));   // verilog/motorControl.v(33[10:34])
    defparam i33601_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32631_4_lut (.I0(n48741), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[14]), .O(n48133));   // verilog/motorControl.v(33[10:34])
    defparam i32631_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33723_4_lut (.I0(n48133), .I1(n49103), .I2(n50455), .I3(n47872), 
            .O(n49225));   // verilog/motorControl.v(33[10:34])
    defparam i33723_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33724_3_lut (.I0(n49225), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n49226));   // verilog/motorControl.v(33[10:34])
    defparam i33724_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32943_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(IntegralLimit[21]), 
            .I2(IntegralLimit[22]), .I3(n49245), .O(n48445));
    defparam i32943_4_lut.LUT_INIT = 16'h7eff;
    SB_LUT4 i33509_4_lut (.I0(n48131), .I1(n48761), .I2(n50420), .I3(n47862), 
            .O(n49011));   // verilog/motorControl.v(33[10:34])
    defparam i33509_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32637_4_lut (.I0(n49226), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[19]), .O(n48139));   // verilog/motorControl.v(33[10:34])
    defparam i32637_4_lut.LUT_INIT = 16'h8f0e;
    SB_LUT4 i33626_3_lut (.I0(n49127), .I1(n67[23]), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(GND_net), .O(n49128));   // verilog/motorControl.v(33[38:63])
    defparam i33626_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i33623_3_lut (.I0(n48139), .I1(n49011), .I2(n48445), .I3(GND_net), 
            .O(n49125));   // verilog/motorControl.v(33[10:34])
    defparam i33623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_1443 (.I0(n49125), .I1(n49128), .I2(\PID_CONTROLLER.integral [9]), 
            .I3(IntegralLimit[23]), .O(n55_adj_3646));   // verilog/motorControl.v(33[10:63])
    defparam i8_4_lut_adj_1443.LUT_INIT = 16'h80c8;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[22]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32225_3_lut_3_lut (.I0(n63[10]), .I1(n421), .I2(\PID_CONTROLLER.result [21]), 
            .I3(GND_net), .O(n47184));   // verilog/motorControl.v(40[28:37])
    defparam i32225_3_lut_3_lut.LUT_INIT = 16'hb8b8;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n75[23]));   // verilog/motorControl.v(32[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_12_i93_2_lut (.I0(\Kd[1] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n137_adj_3643));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i93_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i30_2_lut (.I0(\Kd[0] ), .I1(n61[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_3642));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i158_2_lut (.I0(\Kd[2] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n234_adj_3641));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i158_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i223_2_lut (.I0(\Kd[3] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n331_adj_3640));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i223_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i49_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n72));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i49_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_12_i288_2_lut (.I0(\Kd[4] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n428_adj_3639));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i288_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i98_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n145_adj_3638));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i98_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_12_i353_2_lut (.I0(\Kd[5] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n525_adj_3637));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i147_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n218_adj_3636));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i147_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i32190_3_lut_4_lut (.I0(\PWMLimit[3] ), .I1(\PID_CONTROLLER.result [3]), 
            .I2(\PID_CONTROLLER.result [2]), .I3(\PWMLimit[2] ), .O(n47692));   // verilog/motorControl.v(38[12:27])
    defparam i32190_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_12_i418_2_lut (.I0(\Kd[6] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n622_adj_3635));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3634));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[4] ), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3633));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [4]), 
            .I1(\PID_CONTROLLER.result [8]), .I2(\deadband[8] ), .I3(GND_net), 
            .O(n8_adj_3937));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i8_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut  (.I0(\PID_CONTROLLER.result [2]), 
            .I1(\PID_CONTROLLER.result [3]), .I2(\deadband[3] ), .I3(GND_net), 
            .O(n6_adj_3935));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i6_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut  (.I0(\PID_CONTROLLER.result[5] ), 
            .I1(\PID_CONTROLLER.result[6] ), .I2(\deadband[6] ), .I3(GND_net), 
            .O(n10_adj_3939));   // verilog/motorControl.v(37[10:27])
    defparam \PID_CONTROLLER.result_31__I_0_i10_3_lut_3_lut .LUT_INIT = 16'h8e8e;
    SB_LUT4 i6309_2_lut_3_lut (.I0(hall3), .I1(hall1), .I2(n878), .I3(GND_net), 
            .O(n19615));   // verilog/motorControl.v(96[14] 98[8])
    defparam i6309_2_lut_3_lut.LUT_INIT = 16'h2f2f;
    SB_LUT4 i28515_2_lut_3_lut (.I0(hall3), .I1(hall2), .I2(hall1), .I3(GND_net), 
            .O(n44011));
    defparam i28515_2_lut_3_lut.LUT_INIT = 16'h7474;
    SB_LUT4 i10239_2_lut_3_lut (.I0(n19600), .I1(hall2), .I2(n19608), 
            .I3(GND_net), .O(PHASES_5__N_3039[2]));   // verilog/motorControl.v(74[7] 76[10])
    defparam i10239_2_lut_3_lut.LUT_INIT = 16'h7575;
    SB_LUT4 i28584_2_lut_4_lut (.I0(hall3), .I1(hall1), .I2(n19292), .I3(n880), 
            .O(n44081));
    defparam i28584_2_lut_4_lut.LUT_INIT = 16'hfff2;
    SB_LUT4 i32406_2_lut_4_lut (.I0(n911), .I1(hall3), .I2(hall1), .I3(n878), 
            .O(n47229));
    defparam i32406_2_lut_4_lut.LUT_INIT = 16'h4500;
    SB_LUT4 mult_12_i483_2_lut (.I0(\Kd[7] ), .I1(n61[13]), .I2(GND_net), 
            .I3(GND_net), .O(n719_adj_3632));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i483_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23323_3_lut_4_lut (.I0(n10114[2]), .I1(\Kd[4] ), .I2(n61[25]), 
            .I3(n6_adj_3958), .O(n8_adj_3918));   // verilog/motorControl.v(36[26:45])
    defparam i23323_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i2_3_lut_4_lut_adj_1444 (.I0(\Kd[5] ), .I1(n61[25]), .I2(\Kd[4] ), 
            .I3(n6_adj_3958), .O(n8_adj_3919));   // verilog/motorControl.v(36[26:45])
    defparam i2_3_lut_4_lut_adj_1444.LUT_INIT = 16'hb748;
    SB_LUT4 i23315_3_lut_4_lut (.I0(n11529[1]), .I1(\Kd[3] ), .I2(n61[25]), 
            .I3(n4_adj_3910), .O(n6_adj_3958));   // verilog/motorControl.v(36[26:45])
    defparam i23315_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i23294_2_lut_3_lut (.I0(\Kd[0] ), .I1(n61[25]), .I2(\Kd[1] ), 
            .I3(GND_net), .O(n36732));   // verilog/motorControl.v(36[26:45])
    defparam i23294_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i32402_2_lut_3_lut (.I0(hall3), .I1(hall2), .I2(n878), .I3(GND_net), 
            .O(n47234));
    defparam i32402_2_lut_3_lut.LUT_INIT = 16'hb0b0;
    SB_LUT4 i2_3_lut_4_lut_adj_1445 (.I0(hall1), .I1(n19292), .I2(hall2), 
            .I3(n19608), .O(n44840));
    defparam i2_3_lut_4_lut_adj_1445.LUT_INIT = 16'hdfda;
    SB_LUT4 i1_3_lut_4_lut_adj_1446 (.I0(n10114[2]), .I1(\Kd[4] ), .I2(n61[25]), 
            .I3(n6_adj_3958), .O(n10114[3]));   // verilog/motorControl.v(36[26:45])
    defparam i1_3_lut_4_lut_adj_1446.LUT_INIT = 16'h956a;
    SB_LUT4 i3660_2_lut_3_lut (.I0(hall1), .I1(hall2), .I2(n19608), .I3(GND_net), 
            .O(n16801));   // verilog/motorControl.v(74[7] 76[10])
    defparam i3660_2_lut_3_lut.LUT_INIT = 16'h7474;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\Kd[3] ), .I1(n61[25]), .I2(n4_adj_3910), 
            .I3(n11529[1]), .O(n10114[2]));   // verilog/motorControl.v(36[26:45])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1447 (.I0(hall1), .I1(hall2), .I2(n878), 
            .I3(n19608), .O(n20352));   // verilog/motorControl.v(96[14] 98[8])
    defparam i2_3_lut_4_lut_adj_1447.LUT_INIT = 16'h7f4f;
    SB_LUT4 mult_14_i196_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n291));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i196_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_14_i245_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n364_adj_3630));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i245_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_2_lut_3_lut (.I0(hall1), .I1(hall2), .I2(hall3), .I3(GND_net), 
            .O(n6_adj_3917));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i14976_3_lut_4_lut (.I0(n880), .I1(hall3), .I2(hall1), .I3(hall2), 
            .O(PHASES_5__N_3039[1]));   // verilog/motorControl.v(74[7] 76[10])
    defparam i14976_3_lut_4_lut.LUT_INIT = 16'h0c2e;
    SB_LUT4 i1_4_lut_4_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n6_adj_3904), .I3(n38898), .O(n7_adj_3906));   // verilog/motorControl.v(36[17:23])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h78b4;
    SB_LUT4 i23175_3_lut_4_lut (.I0(n16653[1]), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n4_adj_3959), .O(n6_adj_3904));   // verilog/motorControl.v(36[17:23])
    defparam i23175_3_lut_4_lut.LUT_INIT = 16'hea80;
    SB_LUT4 i23386_2_lut_3_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(\Kp[1] ), .I3(GND_net), .O(n36452));   // verilog/motorControl.v(36[17:23])
    defparam i23386_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut (.I0(n16653[1]), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err[31] ), 
            .I3(n4_adj_3959), .O(n16647[2]));   // verilog/motorControl.v(36[17:23])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h956a;
    SB_LUT4 i1_2_lut_3_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n4_adj_3959), .I3(GND_net), .O(n43578));   // verilog/motorControl.v(36[17:23])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i23199_4_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[31] ), 
            .I2(n16640[0]), .I3(n36452), .O(n4_adj_3959));   // verilog/motorControl.v(36[17:23])
    defparam i23199_4_lut_4_lut.LUT_INIT = 16'hf8a0;
    SB_LUT4 mult_14_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3629));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i294_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n437_adj_3628));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i294_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_3627));   // verilog/motorControl.v(36[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_12_i337_2_lut (.I0(\Kd[5] ), .I1(n61[5]), .I2(GND_net), 
            .I3(GND_net), .O(n501));   // verilog/motorControl.v(36[26:45])
    defparam mult_12_i337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22995_3_lut_4_lut_4_lut_4_lut (.I0(\PID_CONTROLLER.err[31] ), 
            .I1(\Kp[0] ), .I2(\Kp[1] ), .I3(\Kp[2] ), .O(n16653[1]));   // verilog/motorControl.v(36[17:23])
    defparam i22995_3_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'h02a8;
    SB_LUT4 mult_14_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_3626));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_14_i343_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n510));   // verilog/motorControl.v(36[48:59])
    defparam mult_14_i343_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i32206_2_lut_4_lut (.I0(\PID_CONTROLLER.result [8]), .I1(pwm_23__N_2951[8]), 
            .I2(\PID_CONTROLLER.result [4]), .I3(pwm_23__N_2951[4]), .O(n47708));
    defparam i32206_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_2_lut_4_lut_adj_1448 (.I0(\PID_CONTROLLER.result [28]), .I1(\PID_CONTROLLER.result [30]), 
            .I2(\PID_CONTROLLER.result [29]), .I3(n56_adj_3392), .O(n43147));   // verilog/motorControl.v(38[12:27])
    defparam i1_2_lut_4_lut_adj_1448.LUT_INIT = 16'h8000;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=47, LSE_LCOL=12, LSE_RCOL=39, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[12] 38[39])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n24341, encoder1_position, clk32MHz, 
            n24340, n24339, n24353, n24352, n24351, n24350, n24349, 
            n24348, n24347, n24346, n24345, n24344, n24343, n24342, 
            n24338, n24337, data_o, n24336, n24335, n24334, n24333, 
            n24332, n2241, GND_net, n24321, n23746, count_enable, 
            n24385, n44576, reg_B, PIN_18_c_1, PIN_19_c_0, n23752) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n24341;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n24340;
    input n24339;
    input n24353;
    input n24352;
    input n24351;
    input n24350;
    input n24349;
    input n24348;
    input n24347;
    input n24346;
    input n24345;
    input n24344;
    input n24343;
    input n24342;
    input n24338;
    input n24337;
    output [1:0]data_o;
    input n24336;
    input n24335;
    input n24334;
    input n24333;
    input n24332;
    output [23:0]n2241;
    input GND_net;
    input n24321;
    input n23746;
    output count_enable;
    input n24385;
    output n44576;
    output [1:0]reg_B;
    input PIN_18_c_1;
    input PIN_19_c_0;
    input n23752;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire B_delayed, A_delayed, n2233, n37121, n37120, n37119, n37118, 
        n37117, n37116, n37115, n37114, n37113, n37112, n37111, 
        n37110, n37109, n37108, n37107, n37106, n37105, n37104, 
        n37103, n37102, n37101, n37100, n37099, count_direction, 
        n37098;
    
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n24341));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n24340));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n24339));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n24353));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n24352));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n24351));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n24350));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n24349));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n24348));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n24347));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n24346));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n24345));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n24344));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n24343));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n24342));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n24338));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n24337));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n24336));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n24335));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n24334));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n24333));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n24332));   // quad.v(35[10] 41[6])
    SB_LUT4 add_523_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2233), 
            .I3(n37121), .O(n2241[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_523_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2233), 
            .I3(n37120), .O(n2241[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_24 (.CI(n37120), .I0(encoder1_position[22]), .I1(n2233), 
            .CO(n37121));
    SB_LUT4 add_523_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2233), 
            .I3(n37119), .O(n2241[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_23 (.CI(n37119), .I0(encoder1_position[21]), .I1(n2233), 
            .CO(n37120));
    SB_LUT4 add_523_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2233), 
            .I3(n37118), .O(n2241[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_22 (.CI(n37118), .I0(encoder1_position[20]), .I1(n2233), 
            .CO(n37119));
    SB_LUT4 add_523_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2233), 
            .I3(n37117), .O(n2241[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_21 (.CI(n37117), .I0(encoder1_position[19]), .I1(n2233), 
            .CO(n37118));
    SB_LUT4 add_523_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2233), 
            .I3(n37116), .O(n2241[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_20 (.CI(n37116), .I0(encoder1_position[18]), .I1(n2233), 
            .CO(n37117));
    SB_LUT4 add_523_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2233), 
            .I3(n37115), .O(n2241[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_19 (.CI(n37115), .I0(encoder1_position[17]), .I1(n2233), 
            .CO(n37116));
    SB_LUT4 add_523_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2233), 
            .I3(n37114), .O(n2241[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_18 (.CI(n37114), .I0(encoder1_position[16]), .I1(n2233), 
            .CO(n37115));
    SB_LUT4 add_523_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2233), 
            .I3(n37113), .O(n2241[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_17 (.CI(n37113), .I0(encoder1_position[15]), .I1(n2233), 
            .CO(n37114));
    SB_LUT4 add_523_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2233), 
            .I3(n37112), .O(n2241[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_16 (.CI(n37112), .I0(encoder1_position[14]), .I1(n2233), 
            .CO(n37113));
    SB_LUT4 add_523_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2233), 
            .I3(n37111), .O(n2241[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_15 (.CI(n37111), .I0(encoder1_position[13]), .I1(n2233), 
            .CO(n37112));
    SB_LUT4 add_523_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2233), 
            .I3(n37110), .O(n2241[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_14 (.CI(n37110), .I0(encoder1_position[12]), .I1(n2233), 
            .CO(n37111));
    SB_LUT4 add_523_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2233), 
            .I3(n37109), .O(n2241[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_13 (.CI(n37109), .I0(encoder1_position[11]), .I1(n2233), 
            .CO(n37110));
    SB_LUT4 add_523_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2233), 
            .I3(n37108), .O(n2241[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_12 (.CI(n37108), .I0(encoder1_position[10]), .I1(n2233), 
            .CO(n37109));
    SB_LUT4 add_523_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2233), 
            .I3(n37107), .O(n2241[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_11 (.CI(n37107), .I0(encoder1_position[9]), .I1(n2233), 
            .CO(n37108));
    SB_LUT4 add_523_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2233), 
            .I3(n37106), .O(n2241[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_10 (.CI(n37106), .I0(encoder1_position[8]), .I1(n2233), 
            .CO(n37107));
    SB_LUT4 add_523_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2233), 
            .I3(n37105), .O(n2241[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_9 (.CI(n37105), .I0(encoder1_position[7]), .I1(n2233), 
            .CO(n37106));
    SB_LUT4 add_523_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2233), 
            .I3(n37104), .O(n2241[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_8 (.CI(n37104), .I0(encoder1_position[6]), .I1(n2233), 
            .CO(n37105));
    SB_LUT4 add_523_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2233), 
            .I3(n37103), .O(n2241[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_7 (.CI(n37103), .I0(encoder1_position[5]), .I1(n2233), 
            .CO(n37104));
    SB_LUT4 add_523_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2233), 
            .I3(n37102), .O(n2241[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_6 (.CI(n37102), .I0(encoder1_position[4]), .I1(n2233), 
            .CO(n37103));
    SB_LUT4 add_523_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2233), 
            .I3(n37101), .O(n2241[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_5 (.CI(n37101), .I0(encoder1_position[3]), .I1(n2233), 
            .CO(n37102));
    SB_LUT4 add_523_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2233), 
            .I3(n37100), .O(n2241[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_4 (.CI(n37100), .I0(encoder1_position[2]), .I1(n2233), 
            .CO(n37101));
    SB_LUT4 add_523_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2233), 
            .I3(n37099), .O(n2241[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_3 (.CI(n37099), .I0(encoder1_position[1]), .I1(n2233), 
            .CO(n37100));
    SB_LUT4 add_523_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n37098), .O(n2241[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_523_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_523_2 (.CI(n37098), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n37099));
    SB_CARRY add_523_1 (.CI(GND_net), .I0(n2233), .I1(n2233), .CO(n37098));
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n24321));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n23746));   // quad.v(35[10] 41[6])
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i719_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2233));   // quad.v(37[5] 40[8])
    defparam i719_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n24385(n24385), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .n44576(n44576), .GND_net(GND_net), .reg_B({reg_B}), .PIN_18_c_1(PIN_18_c_1), 
            .PIN_19_c_0(PIN_19_c_0), .n23752(n23752)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n24385, data_o, clk32MHz, n44576, GND_net, 
            reg_B, PIN_18_c_1, PIN_19_c_0, n23752) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n24385;
    output [1:0]data_o;
    input clk32MHz;
    output n44576;
    input GND_net;
    output [1:0]reg_B;
    input PIN_18_c_1;
    input PIN_19_c_0;
    input n23752;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    
    wire cnt_next_2__N_3104, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n24385));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n44576));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1050__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_18_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_19_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n23752));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1050__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1050__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i23371_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23371_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i23364_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23364_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n44576), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3104));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i23362_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i23362_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, \data_in_frame[13] , \data_in_frame[11] , GND_net, 
            gearBoxRatio, n10, n24253, \data_in[0] , n24252, n24251, 
            \data_in_frame[14] , \data_in_frame[19] , n24250, rx_data, 
            \deadband[9] , \deadband[8] , \deadband[7] , \deadband[6] , 
            \deadband[5] , \deadband[4] , \deadband[3] , \deadband[2] , 
            \deadband[1] , n24412, setpoint, n24411, n24410, n42279, 
            n24408, n24407, n24406, n24405, n24404, n24403, n24402, 
            n24401, n24400, n24399, n24398, n24397, n24396, n24395, 
            n24394, n24393, n24392, n24391, n24390, n24388, VCC_net, 
            byte_transmit_counter, n23822, n24236, \data_in[2] , n24234, 
            n24233, n24228, \data_in[3][2] , n24227, \data_in[3][3] , 
            n24226, \data_in[3][4] , n24225, \data_in[3][5] , n24223, 
            \data_in[3][7] , n24222, \data_out_frame[0][2] , n24221, 
            \data_out_frame[0][3] , n24220, \data_out_frame[0][4] , n24217, 
            \data_out_frame[5][2] , IntegralLimit, \Kp[1] , \Kp[2] , 
            n24249, n24248, rx_data_ready, n24245, \data_in[1][1] , 
            n24244, \data_in[1][2] , \Kp[3] , \Kp[4] , \FRAME_MATCHER.state , 
            n47, n3839, n29726, \Kp[5] , n43231, n43238, n43253, 
            \data_in_frame[1][4] , n24068, \data_in_frame[3] , n24067, 
            n24066, n24065, n24064, n24063, n24062, n24061, n24243, 
            \data_in[1][3] , \data_in_frame[5] , n24052, n24051, n24050, 
            n24049, n23533, n24048, n24047, n24046, n24045, \Kp[6] , 
            \Kp[7] , \Ki[1] , n24036, \data_in_frame[7] , n24035, 
            n24034, n24033, n24032, n24031, n24030, n24029, n24242, 
            \data_in[1][4] , n23825, \data_in_frame[10][6] , n24004, 
            n24003, n24002, n24001, n24000, n23999, n23998, n23997, 
            n23988, n23987, n23986, n23985, n23984, n23983, n23982, 
            n20342, n23981, \data_in_frame[14][0] , n24241, \data_in[1][5] , 
            n23972, \data_in_frame[15] , n23971, n23970, n23969, n23968, 
            n23967, n23966, n23965, n23838, n22456, n43255, \data_in_frame[16][1] , 
            n23835, n23832, n23823, n23820, n2241, \data_in_frame[18][0] , 
            \data_in_frame[18][2] , Kp_23__N_865, n43441, n23940, n23939, 
            n23938, n103, n23937, n23936, n23935, n23934, n23933, 
            Kp_23__N_515, n45225, n122, n44586, n23924, \data_in_frame[21] , 
            n23923, n23922, n23921, n23920, n23919, n23918, n23917, 
            control_mode, \PWMLimit[1] , \PWMLimit[2] , \PWMLimit[3] , 
            \PWMLimit[4] , \PWMLimit[5] , \PWMLimit[6] , \PWMLimit[7] , 
            \PWMLimit[8] , \PWMLimit[9] , n50101, n23834, n23837, 
            n23840, \Ki[2] , \Ki[3] , \Ki[4] , n24240, \data_in[1][6] , 
            \Ki[5] , \data_in[2][1] , \Ki[6] , \Ki[7] , \Kd[1] , \Kd[2] , 
            \Kd[3] , n43459, \Kd[4] , \Kd[5] , \Kd[6] , \Kd[7] , 
            \deadband[0] , n23756, n42561, \PWMLimit[0] , \Kd[0] , 
            \Ki[0] , \Kp[0] , n22, n22833, n40155, n44311, n43709, 
            n3799, n3800, n3801, n3802, n3803, n3804, n3805, n22429, 
            encoder0_position, n3806, n3807, displacement, n3808, 
            encoder1_position, n3809, n3810, n3811, n3812, n3813, 
            pwm, n3814, n44238, n3815, n5022, n23563, n3817, n3818, 
            n3822, n3816, n3820, n3821, n7, n5, n5_adj_3, n44019, 
            n22458, n20136, n44009, n43229, n43236, n43251, n23776, 
            n23779, n23778, n23781, n23784, n23787, n23790, n23793, 
            n23796, n23799, n23803, r_Bit_Index, n23806, n23782, 
            n23785, n23788, n23602, n23716, n4037, n23845, n23791, 
            n23794, n23797, n23844, n23846, n23849, tx_o, tx_enable, 
            n23809, r_Bit_Index_adj_9, n23812, n28794, \r_SM_Main[1] , 
            n24357, r_Rx_Data, LED_c, \r_SM_Main[2] , n23596, n23714, 
            n4015, n23819, n23818, n23817, n23816, n23853, n23815, 
            n23814, n23813, n23751, n28760, n1, n28350, n4, n4_adj_7, 
            n22470, n22462, n4_adj_8, n47207, n47206) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[11] ;
    input GND_net;
    output [23:0]gearBoxRatio;
    input n10;
    input n24253;
    output [7:0]\data_in[0] ;
    input n24252;
    input n24251;
    output [7:0]\data_in_frame[14] ;
    output [7:0]\data_in_frame[19] ;
    input n24250;
    output [7:0]rx_data;
    output \deadband[9] ;
    output \deadband[8] ;
    output \deadband[7] ;
    output \deadband[6] ;
    output \deadband[5] ;
    output \deadband[4] ;
    output \deadband[3] ;
    output \deadband[2] ;
    output \deadband[1] ;
    input n24412;
    output [23:0]setpoint;
    input n24411;
    input n24410;
    input n42279;
    input n24408;
    input n24407;
    input n24406;
    input n24405;
    input n24404;
    input n24403;
    input n24402;
    input n24401;
    input n24400;
    input n24399;
    input n24398;
    input n24397;
    input n24396;
    input n24395;
    input n24394;
    input n24393;
    input n24392;
    input n24391;
    input n24390;
    input n24388;
    input VCC_net;
    output [7:0]byte_transmit_counter;
    input n23822;
    input n24236;
    output [7:0]\data_in[2] ;
    input n24234;
    input n24233;
    input n24228;
    output \data_in[3][2] ;
    input n24227;
    output \data_in[3][3] ;
    input n24226;
    output \data_in[3][4] ;
    input n24225;
    output \data_in[3][5] ;
    input n24223;
    output \data_in[3][7] ;
    input n24222;
    output \data_out_frame[0][2] ;
    input n24221;
    output \data_out_frame[0][3] ;
    input n24220;
    output \data_out_frame[0][4] ;
    input n24217;
    output \data_out_frame[5][2] ;
    output [23:0]IntegralLimit;
    output \Kp[1] ;
    output \Kp[2] ;
    input n24249;
    input n24248;
    output rx_data_ready;
    input n24245;
    output \data_in[1][1] ;
    input n24244;
    output \data_in[1][2] ;
    output \Kp[3] ;
    output \Kp[4] ;
    output [31:0]\FRAME_MATCHER.state ;
    output n47;
    output n3839;
    output n29726;
    output \Kp[5] ;
    output n43231;
    output n43238;
    output n43253;
    output \data_in_frame[1][4] ;
    input n24068;
    output [7:0]\data_in_frame[3] ;
    input n24067;
    input n24066;
    input n24065;
    input n24064;
    input n24063;
    input n24062;
    input n24061;
    input n24243;
    output \data_in[1][3] ;
    output [7:0]\data_in_frame[5] ;
    input n24052;
    input n24051;
    input n24050;
    input n24049;
    output n23533;
    input n24048;
    input n24047;
    input n24046;
    input n24045;
    output \Kp[6] ;
    output \Kp[7] ;
    output \Ki[1] ;
    input n24036;
    output [7:0]\data_in_frame[7] ;
    input n24035;
    input n24034;
    input n24033;
    input n24032;
    input n24031;
    input n24030;
    input n24029;
    input n24242;
    output \data_in[1][4] ;
    input n23825;
    output \data_in_frame[10][6] ;
    input n24004;
    input n24003;
    input n24002;
    input n24001;
    input n24000;
    input n23999;
    input n23998;
    input n23997;
    input n23988;
    input n23987;
    input n23986;
    input n23985;
    input n23984;
    input n23983;
    input n23982;
    output n20342;
    input n23981;
    output \data_in_frame[14][0] ;
    input n24241;
    output \data_in[1][5] ;
    input n23972;
    output [7:0]\data_in_frame[15] ;
    input n23971;
    input n23970;
    input n23969;
    input n23968;
    input n23967;
    input n23966;
    input n23965;
    output n23838;
    output n22456;
    output n43255;
    output \data_in_frame[16][1] ;
    output n23835;
    output n23832;
    output n23823;
    output n23820;
    output n2241;
    output \data_in_frame[18][0] ;
    output \data_in_frame[18][2] ;
    output Kp_23__N_865;
    output n43441;
    input n23940;
    input n23939;
    input n23938;
    output n103;
    input n23937;
    input n23936;
    input n23935;
    input n23934;
    input n23933;
    input Kp_23__N_515;
    output n45225;
    output n122;
    output n44586;
    input n23924;
    output [7:0]\data_in_frame[21] ;
    input n23923;
    input n23922;
    input n23921;
    input n23920;
    input n23919;
    input n23918;
    input n23917;
    output [7:0]control_mode;
    output \PWMLimit[1] ;
    output \PWMLimit[2] ;
    output \PWMLimit[3] ;
    output \PWMLimit[4] ;
    output \PWMLimit[5] ;
    output \PWMLimit[6] ;
    output \PWMLimit[7] ;
    output \PWMLimit[8] ;
    output \PWMLimit[9] ;
    input n50101;
    input n23834;
    input n23837;
    input n23840;
    output \Ki[2] ;
    output \Ki[3] ;
    output \Ki[4] ;
    input n24240;
    output \data_in[1][6] ;
    output \Ki[5] ;
    output \data_in[2][1] ;
    output \Ki[6] ;
    output \Ki[7] ;
    output \Kd[1] ;
    output \Kd[2] ;
    output \Kd[3] ;
    input n43459;
    output \Kd[4] ;
    output \Kd[5] ;
    output \Kd[6] ;
    output \Kd[7] ;
    output \deadband[0] ;
    input n23756;
    input n42561;
    output \PWMLimit[0] ;
    output \Kd[0] ;
    output \Ki[0] ;
    output \Kp[0] ;
    input n22;
    output n22833;
    output n40155;
    input n44311;
    input n43709;
    output n3799;
    output n3800;
    output n3801;
    output n3802;
    output n3803;
    output n3804;
    output n3805;
    output n22429;
    input [23:0]encoder0_position;
    output n3806;
    output n3807;
    input [23:0]displacement;
    output n3808;
    input [23:0]encoder1_position;
    output n3809;
    output n3810;
    output n3811;
    output n3812;
    output n3813;
    input [23:0]pwm;
    output n3814;
    output n44238;
    output n3815;
    output n5022;
    output n23563;
    output n3817;
    output n3818;
    output n3822;
    output n3816;
    output n3820;
    output n3821;
    output n7;
    output n5;
    output n5_adj_3;
    output n44019;
    output n22458;
    output n20136;
    input n44009;
    output n43229;
    output n43236;
    output n43251;
    output n23776;
    output n23779;
    input n23778;
    input n23781;
    input n23784;
    input n23787;
    input n23790;
    input n23793;
    input n23796;
    input n23799;
    input n23803;
    output [2:0]r_Bit_Index;
    input n23806;
    output n23782;
    output n23785;
    output n23788;
    output n23602;
    output n23716;
    output n4037;
    output n23845;
    output n23791;
    output n23794;
    output n23797;
    output n23844;
    input n23846;
    input n23849;
    output tx_o;
    output tx_enable;
    input n23809;
    output [2:0]r_Bit_Index_adj_9;
    input n23812;
    input n28794;
    output \r_SM_Main[1] ;
    input n24357;
    output r_Rx_Data;
    input LED_c;
    output \r_SM_Main[2] ;
    output n23596;
    output n23714;
    output n4015;
    input n23819;
    input n23818;
    input n23817;
    input n23816;
    input n23853;
    input n23815;
    input n23814;
    input n23813;
    input n23751;
    output n28760;
    output n1;
    output n28350;
    output n4;
    output n4_adj_7;
    output n22470;
    output n22462;
    output n4_adj_8;
    output n47207;
    output n47206;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n24202;
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(94[12:26])
    
    wire n24201, n24200, n24199, n24198, n43596, n24197, n24276, 
        n24275, n24274, n24273, n24272, n24271, n24270, n24196, 
        n36947;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(112[11:12])
    
    wire n36948, n2, n36946, n1507, n36935, n36936, n40198, n43691, 
        n24195;
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(94[12:26])
    
    wire n2_adj_3110, n36934, n2_adj_3111, n36945, n24194, n24193, 
        n24269, n24192, n24191, n24190, n24189, n24188, n24268, 
        n24267, n24266, n24265, n24264, n24263, n24262, n24261, 
        n24260, n24259, n24258, n24257, n24256, n24255, n24254, 
        n23126, n43751, n6, n43518, n40163, n24187;
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(94[12:26])
    
    wire n24186, n8, n43226;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(93[12:25])
    
    wire n24053, n24421, n24420, n24419, n24418, n24417, n24416, 
        n24415, n24414, n24413;
    wire [7:0]byte_transmit_counter_c;   // verilog/coms.v(99[12:33])
    
    wire n24185, n24184, n27275, n24183, n24182, n24181, n24232, 
        n24180, n24231;
    wire [7:0]\data_in[2]_c ;   // verilog/coms.v(92[12:19])
    
    wire n24179;
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(94[12:26])
    
    wire n24230;
    wire [7:0]\data_in[3] ;   // verilog/coms.v(92[12:19])
    
    wire n24178, n24229, n24177, n24176, n24175, n24174, n24173, 
        n24224, n24172, n24171;
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(94[12:26])
    
    wire n24219;
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(94[12:26])
    
    wire n24218, n24216, n24215, n24214, n24213, n24212, n24303, 
        n24302, n24301, n24300, n24299, n24298, n24297, n24170, 
        n24169, n24168, n24167, n24166, n24211;
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(94[12:26])
    
    wire n24210, n24209, n24208, n24207, n24206, n24165, n24054, 
        n24164, n24205, n24204, n24163;
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(94[12:26])
    
    wire n24296, n24162, n24055, n24161, n24160, n24159, n24158, 
        n24157, n24156, n24155;
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(94[12:26])
    
    wire n24154, n24153, n24152, n24151, n24247;
    wire [7:0]\data_in[0]_c ;   // verilog/coms.v(92[12:19])
    
    wire n24150, n24246;
    wire [7:0]\data_in[1] ;   // verilog/coms.v(92[12:19])
    
    wire n24149, n24148, n24147;
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(94[12:26])
    
    wire n24146, n24145, n24144, n24143, n24142, \FRAME_MATCHER.rx_data_ready_prev , 
        n24141, n24140, n24312, n24139;
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(94[12:26])
    
    wire n24138, n24137, n24136, n24135, n24056, n24311, n24310, 
        n24134, n24133, n24305, n24132, n24057, n24295, n24294, 
        n24131;
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(94[12:26])
    
    wire n24058, n24130, n24129, n24128, n24127, n24126, n24125, 
        n24124, n24123;
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(94[12:26])
    
    wire n24122, n24121, n24120, n24119, n24118, n6_adj_3112, n24117, 
        n2_adj_3113, n36944, n2_adj_3114, n36933, n24059, n24116, 
        n24115;
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(94[12:26])
    
    wire n24114, n24060, n28723, n47090, n29738, n45217, n44005, 
        n24113, n24112, n24111, n24110, n24109, n24108, n24107;
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(94[12:26])
    
    wire n24106, n24293, n24105, n24104, n24103, n24102, n24101, 
        n24100, n24099;
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(94[12:26])
    
    wire n24098, n24097, n24096, n24095, n24094, n24309, n24093, 
        n24092, n24091;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(93[12:25])
    
    wire n24090, n24089, n24088, n43235, n24087, n24086, n43247, 
        n24085, n24084;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(93[12:25])
    
    wire n24083, n24082, n24081, n24080, n24079, n22453, n28434, 
        n2123, n24078, n24077, n24076;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(93[12:25])
    
    wire n24075, n24074, n24073, n24304, n24072, n24071, n24070, 
        n24069, n20432, Kp_23__N_458, Kp_23__N_1179, n7_c, n23385, 
        n22796, n16, n22801, n22_c, n23176, n22928, n6_adj_3115, 
        n15, n39466, n10_adj_3116, n23242, n20, n8_adj_3117, n23183, 
        n24, n22953, n23367, n16_adj_3118, n24044;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(93[12:25])
    
    wire n24043, n24042, n24041, n24040, n24039, n24038, n24037, 
        n24292, n22334, n22451, n24291, n24290, n24308, n8_adj_3119, 
        n24028;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(93[12:25])
    
    wire n24027, n24026, n24025, n24024, n24023, n24022, n24021, 
        n24020;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(93[12:25])
    
    wire n24019, n24018, n24017, n24016, n24015, n24014, n24013, 
        n24012;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(93[12:25])
    
    wire n24011, n22343, n2854, n24010, n2_adj_3120, n36943, n10_adj_3121, 
        n50095, n50098, n23828, n50083, n50086;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(93[12:25])
    
    wire n23989, n24009, n24008, n19, n47245, n50089, n24007, 
        n17, n16_adj_3122, n50092, n24006, n24005, n47217, n5_c, 
        n45342, n45343, n50077, n45340, n45339, n50080, n45348, 
        n45349, n50071, n45346, n45345, n50074, n23996, n50065, 
        n23995, n50068, n23994, n23993, n50059, n23992, n50062, 
        n23991, n23990, n50053, n50056, n50047, n50050, n50041, 
        n50044;
    wire [7:0]\data_in_frame[14]_c ;   // verilog/coms.v(93[12:25])
    
    wire n23973, n23974, n23975, n23976, n23977, n23978, n23979, 
        n23980, n59, n54, n44574;
    wire [31:0]\FRAME_MATCHER.state_c ;   // verilog/coms.v(109[11:16])
    
    wire n42473, n8_adj_3123, n22442, n2_adj_3124, n20099, n42605, 
        n2_adj_3125, n36942, n42607, n28314, n42609, n42611, n28316, 
        n2_adj_3126, n36932, n75, n42613, n50035, n50038, n7_adj_3127, 
        n42603, n42551, n28291, n28289, n42481, n42663, n42519, 
        n42661, n42507, n7_adj_3128, n8_adj_3129, n42601, n42555, 
        n42599, n42427, n42593, n42553, n42597, n42589, n42681, 
        n42509, n42677, n42557, n42627, n42559, n42625, n42511, 
        n42623, n42501, n42621, n42563, n42619, n42565, n42617, 
        n42567, n42615, n42569, n42571, n42573, n42575, n42577, 
        n28698, n42579, n42581, n42675, n42493, n42491, n42727, 
        n42487, n50100, n43398, n23557;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(94[12:26])
    
    wire n44472, n22915, n43410, n44636, n44772, n43282, n43283, 
        n45019;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(94[12:26])
    
    wire n44400, n44383, n44979, n44983, n45043, n44955, n44821, 
        n36967, n2_adj_3130, n36941, n23964;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(93[12:25])
    
    wire n2_adj_3131, n36940, n2_adj_3132, n3, n43132, n43245, n6_adj_3133, 
        n43127, n43273, n43271, n10_adj_3134, n14, n10_adj_3135, 
        n14_adj_3136, n43635, n43287, n40234, n45002, Kp_23__N_804, 
        n43391, n43712, n16_adj_3137, n39479, n39570, n17_adj_3138;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(93[12:25])
    
    wire n15_adj_3139, n43426, n43678, n43684, n12, n43827, n44630, 
        n43587, n43512;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(93[12:25])
    
    wire n16_adj_3140, n43849, n43739, n17_adj_3141, n22827, n43789, 
        n23346, n6_adj_3142, n43733, n43852, n22728, n43614, n43885, 
        n43727, n43508, n16_adj_3143, n43381, n17_adj_3144, n22750, 
        n43843, n43730, n43490, n43801, n18, n43675, n20_adj_3145, 
        n43867, n16_adj_3146, n40149, n2_adj_3147, n3_adj_3148, n2_adj_3149, 
        n3_adj_3150, n2_adj_3151, n3_adj_3152, n2_adj_3153, n3_adj_3154, 
        n2_adj_3155, n3_adj_3156, n2_adj_3157, n3_adj_3158, n2_adj_3159, 
        n3_adj_3160, n2_adj_3161, n3_adj_3162, n2_adj_3163, n3_adj_3164, 
        n2_adj_3165, n3_adj_3166, n2_adj_3167, n3_adj_3168, n2_adj_3169, 
        n3_adj_3170, n2_adj_3171, n3_adj_3172, n3_adj_3173, n3_adj_3174, 
        n3_adj_3175, n3_adj_3176, n3_adj_3177, n3_adj_3178, n3_adj_3179, 
        n2_adj_3180, n3_adj_3181, n2_adj_3182, n3_adj_3183, n2_adj_3184, 
        n3_adj_3185, n2_adj_3186, n3_adj_3187, n2_adj_3188, n3_adj_3189, 
        n3_adj_3190, n3_adj_3191, n3_adj_3192, n2_adj_3193, n3_adj_3194, 
        n2_adj_3195, n3_adj_3196, n23963, n23219, n40161, n40127, 
        n40169, n22_adj_3197, n20_adj_3198, n36966, n36939, n36965, 
        n36931, n23829, n36964, n36930, n16_adj_3199, n24_adj_3200, 
        n23826, n36963, n36938, n24307, n23962, n23961, n23960, 
        n23959, n43724, n43501, n23078, n43528, n8_adj_3201, n36962, 
        n10_adj_3202, n23958, n43278, n23212, n23957, n23956, n23955, 
        n43471, n23169, n23954, n23953, n43557, n36961, n43367;
    wire [2:0]r_SM_Main_2__N_2747;
    
    wire tx_active, n7_adj_3203, tx_transmit_N_2639, n10_adj_3204, n43569, 
        n23952, n23951, n23950, n23949, n23948, n23947, n23946, 
        n23945, n43343, n23209, n23944, n23943, n23942, n23941, 
        n43879, n50029, n744, n43873, n43706, n4_c, n737, n22443, 
        n20098, n3758, n43833, n43802, n139, n43263, n8_adj_3205, 
        n36960, n36959, n23932;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(93[12:25])
    
    wire n23931, n23930, n23929, n23928, n23927, n36958, n43301, 
        n43644, n10_adj_3206, n12_adj_3207, n50032, n43894, n43754, 
        n43855, n10_adj_3208, n40131, n43462, n10_adj_3209, Kp_23__N_325, 
        n43474, n22454, n39443, n6_adj_3210, n39561, n28284, n23926, 
        n23925, n36937, n23916, n23915, n23914, n23913, n23912, 
        n23911, n23910, n23909, n23908, n23907, n23906, n23905, 
        n28060, n36957, n23903, n23902, n23901, n22501, n43563, 
        n43538, n43770, n10_adj_3211, n40129, n42, n36956, n8_adj_3212, 
        n6_adj_3213, n36955, n36954, n36953, n43352, n39500, n43308, 
        n20125, n37, n44497, n44479, n6_adj_3214, n40137, n43718, 
        n6_adj_3215, n43888, n24289, n43453, n22605, n24288, n43477, 
        n23251, n39281, n24287, n50023, n50026, n24239;
    wire [0:0]n2416;
    
    wire n44089, n36952, n43703, n24286, n23254, n10_adj_3216, n39470, 
        n24238, n43397, n10_adj_3217, n22721, n27276, n24285, n24320, 
        n24319, n24318, n24317, n5_adj_3218, n4_adj_3219, n24284, 
        n12_adj_3220, n24283, n43837, n22771, n43767, n24282, n24281, 
        n6_adj_3221, n24306, n43830, n43821, n43566, n43748, n52, 
        n6_adj_3222, n59_adj_3223, n43858, n56, n43375, n43804, 
        n54_adj_3224, n55, n43870, n43299, n53, n43388, n58, n64, 
        n43626, n57, n65, n43783, n10_adj_3225, n23436, n43742, 
        n43525, n43541, n6_adj_3226, n21061, n24280, n43429, n43355, 
        n43861, n22746, n43694, n43641, n36951, n36950, n24279, 
        n24278, n24277, n43882, n23757, n24203, n2_adj_3227, n3_adj_3228, 
        n11, n12_adj_3229, n50011, n24316, n24315, n24314, n24313, 
        n43846, n12_adj_3230, n23742, n23741, n23740, n23739, n23738, 
        n23737, n23736, Kp_23__N_785, n43349, n26, n23735, n23734, 
        n9, n8_adj_3231, n50014, n24_adj_3232, n43593, n25, n23, 
        n36949, n161, n40194, n8_adj_3233, n43671, n43824, n12_adj_3234, 
        n8_adj_3235, n43415, n12_adj_3236, n43795, n43371, n43544, 
        n14_adj_3237, n15_adj_3239, n43423, n6_adj_3240, n43758, n23358, 
        n23468, Kp_23__N_328, n43495, n43480, n18_adj_3241, n30, 
        n43378, n28, n43655, n43780, n29, n43394, n27, n50005, 
        n15_adj_3242, n14_adj_3243, n23202, n43318, n43584, n12_adj_3244, 
        n7_adj_3245, n12_adj_3246, n44324, n8_adj_3247, n12_adj_3248, 
        n44580, n45075, n44856, n50008, n107, n44965, n14_adj_3249, 
        n15_adj_3250, n44172, n8_adj_3251, n18_adj_3252, n44367, n26_adj_3253, 
        n44888, n24_adj_3254, n30_adj_3255, n44977, n8_adj_3256, n7_adj_3257, 
        n20_adj_3258, n28_adj_3259, n32, n19_adj_3260, n8_adj_3261, 
        n47239, n19_adj_3262, n47504, n5_adj_3263, n45301, n45302, 
        n45273, n45275, n45274, n49999, n50002, n18_adj_3264, n16_adj_3265, 
        n20_adj_3266, n6_adj_3267, n4_adj_3268, n45252, n38, n39, 
        n37_adj_3269, n45248, n46, n45250;
    wire [31:0]\FRAME_MATCHER.state_31__N_1924 ;
    
    wire n23530;
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n25425, n5024, n19_adj_3270, n45271, n47677, n5_adj_3271, 
        n45272, n47022, n45297, n45299, n19_adj_3272, n45268, n47670, 
        n5_adj_3273, n49996, n45269, n45294, n45296, n19_adj_3274, 
        n47665, n5_adj_3275, n45265, n49990, n45266, n45291, n45293, 
        n49966, n45292, n19_adj_3276, n45262, n49984, n45263, n48879;
    wire [7:0]tx_data;   // verilog/coms.v(102[13:20])
    
    wire n47202, n6_adj_3277, n5_adj_3278, n45282, n45284, n49978, 
        n49972, n45283, n47199, n19_adj_3279, n6_adj_3280, n5_adj_3281, 
        n45307, n45308, n45279, n45281, n45280, n19_adj_3282, n47645, 
        n5_adj_3283, n45304, n45305, n45276, n45278, n45277, n47095, 
        n23_adj_3284, n31, n63, n22133, n43450, n8_adj_3287, n22984, 
        n23259, n39498, n43284, n7_adj_3288, n44835, n43608, n43652, 
        n6_adj_3289, n1713, n43314, n39866, n23282, n43620, n49993, 
        n43786, n43611, n43605, n49987, n22809, n44887, n49981, 
        n43581, n43777, n43590, n1692, n43688, n39462, n10_adj_3290, 
        n10_adj_3291, n40119, n43697, n14_adj_3292, n39990, n23405, 
        n44973, n6_adj_3293, n1784, n43599, n43326, n39781, n12_adj_3294, 
        n43813, n43385, n39404, n43807, n43465, n20_adj_3295, n23381, 
        n43647, n19_adj_3296, n22146, n21, n44765, n12_adj_3297, 
        n43409, n14_adj_3298, n43295, n22166, n43638, n43810, n24_adj_3299, 
        n22190, n17_adj_3300, n43864, n43329, n22_adj_3301, n40167, 
        n43891, n26_adj_3302, n22126, n10_adj_3303, n43554, n14_adj_3304, 
        n43617, n1592, n43403, n22596, n39504, n12_adj_3305, n39844, 
        n43292, n6_adj_3306, n43419, n1503, n23337, n43447, n43412, 
        n23331, n52_adj_3307, n56_adj_3308, n58_adj_3309, n43764, 
        n59_adj_3310, n43438, n57_adj_3311, n23110, n43681, n43456, 
        n54_adj_3312, n7_adj_3313, n62, n60, n66, n43876, n43340, 
        n43484, n22142, n53_adj_3314, n43325, n23081, n23119, n23327, 
        n10_adj_3315, n14_adj_3316, n22599, n16_adj_3317, n43332, 
        n43572, n22_adj_3318, n43487, n14_adj_3319, n49269, n43773, 
        n24_adj_3320, n23_adj_3321, n16_adj_3322, n1512, n43400, n22_adj_3323, 
        n43363, n20_adj_3324, n24_adj_3325, n43305, n43623, n40144, 
        n23085, n43522, n43667, n20_adj_3326, n43818, n19_adj_3327, 
        n21_adj_3328, n39476, n43792, n44734, n40117, n6_adj_3329, 
        n22972, n6_adj_3330, n23323, n43660, n16_adj_3331, n17_adj_3332, 
        n43798, n43498, n22994, n43629, n40171, n43505, n43700, 
        n14_adj_3333, n43840, n15_adj_3334, n43346, n43663, n43468, 
        n6_adj_3335, n14_adj_3336, n15_adj_3337, n43721, n43358, n6_adj_3338, 
        n14_adj_3339, n10_adj_3340, n12_adj_3341, n63_adj_3342, n2119, 
        n22448, n49975, n7_adj_3344;
    wire [31:0]\FRAME_MATCHER.state_31__N_1860 ;
    wire [31:0]\FRAME_MATCHER.state_31__N_1892 ;
    
    wire n6_adj_3345, n7_adj_3346, n7_adj_3347, n4_adj_3348, n22441, 
        n43218, n44728, n4_adj_3349, n10_adj_3350, n22447, n27228, 
        n12_adj_3351, n8_adj_3352, n26_adj_3353, n36, n44869, n34, 
        n40, n38_adj_3354, n39_adj_3355, n37_adj_3356, n15_adj_3357, 
        n6_adj_3358, n6_adj_3359, n44946, n22475, n10_adj_3360, n22564, 
        n16_adj_3361, n17_adj_3362, n22432, n10_adj_3363, n14_adj_3364, 
        n45152, n12_adj_3365, n18_adj_3366, n45254, n12_adj_3367, 
        n25797, n21_adj_3368, n49969, n49963;
    
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n24202));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n24201));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n24200));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n24199));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n24198));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n43596));   // verilog/coms.v(67[16:27])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n24197));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n24276));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n24275));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n24274));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n24273));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n24272));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n24271));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n24270));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n24196));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_20 (.CI(n36947), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n36948));
    SB_LUT4 add_41_19_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n36946), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_8 (.CI(n36935), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n36936));
    SB_CARRY add_41_19 (.CI(n36946), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n36947));
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n10), .I3(n40198), .O(n43691));   // verilog/coms.v(67[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n24195));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_7_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n36934), .O(n2_adj_3110)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_7 (.CI(n36934), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n36935));
    SB_LUT4 add_41_18_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n36945), .O(n2_adj_3111)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_18 (.CI(n36945), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n36946));
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n24194));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n24193));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n24269));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n24192));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n24191));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n24190));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n24189));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n24188));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n24268));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n24267));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n24266));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n24265));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n24264));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n24263));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n24262));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n24261));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n24260));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n24259));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n24258));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n24257));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n24256));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n24255));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n24254));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n24253));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n24252));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n24251));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_4_lut (.I0(n23126), .I1(n43751), .I2(\data_in_frame[14] [4]), 
            .I3(\data_in_frame[19] [2]), .O(n6));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_828 (.I0(n23126), .I1(n43751), .I2(\data_in_frame[14] [4]), 
            .I3(n43518), .O(n40163));
    defparam i1_2_lut_4_lut_adj_828.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n24250));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n24187));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n24186));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10638_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n24053));
    defparam i10638_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF deadband_i0_i9 (.Q(\deadband[9] ), .C(clk32MHz), .D(n24421));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i8 (.Q(\deadband[8] ), .C(clk32MHz), .D(n24420));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i7 (.Q(\deadband[7] ), .C(clk32MHz), .D(n24419));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i6 (.Q(\deadband[6] ), .C(clk32MHz), .D(n24418));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i5 (.Q(\deadband[5] ), .C(clk32MHz), .D(n24417));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i4 (.Q(\deadband[4] ), .C(clk32MHz), .D(n24416));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i3 (.Q(\deadband[3] ), .C(clk32MHz), .D(n24415));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i2 (.Q(\deadband[2] ), .C(clk32MHz), .D(n24414));   // verilog/coms.v(125[12] 284[6])
    SB_DFF deadband_i0_i1 (.Q(\deadband[1] ), .C(clk32MHz), .D(n24413));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n24412));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n24411));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n24410));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n42279));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n24408));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n24407));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n24406));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n24405));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n24404));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n24403));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n24402));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n24401));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n24400));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n24399));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n24398));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n24397));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n24396));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n24395));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n24394));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n24393));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n24392));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n24391));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n24390));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(VCC_net), .D(n24388));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter_c[1]), .C(clk32MHz), 
           .D(n23822));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n24185));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n24236));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n24184));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n27275));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n24183));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n24234));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n24182));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n24233));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n24181));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n24232));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n24180));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2]_c [7]), .C(clk32MHz), .D(n24231));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n24179));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n24230));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n24178));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n24229));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n24177));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3][2] ), .C(clk32MHz), .D(n24228));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n24176));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3][3] ), .C(clk32MHz), .D(n24227));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n24175));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3][4] ), .C(clk32MHz), .D(n24226));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n24174));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3][5] ), .C(clk32MHz), .D(n24225));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n24173));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n24224));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n24172));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3][7] ), .C(clk32MHz), .D(n24223));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n24171));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i3 (.Q(\data_out_frame[0][2] ), .C(clk32MHz), 
           .D(n24222));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk32MHz), 
           .D(n24221));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk32MHz), 
           .D(n24220));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n24219));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n24218));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5][2] ), .C(clk32MHz), 
           .D(n24217));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n24216));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n24215));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n24214));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n24213));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n24212));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n24303));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n24302));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n24301));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n24300));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n24299));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n24298));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n24297));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n24170));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n24169));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n24168));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n24167));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n24166));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n24211));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n24210));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n24209));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n24208));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n24207));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n24206));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n24165));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10639_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n24054));
    defparam i10639_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n24164));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n24205));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n24204));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n24163));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n24296));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n24162));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n24249));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10640_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n24055));
    defparam i10640_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n24161));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n24160));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n24248));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n24159));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n24158));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n24157));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n24156));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n24155));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n24154));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n24153));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n24152));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n24151));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0]_c [7]), .C(clk32MHz), .D(n24247));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n24150));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n24246));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n24149));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n24148));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n24147));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n24146));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n24145));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n24144));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n24143));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n24142));   // verilog/coms.v(125[12] 284[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3221  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n24141));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n24140));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n24312));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n24139));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n24138));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n24137));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n24136));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1][1] ), .C(clk32MHz), .D(n24245));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n24135));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10641_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n24056));
    defparam i10641_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n24311));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1][2] ), .C(clk32MHz), .D(n24244));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n24310));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n24134));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n24133));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n24305));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n24132));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10642_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n24057));
    defparam i10642_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n24295));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n24294));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n24131));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10643_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n24058));
    defparam i10643_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n24130));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n24129));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n24128));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n24127));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n24126));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n24125));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n24124));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n24123));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n24122));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n24121));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n24120));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n24119));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n24118));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3112));
    defparam i2_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n24117));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_17_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n36944), .O(n2_adj_3113)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_41_6_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n36933), .O(n2_adj_3114)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_17 (.CI(n36944), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n36945));
    SB_LUT4 i10644_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n24059));
    defparam i10644_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n24116));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n24115));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n24114));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10645_3_lut_4_lut (.I0(n8), .I1(n43226), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n24060));
    defparam i10645_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32399_4_lut (.I0(n47), .I1(n6_adj_3112), .I2(n28723), .I3(\FRAME_MATCHER.state [0]), 
            .O(n47090));   // verilog/coms.v(109[11:16])
    defparam i32399_4_lut.LUT_INIT = 16'hfcfe;
    SB_LUT4 i29717_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n29738), .I3(GND_net), .O(n45217));
    defparam i29717_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 i16377_4_lut (.I0(n45217), .I1(n47090), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n44005), .O(n3839));   // verilog/coms.v(109[11:16])
    defparam i16377_4_lut.LUT_INIT = 16'hcfc5;
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n24113));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n24112));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n24111));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n3839), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n29726));   // verilog/coms.v(109[11:16])
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n24110));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n24109));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n24108));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n24107));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n24106));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n24293));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n24105));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n24104));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n24103));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 equal_64_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(149[7:23])
    defparam equal_64_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n24102));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n24101));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n24100));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n24099));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n24098));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n24097));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n24096));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n24095));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43226), .I3(\FRAME_MATCHER.i [0]), .O(n43231));   // verilog/coms.v(149[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n24094));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n24309));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n24093));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n24092));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n24091));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n24090));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n24089));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n24088));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_829 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43235), .I3(\FRAME_MATCHER.i [0]), .O(n43238));   // verilog/coms.v(149[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_829.LUT_INIT = 16'hfbff;
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n24087));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n24086));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_830 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43247), .I3(\FRAME_MATCHER.i [0]), .O(n43253));   // verilog/coms.v(149[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_830.LUT_INIT = 16'hfbff;
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n24085));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n24084));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n24083));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n24082));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n24081));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1][4] ), .C(clk32MHz), 
           .D(n24080));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n24079));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i15291_3_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n22453), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n28434), .O(n2123));   // verilog/coms.v(248[5:27])
    defparam i15291_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n24078));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n24077));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n24076));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n24075));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n24074));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n24073));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n24304));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n24072));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n24071));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n24070));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n24069));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n24068));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n24067));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n24066));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n24065));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n24064));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n24063));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n24062));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n24061));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n24060));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n24059));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1][3] ), .C(clk32MHz), .D(n24243));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n24058));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n24057));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n24056));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_4_lut (.I0(n20432), .I1(Kp_23__N_458), .I2(Kp_23__N_1179), 
            .I3(\data_in_frame[5] [6]), .O(n7_c));
    defparam i2_4_lut.LUT_INIT = 16'h3bce;
    SB_LUT4 i9_4_lut (.I0(n23385), .I1(n22796), .I2(n16), .I3(n22801), 
            .O(n22_c));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_831 (.I0(n23176), .I1(n7_c), .I2(n22928), .I3(n6_adj_3115), 
            .O(n15));
    defparam i2_4_lut_adj_831.LUT_INIT = 16'hffef;
    SB_LUT4 i7_3_lut (.I0(n39466), .I1(n10_adj_3116), .I2(n23242), .I3(GND_net), 
            .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n15), .I1(n22_c), .I2(n8_adj_3117), .I3(n23183), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n22953), .I1(n24), .I2(n20), .I3(n23367), 
            .O(n47));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_3_lut (.I0(n29738), .I1(n47), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n16_adj_3118));   // verilog/coms.v(109[11:16])
    defparam i22_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n24055));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n24054));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n24053));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n24052));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n24051));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n24050));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n24049));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n16_adj_3118), .I3(n44005), .O(n23533));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n24048));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n24047));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n24046));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n24045));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n24044));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n24043));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n24042));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n24041));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n24040));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n24039));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n24038));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n24037));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n24292));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22334), 
            .I2(\FRAME_MATCHER.state [0]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n22451));   // verilog/coms.v(156[5:29])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n24291));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n24290));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n24308));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n24036));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n24035));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10622_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n24037));
    defparam i10622_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n24034));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n24033));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n24032));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n24031));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10623_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n24038));
    defparam i10623_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10624_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n24039));
    defparam i10624_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n24030));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n24029));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n24028));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n24027));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n24026));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n24025));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n24024));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n24023));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n24022));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n24021));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n24020));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n24019));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n24018));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n24017));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n24016));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10625_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n24040));
    defparam i10625_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10626_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n24041));
    defparam i10626_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10627_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n24042));
    defparam i10627_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n24015));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n24014));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10628_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n24043));
    defparam i10628_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n24013));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n24012));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10629_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43226), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n24044));
    defparam i10629_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n24011));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i15038_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n22343), .I3(\FRAME_MATCHER.i [31]), .O(n2854));
    defparam i15038_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n24010));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_16_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n36943), .O(n2_adj_3120)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1842_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_3121));
    defparam i1842_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_DFF data_in_0___i13 (.Q(\data_in[1][4] ), .C(clk32MHz), .D(n24242));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_6 (.CI(n36933), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n36934));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n50095));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n50095_bdd_4_lut (.I0(n50095), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n50098));
    defparam n50095_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_41_16 (.CI(n36943), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n36944));
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter_c[2]), .C(clk32MHz), 
           .D(n23825));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter_c[3]), .C(clk32MHz), 
           .D(n23828));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50083_bdd_4_lut_4_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter_c[2]), .I3(n50083), .O(n50086));
    defparam n50083_bdd_4_lut_4_lut.LUT_INIT = 16'hfc02;
    SB_LUT4 i10574_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n23989));
    defparam i10574_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n24009));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n24008));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter_c[1]), 
            .I1(n19), .I2(n47245), .I3(byte_transmit_counter_c[2]), .O(n50089));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n24007));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50089_bdd_4_lut (.I0(n50089), .I1(n17), .I2(n16_adj_3122), 
            .I3(byte_transmit_counter_c[2]), .O(n50092));
    defparam n50089_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10][6] ), .C(clk32MHz), 
           .D(n24006));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n24005));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_34568 (.I0(byte_transmit_counter_c[1]), 
            .I1(n47217), .I2(n5_c), .I3(byte_transmit_counter_c[2]), .O(n50083));
    defparam byte_transmit_counter_1__bdd_4_lut_34568.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n24004));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n24003));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n24002));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_34563 (.I0(byte_transmit_counter_c[1]), 
            .I1(n45342), .I2(n45343), .I3(byte_transmit_counter_c[2]), 
            .O(n50077));
    defparam byte_transmit_counter_1__bdd_4_lut_34563.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n24001));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50077_bdd_4_lut (.I0(n50077), .I1(n45340), .I2(n45339), .I3(byte_transmit_counter_c[2]), 
            .O(n50080));
    defparam n50077_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n24000));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n23999));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_34558 (.I0(byte_transmit_counter_c[1]), 
            .I1(n45348), .I2(n45349), .I3(byte_transmit_counter_c[2]), 
            .O(n50071));
    defparam byte_transmit_counter_1__bdd_4_lut_34558.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n23998));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50071_bdd_4_lut (.I0(n50071), .I1(n45346), .I2(n45345), .I3(byte_transmit_counter_c[2]), 
            .O(n50074));
    defparam n50071_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n23997));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n23996));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34573 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n50065));
    defparam byte_transmit_counter_0__bdd_4_lut_34573.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n23995));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50065_bdd_4_lut (.I0(n50065), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n50068));
    defparam n50065_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n23994));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n23993));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34548 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n50059));
    defparam byte_transmit_counter_0__bdd_4_lut_34548.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n23992));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50059_bdd_4_lut (.I0(n50059), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n50062));
    defparam n50059_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n23991));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n23990));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34543 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n50053));
    defparam byte_transmit_counter_0__bdd_4_lut_34543.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n23989));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50053_bdd_4_lut (.I0(n50053), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n50056));
    defparam n50053_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n23988));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n23987));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34538 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n50047));
    defparam byte_transmit_counter_0__bdd_4_lut_34538.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n23986));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50047_bdd_4_lut (.I0(n50047), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n50050));
    defparam n50047_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n23985));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10575_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n23990));
    defparam i10575_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n23984));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34533 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n50041));
    defparam byte_transmit_counter_0__bdd_4_lut_34533.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n23983));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50041_bdd_4_lut (.I0(n50041), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n50044));
    defparam n50041_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n23982));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10576_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n23991));
    defparam i10576_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10577_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n23992));
    defparam i10577_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10578_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n23993));
    defparam i10578_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10579_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n23994));
    defparam i10579_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_62_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3119));
    defparam equal_62_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i10580_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n23995));
    defparam i10580_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_832 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43226), .I3(\FRAME_MATCHER.i [0]), .O(n20342));
    defparam i1_2_lut_3_lut_4_lut_adj_832.LUT_INIT = 16'hf7ff;
    SB_LUT4 i10581_3_lut_4_lut (.I0(n8), .I1(n43247), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n23996));
    defparam i10581_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n23981));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10558_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[7]), 
            .I3(\data_in_frame[14]_c [7]), .O(n23973));
    defparam i10558_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10559_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[6]), 
            .I3(\data_in_frame[14]_c [6]), .O(n23974));
    defparam i10559_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10560_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[5]), 
            .I3(\data_in_frame[14]_c [5]), .O(n23975));
    defparam i10560_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10561_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n23976));
    defparam i10561_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10562_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[3]), 
            .I3(\data_in_frame[14]_c [3]), .O(n23977));
    defparam i10562_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10563_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[2]), 
            .I3(\data_in_frame[14]_c [2]), .O(n23978));
    defparam i10563_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10564_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[1]), 
            .I3(\data_in_frame[14]_c [1]), .O(n23979));
    defparam i10564_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10565_3_lut_4_lut (.I0(n8_adj_3119), .I1(n43247), .I2(rx_data[0]), 
            .I3(\data_in_frame[14][0] ), .O(n23980));
    defparam i10565_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_833 (.I0(n59), .I1(n54), .I2(n44574), .I3(\FRAME_MATCHER.state_c [29]), 
            .O(n42473));
    defparam i1_2_lut_4_lut_adj_833.LUT_INIT = 16'hfe00;
    SB_LUT4 i80_2_lut_4_lut (.I0(n59), .I1(n54), .I2(n44574), .I3(\FRAME_MATCHER.state_c [31]), 
            .O(n8_adj_3123));
    defparam i80_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_834 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [5]), .O(n42605));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_834.LUT_INIT = 16'hdc00;
    SB_LUT4 add_41_15_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n36942), .O(n2_adj_3125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_835 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [6]), .O(n42607));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_835.LUT_INIT = 16'hdc00;
    SB_LUT4 i14915_2_lut_4_lut (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [7]), .O(n28314));   // verilog/coms.v(112[11:12])
    defparam i14915_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_836 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [8]), .O(n42609));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_836.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_837 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [9]), .O(n42611));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_837.LUT_INIT = 16'hdc00;
    SB_LUT4 i14916_2_lut_4_lut (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [10]), .O(n28316));   // verilog/coms.v(112[11:12])
    defparam i14916_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14][0] ), .C(clk32MHz), 
           .D(n23980));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_5_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n36932), .O(n2_adj_3126)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14]_c [1]), .C(clk32MHz), 
           .D(n23979));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter_c[4]), .C(clk32MHz), 
           .D(n75));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_4_lut_adj_838 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [11]), .O(n42613));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_838.LUT_INIT = 16'hdc00;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34528 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n50035));
    defparam byte_transmit_counter_0__bdd_4_lut_34528.LUT_INIT = 16'he4aa;
    SB_DFF data_in_0___i14 (.Q(\data_in[1][5] ), .C(clk32MHz), .D(n24241));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50035_bdd_4_lut (.I0(n50035), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n50038));
    defparam n50035_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(clk32MHz), 
            .D(n7_adj_3127), .S(n8_adj_3123));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(clk32MHz), 
            .D(n42603), .S(n42551));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(clk32MHz), 
            .D(n28291), .S(n42473));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(clk32MHz), 
            .D(n28289), .S(n42481));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(clk32MHz), 
            .D(n42663), .S(n42519));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(clk32MHz), 
            .D(n42661), .S(n42507));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(clk32MHz), 
            .D(n7_adj_3128), .S(n8_adj_3129));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(clk32MHz), 
            .D(n42601), .S(n42555));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(clk32MHz), 
            .D(n42599), .S(n42427));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(clk32MHz), 
            .D(n42593), .S(n42553));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(clk32MHz), 
            .D(n42597), .S(n42589));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(clk32MHz), 
            .D(n42681), .S(n42509));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(clk32MHz), 
            .D(n42677), .S(n42557));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(clk32MHz), 
            .D(n42627), .S(n42559));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(clk32MHz), 
            .D(n42625), .S(n42511));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(clk32MHz), 
            .D(n42623), .S(n42501));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(clk32MHz), 
            .D(n42621), .S(n42563));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(clk32MHz), 
            .D(n42619), .S(n42565));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(clk32MHz), 
            .D(n42617), .S(n42567));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(clk32MHz), 
            .D(n42615), .S(n42569));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(clk32MHz), 
            .D(n42613), .S(n42571));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(clk32MHz), 
            .D(n28316), .S(n42573));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(clk32MHz), 
            .D(n42611), .S(n42575));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(clk32MHz), 
            .D(n42609), .S(n42577));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(clk32MHz), 
            .D(n28314), .S(n28698));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(clk32MHz), 
            .D(n42607), .S(n42579));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(clk32MHz), 
            .D(n42605), .S(n42581));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(clk32MHz), 
            .D(n42675), .S(n42493));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n42491), .S(n42727));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n42487), .S(n50100));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14]_c [2]), .C(clk32MHz), 
           .D(n23978));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_15 (.CI(n36942), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n36943));
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14]_c [3]), .C(clk32MHz), 
           .D(n23977));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n23976));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14]_c [5]), .C(clk32MHz), 
           .D(n23975));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14]_c [6]), .C(clk32MHz), 
           .D(n23974));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14]_c [7]), .C(clk32MHz), 
           .D(n23973));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n23972));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n23971));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_4_lut_adj_839 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [12]), .O(n42615));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_839.LUT_INIT = 16'hdc00;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n23970));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n23969));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n23968));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n23967));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n23966));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_4_lut_adj_840 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [13]), .O(n42617));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_840.LUT_INIT = 16'hdc00;
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n23557), .D(n43398));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_4_lut_adj_841 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [14]), .O(n42619));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_841.LUT_INIT = 16'hdc00;
    SB_LUT4 i15035_1_lut (.I0(n28434), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1507));
    defparam i15035_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n23557), .D(n44472));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n23557), .D(n22915));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n23557), .D(n43410));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n23557), .D(n44636));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n23557), .D(n44772));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n23557), .D(n43282));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n23557), .D(n43283));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n23557), .D(n45019));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n23557), .D(n44400));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n23557), .D(n44383));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n23557), .D(n44979));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n23557), .D(n44983));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n23557), .D(n45043));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n23557), .D(n44955));   // verilog/coms.v(125[12] 284[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n23557), .D(n44821));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n23965));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_563_9_lut (.I0(byte_transmit_counter_c[7]), .I1(byte_transmit_counter_c[7]), 
            .I2(n3839), .I3(n36967), .O(n23838)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_9_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_41_5 (.CI(n36932), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n36933));
    SB_LUT4 i1_2_lut_4_lut_adj_842 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [15]), .O(n42621));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_842.LUT_INIT = 16'hdc00;
    SB_LUT4 add_41_14_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n36941), .O(n2_adj_3130)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_843 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [16]), .O(n42623));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_843.LUT_INIT = 16'hdc00;
    SB_CARRY add_41_14 (.CI(n36941), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n36942));
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n23964));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_13_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n36940), .O(n2_adj_3131)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_844 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [17]), .O(n42625));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_844.LUT_INIT = 16'hdc00;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_3132), .S(n3));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut (.I0(n43132), .I1(n43245), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_3133));   // verilog/coms.v(147[5:27])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(n43127), .I1(n43273), .I2(n43271), .I3(n6_adj_3133), 
            .O(n22456));   // verilog/coms.v(147[5:27])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_845 (.I0(\FRAME_MATCHER.state [3]), .I1(n22456), 
            .I2(GND_net), .I3(GND_net), .O(n22334));   // verilog/coms.v(147[5:27])
    defparam i1_2_lut_adj_845.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_846 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [18]), .O(n42627));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_846.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_847 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [21]), .O(n42597));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_847.LUT_INIT = 16'hdc00;
    SB_LUT4 i2_2_lut_adj_848 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3134));
    defparam i2_2_lut_adj_848.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i7_4_lut (.I0(\data_in_frame[0] [0]), .I1(n14), .I2(n10_adj_3134), 
            .I3(\data_in_frame[0] [3]), .O(Kp_23__N_1179));
    defparam i7_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_2_lut_adj_849 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3135));   // verilog/coms.v(227[13:35])
    defparam i2_2_lut_adj_849.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_850 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_3136));   // verilog/coms.v(227[13:35])
    defparam i6_4_lut_adj_850.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_851 (.I0(\data_in_frame[0] [0]), .I1(n14_adj_3136), 
            .I2(n10_adj_3135), .I3(\data_in_frame[0] [3]), .O(n20432));   // verilog/coms.v(227[13:35])
    defparam i7_4_lut_adj_851.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_852 (.I0(n40198), .I1(n43635), .I2(n43287), .I3(n40234), 
            .O(n45002));
    defparam i3_4_lut_adj_852.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_853 (.I0(Kp_23__N_804), .I1(n43391), .I2(n43712), 
            .I3(n43518), .O(n16_adj_3137));
    defparam i6_4_lut_adj_853.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_854 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [23]), .O(n42599));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_854.LUT_INIT = 16'hdc00;
    SB_LUT4 i7_4_lut_adj_855 (.I0(\data_in_frame[16] [5]), .I1(n45002), 
            .I2(n39479), .I3(n39570), .O(n17_adj_3138));
    defparam i7_4_lut_adj_855.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[18] [1]), .I1(n17_adj_3138), .I2(n15_adj_3139), 
            .I3(n16_adj_3137), .O(n43426));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut (.I0(n43678), .I1(n43684), .I2(\data_in_frame[8] [7]), 
            .I3(\data_in_frame[6] [6]), .O(n12));   // verilog/coms.v(68[16:27])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_856 (.I0(\data_in_frame[9] [0]), .I1(n12), .I2(n43827), 
            .I3(\data_in_frame[8] [5]), .O(n44630));   // verilog/coms.v(68[16:27])
    defparam i6_4_lut_adj_856.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_857 (.I0(\data_in_frame[19] [5]), .I1(n43587), 
            .I2(n43512), .I3(\data_in_frame[17] [4]), .O(n16_adj_3140));   // verilog/coms.v(68[16:27])
    defparam i6_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_858 (.I0(n44630), .I1(n43849), .I2(\data_in_frame[17] [3]), 
            .I3(n43739), .O(n17_adj_3141));   // verilog/coms.v(68[16:27])
    defparam i7_4_lut_adj_858.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_859 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43247), .I3(\FRAME_MATCHER.i [0]), .O(n43255));
    defparam i1_2_lut_3_lut_4_lut_adj_859.LUT_INIT = 16'hf7ff;
    SB_LUT4 i1_2_lut_4_lut_adj_860 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [24]), .O(n42601));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_860.LUT_INIT = 16'hdc00;
    SB_LUT4 i9_4_lut_adj_861 (.I0(n17_adj_3141), .I1(n8_adj_3117), .I2(n16_adj_3140), 
            .I3(n22827), .O(n43789));   // verilog/coms.v(68[16:27])
    defparam i9_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_862 (.I0(\data_in_frame[19] [4]), .I1(n23346), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3142));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_862.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_863 (.I0(n43733), .I1(n43852), .I2(n22728), .I3(n6_adj_3142), 
            .O(n43614));   // verilog/coms.v(68[16:27])
    defparam i4_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[14]_c [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43885));
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_865 (.I0(n43727), .I1(\data_in_frame[5] [7]), .I2(n43508), 
            .I3(\data_in_frame[1] [5]), .O(n16_adj_3143));   // verilog/coms.v(68[16:27])
    defparam i6_4_lut_adj_865.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_866 (.I0(\data_in_frame[8] [2]), .I1(n43381), .I2(\data_in_frame[4] [0]), 
            .I3(\data_in_frame[3] [4]), .O(n17_adj_3144));   // verilog/coms.v(68[16:27])
    defparam i7_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_867 (.I0(n17_adj_3144), .I1(\data_in_frame[3] [7]), 
            .I2(n16_adj_3143), .I3(n22750), .O(n43852));   // verilog/coms.v(68[16:27])
    defparam i9_4_lut_adj_867.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_868 (.I0(n43852), .I1(n43843), .I2(n43885), .I3(n6), 
            .O(n43730));
    defparam i4_4_lut_adj_868.LUT_INIT = 16'h6996;
    SB_LUT4 i14893_2_lut_4_lut (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [29]), .O(n28291));   // verilog/coms.v(112[11:12])
    defparam i14893_2_lut_4_lut.LUT_INIT = 16'hdc00;
    SB_LUT4 i7_4_lut_adj_869 (.I0(\data_in_frame[14]_c [6]), .I1(n43490), 
            .I2(n43801), .I3(\data_in_frame[15] [1]), .O(n18));
    defparam i7_4_lut_adj_869.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_870 (.I0(\data_in_frame[17] [2]), .I1(n18), .I2(n43675), 
            .I3(n43885), .O(n20_adj_3145));
    defparam i9_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n43867), .I1(n20_adj_3145), .I2(n16_adj_3146), 
            .I3(n43739), .O(n40149));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_871 (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43843));
    defparam i1_2_lut_adj_871.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[10] [3]), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[6] [0]), .I3(GND_net), .O(n43849));   // verilog/coms.v(82[17:28])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_3147), .S(n3_adj_3148));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_3149), .S(n3_adj_3150));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_3151), .S(n3_adj_3152));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_3153), .S(n3_adj_3154));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_3155), .S(n3_adj_3156));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_3157), .S(n3_adj_3158));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_3159), .S(n3_adj_3160));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_3161), .S(n3_adj_3162));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_3163), .S(n3_adj_3164));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_3165), .S(n3_adj_3166));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_3167), .S(n3_adj_3168));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_3169), .S(n3_adj_3170));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_3171), .S(n3_adj_3172));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_3173));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3111), .S(n3_adj_3174));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3113), .S(n3_adj_3175));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3120), .S(n3_adj_3176));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3125), .S(n3_adj_3177));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3130), .S(n3_adj_3178));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3131), .S(n3_adj_3179));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3180), .S(n3_adj_3181));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3182), .S(n3_adj_3183));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3184), .S(n3_adj_3185));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3186), .S(n3_adj_3187));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3188), .S(n3_adj_3189));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3110), .S(n3_adj_3190));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3114), .S(n3_adj_3191));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3126), .S(n3_adj_3192));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3193), .S(n3_adj_3194));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3195), .S(n3_adj_3196));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16][1] ), .C(clk32MHz), 
           .D(n23963));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_872 (.I0(n23219), .I1(n40161), .I2(n40127), .I3(n40169), 
            .O(n43712));
    defparam i3_4_lut_adj_872.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_873 (.I0(n43712), .I1(\data_in_frame[14]_c [6]), 
            .I2(\data_in_frame[15] [5]), .I3(n43849), .O(n22_adj_3197));   // verilog/coms.v(82[17:28])
    defparam i9_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_adj_874 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[18] [7]), .I3(GND_net), .O(n20_adj_3198));   // verilog/coms.v(82[17:28])
    defparam i7_3_lut_adj_874.LUT_INIT = 16'h9696;
    SB_CARRY add_41_13 (.CI(n36940), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n36941));
    SB_LUT4 add_563_8_lut (.I0(byte_transmit_counter_c[6]), .I1(byte_transmit_counter_c[6]), 
            .I2(n3839), .I3(n36966), .O(n23835)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_8_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_41_12_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n36939), .O(n2_adj_3180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_563_8 (.CI(n36966), .I0(byte_transmit_counter_c[6]), .I1(n3839), 
            .CO(n36967));
    SB_LUT4 add_563_7_lut (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[5]), 
            .I2(n3839), .I3(n36965), .O(n23832)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_563_7 (.CI(n36965), .I0(byte_transmit_counter_c[5]), .I1(n3839), 
            .CO(n36966));
    SB_LUT4 add_41_4_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n36931), .O(n2_adj_3193)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_563_6_lut (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter_c[4]), 
            .I2(n3839), .I3(n36964), .O(n23829)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_6_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_4_lut_adj_875 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [30]), .O(n42603));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_875.LUT_INIT = 16'hdc00;
    SB_CARRY add_41_4 (.CI(n36931), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n36932));
    SB_CARRY add_41_12 (.CI(n36939), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n36940));
    SB_LUT4 add_41_3_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n36930), .O(n2_adj_3195)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_563_6 (.CI(n36964), .I0(byte_transmit_counter_c[4]), .I1(n3839), 
            .CO(n36965));
    SB_LUT4 i11_4_lut_adj_876 (.I0(n22728), .I1(n22_adj_3197), .I2(n16_adj_3199), 
            .I3(n43843), .O(n24_adj_3200));   // verilog/coms.v(82[17:28])
    defparam i11_4_lut_adj_876.LUT_INIT = 16'h6996;
    SB_LUT4 add_563_5_lut (.I0(byte_transmit_counter_c[3]), .I1(byte_transmit_counter_c[3]), 
            .I2(n3839), .I3(n36963), .O(n23826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_5_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_41_11_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n36938), .O(n2_adj_3182)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_11_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n24307));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n23962));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n23961));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n23960));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n23959));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i12_4_lut_adj_877 (.I0(n43724), .I1(n24_adj_3200), .I2(n20_adj_3198), 
            .I3(\data_in_frame[6] [1]), .O(n43501));   // verilog/coms.v(82[17:28])
    defparam i12_4_lut_adj_877.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_878 (.I0(n43501), .I1(n23078), .I2(n43528), .I3(GND_net), 
            .O(n8_adj_3201));
    defparam i2_3_lut_adj_878.LUT_INIT = 16'h9696;
    SB_CARRY add_563_5 (.CI(n36963), .I0(byte_transmit_counter_c[3]), .I1(n3839), 
            .CO(n36964));
    SB_LUT4 add_563_4_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[2]), 
            .I2(n3839), .I3(n36962), .O(n23823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_4_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i4_4_lut_adj_879 (.I0(\data_in_frame[19] [3]), .I1(n8_adj_3201), 
            .I2(n40149), .I3(n43730), .O(n10_adj_3202));
    defparam i4_4_lut_adj_879.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n23958));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i5_4_lut_adj_880 (.I0(n43614), .I1(n10_adj_3202), .I2(n43278), 
            .I3(n43789), .O(n23212));
    defparam i5_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_881 (.I0(n22442), .I1(n2_adj_3124), .I2(n20099), 
            .I3(\FRAME_MATCHER.state_c [31]), .O(n7_adj_3127));   // verilog/coms.v(112[11:12])
    defparam i1_2_lut_4_lut_adj_881.LUT_INIT = 16'hdc00;
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n23957));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n23956));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n23955));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_882 (.I0(\data_in_frame[19] [0]), .I1(n43471), 
            .I2(n40163), .I3(\data_in_frame[16] [6]), .O(n23169));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_882.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n23954));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n23953));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_883 (.I0(n43557), .I1(\data_in_frame[6] [4]), .I2(n10_adj_3116), 
            .I3(n22796), .O(n22827));   // verilog/coms.v(71[16:43])
    defparam i3_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_CARRY add_563_4 (.CI(n36962), .I0(byte_transmit_counter_c[2]), .I1(n3839), 
            .CO(n36963));
    SB_LUT4 add_563_3_lut (.I0(byte_transmit_counter_c[1]), .I1(byte_transmit_counter_c[1]), 
            .I2(n3839), .I3(n36961), .O(n23820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43675));
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_885 (.I0(n23176), .I1(n43367), .I2(GND_net), 
            .I3(GND_net), .O(n43827));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i34441_2_lut_3_lut (.I0(r_SM_Main_2__N_2747[0]), .I1(tx_active), 
            .I2(n7_adj_3203), .I3(GND_net), .O(tx_transmit_N_2639));   // verilog/coms.v(125[12] 284[6])
    defparam i34441_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i4_4_lut_adj_886 (.I0(n8_adj_3117), .I1(\data_in_frame[8] [3]), 
            .I2(n43827), .I3(n43675), .O(n10_adj_3204));   // verilog/coms.v(70[16:42])
    defparam i4_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_CARRY add_563_3 (.CI(n36961), .I0(byte_transmit_counter_c[1]), .I1(n3839), 
            .CO(n36962));
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[6] [2]), .I1(n10_adj_3204), .I2(\data_in_frame[6] [3]), 
            .I3(GND_net), .O(n22750));   // verilog/coms.v(70[16:42])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 add_563_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_2639), .I3(GND_net), .O(n2241)) /* synthesis syn_instantiated=1 */ ;
    defparam add_563_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_887 (.I0(\data_in_frame[12] [7]), .I1(n22827), 
            .I2(GND_net), .I3(GND_net), .O(n43569));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_888 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[10] [7]), 
            .I2(n43569), .I3(n22750), .O(n43587));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n23952));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n23951));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n23950));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n23949));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18][0] ), .C(clk32MHz), 
           .D(n23948));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n23947));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18][2] ), .C(clk32MHz), 
           .D(n23946));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n23945));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i3_4_lut_adj_889 (.I0(\data_in_frame[8] [7]), .I1(n43343), .I2(\data_in_frame[8] [6]), 
            .I3(n10_adj_3116), .O(n23209));   // verilog/coms.v(71[16:43])
    defparam i3_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n23944));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n23943));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n23942));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n23941));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_adj_890 (.I0(Kp_23__N_865), .I1(n43441), .I2(n23209), 
            .I3(GND_net), .O(n43879));
    defparam i2_3_lut_adj_890.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n23940));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n23939));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n23938));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34523 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter_c[1]), .O(n50029));
    defparam byte_transmit_counter_0__bdd_4_lut_34523.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_891 (.I0(r_SM_Main_2__N_2747[0]), .I1(tx_active), 
            .I2(n7_adj_3203), .I3(GND_net), .O(n744));   // verilog/coms.v(125[12] 284[6])
    defparam i1_2_lut_3_lut_adj_891.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_adj_892 (.I0(n43873), .I1(n43879), .I2(\data_in_frame[16] [5]), 
            .I3(GND_net), .O(n43706));
    defparam i2_3_lut_adj_892.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_893 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [2]), 
            .I2(\data_in_frame[16][1] ), .I3(\data_in_frame[16] [3]), .O(n23219));   // verilog/coms.v(82[17:63])
    defparam i3_4_lut_adj_893.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n103), .I1(n4_c), .I2(n737), .I3(n22443), 
            .O(n44574));   // verilog/coms.v(92[12:19])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_3_lut_adj_894 (.I0(n103), .I1(n4_c), .I2(n2854), 
            .I3(GND_net), .O(n20098));   // verilog/coms.v(92[12:19])
    defparam i1_2_lut_3_lut_adj_894.LUT_INIT = 16'h0202;
    SB_CARRY add_563_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_2639), 
            .CO(n36961));
    SB_LUT4 i1_2_lut_3_lut_adj_895 (.I0(n103), .I1(n4_c), .I2(n3758), 
            .I3(GND_net), .O(n20099));   // verilog/coms.v(92[12:19])
    defparam i1_2_lut_3_lut_adj_895.LUT_INIT = 16'h0202;
    SB_LUT4 i3_4_lut_adj_896 (.I0(n43833), .I1(n43802), .I2(n23219), .I3(n43518), 
            .O(n43873));
    defparam i3_4_lut_adj_896.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_4_lut (.I0(n139), .I1(n43263), .I2(\data_in[0] [6]), 
            .I3(\data_in[3] [0]), .O(n8_adj_3205));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_adj_897 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43733));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h6666;
    SB_LUT4 add_41_33_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n36960), .O(n2_adj_3132)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_33_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n23937));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_32_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n36959), .O(n2_adj_3147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_32_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n23936));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n23935));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n23934));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n23933));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n23932));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n23931));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n23930));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n23929));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n23928));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_32 (.CI(n36959), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n36960));
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n23927));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_31_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n36958), .O(n2_adj_3149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_898 (.I0(n43301), .I1(n23242), .I2(\data_in_frame[12] [4]), 
            .I3(n43644), .O(n10_adj_3206));   // verilog/coms.v(225[9:81])
    defparam i4_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_899 (.I0(\data_in_frame[10] [3]), .I1(n10_adj_3206), 
            .I2(\data_in_frame[8] [0]), .I3(GND_net), .O(n22728));   // verilog/coms.v(225[9:81])
    defparam i5_3_lut_adj_899.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_900 (.I0(Kp_23__N_458), .I1(\data_in_frame[10] [1]), 
            .I2(n22928), .I3(\data_in_frame[8] [0]), .O(n12_adj_3207));   // verilog/coms.v(82[17:28])
    defparam i5_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_CARRY add_41_11 (.CI(n36938), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n36939));
    SB_LUT4 n50029_bdd_4_lut (.I0(n50029), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter_c[1]), 
            .O(n50032));
    defparam n50029_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_901 (.I0(Kp_23__N_515), .I1(n12_adj_3207), .I2(\data_in_frame[5] [6]), 
            .I3(n43894), .O(n43751));   // verilog/coms.v(82[17:28])
    defparam i6_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_902 (.I0(\data_in_frame[14]_c [5]), .I1(n22728), 
            .I2(GND_net), .I3(GND_net), .O(n43518));
    defparam i1_2_lut_adj_902.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_903 (.I0(\data_in_frame[9] [7]), .I1(n43754), .I2(\data_in_frame[7] [6]), 
            .I3(GND_net), .O(n43855));
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_904 (.I0(n139), .I1(n43263), .I2(n10_adj_3208), 
            .I3(GND_net), .O(n103));
    defparam i1_2_lut_3_lut_adj_904.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_905 (.I0(n40131), .I1(n16), .I2(\data_in_frame[4] [6]), 
            .I3(n43462), .O(n10_adj_3209));
    defparam i4_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_906 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[7] [3]), 
            .I2(n10_adj_3209), .I3(Kp_23__N_325), .O(n43474));
    defparam i1_4_lut_adj_906.LUT_INIT = 16'h9669;
    SB_LUT4 i29725_3_lut_4_lut (.I0(n22443), .I1(n737), .I2(n2854), .I3(n22454), 
            .O(n45225));
    defparam i29725_3_lut_4_lut.LUT_INIT = 16'heee0;
    SB_LUT4 i1_2_lut_adj_907 (.I0(n39443), .I1(n43474), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3210));
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_908 (.I0(n43391), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[14]_c [2]), .I3(n6_adj_3210), .O(n39561));
    defparam i4_4_lut_adj_908.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_909 (.I0(n22443), .I1(n737), .I2(n122), 
            .I3(n103), .O(n44586));
    defparam i2_3_lut_4_lut_adj_909.LUT_INIT = 16'h1000;
    SB_LUT4 i2_3_lut_4_lut_adj_910 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n28284), .O(n43235));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_910.LUT_INIT = 16'hefff;
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n23926));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n23925));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n23924));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n23923));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n23922));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n23921));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n23920));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n23919));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n23918));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_10_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n36937), .O(n2_adj_3184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_31 (.CI(n36958), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n36959));
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n23917));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n23916));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n23915));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n23914));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_3 (.CI(n36930), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n36931));
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n23913));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_10 (.CI(n36937), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n36938));
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n23912));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n23911));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n23910));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i1 (.Q(\PWMLimit[1] ), .C(clk32MHz), .D(n23909));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i2 (.Q(\PWMLimit[2] ), .C(clk32MHz), .D(n23908));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i3 (.Q(\PWMLimit[3] ), .C(clk32MHz), .D(n23907));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i4 (.Q(\PWMLimit[4] ), .C(clk32MHz), .D(n23906));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i5 (.Q(\PWMLimit[5] ), .C(clk32MHz), .D(n23905));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i6 (.Q(\PWMLimit[6] ), .C(clk32MHz), .D(n28060));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_30_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n36957), .O(n2_adj_3151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_30_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i7 (.Q(\PWMLimit[7] ), .C(clk32MHz), .D(n23903));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i8 (.Q(\PWMLimit[8] ), .C(clk32MHz), .D(n23902));   // verilog/coms.v(125[12] 284[6])
    SB_DFF PWMLimit_i0_i9 (.Q(\PWMLimit[9] ), .C(clk32MHz), .D(n23901));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_30 (.CI(n36957), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n36958));
    SB_LUT4 i2_3_lut_4_lut_adj_911 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n22501), .I3(\FRAME_MATCHER.i [4]), .O(n22343));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_911.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_912 (.I0(n43563), .I1(n43538), .I2(\data_in_frame[9] [4]), 
            .I3(n43770), .O(n10_adj_3211));
    defparam i4_4_lut_adj_912.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_913 (.I0(n23183), .I1(n10_adj_3211), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n40129));
    defparam i5_3_lut_adj_913.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_914 (.I0(n2_adj_3124), .I1(n42), .I2(\FRAME_MATCHER.state_c [4]), 
            .I3(GND_net), .O(n42675));
    defparam i1_2_lut_3_lut_adj_914.LUT_INIT = 16'he0e0;
    SB_LUT4 add_41_29_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n36956), .O(n2_adj_3153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_29 (.CI(n36956), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n36957));
    SB_LUT4 i1_2_lut_3_lut_adj_915 (.I0(n2_adj_3124), .I1(n42), .I2(\FRAME_MATCHER.state_c [19]), 
            .I3(GND_net), .O(n42677));
    defparam i1_2_lut_3_lut_adj_915.LUT_INIT = 16'he0e0;
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n50101));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10606_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n24021));
    defparam i10606_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_916 (.I0(n2_adj_3124), .I1(n42), .I2(\FRAME_MATCHER.state_c [20]), 
            .I3(GND_net), .O(n42681));
    defparam i1_2_lut_3_lut_adj_916.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_917 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(n6_adj_3213), .O(n23242));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_28_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n36955), .O(n2_adj_3155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_28 (.CI(n36955), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n36956));
    SB_LUT4 add_41_27_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n36954), .O(n2_adj_3157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_27 (.CI(n36954), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n36955));
    SB_LUT4 add_41_26_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n36953), .O(n2_adj_3159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_918 (.I0(n2_adj_3124), .I1(n42), .I2(\FRAME_MATCHER.state_c [25]), 
            .I3(GND_net), .O(n7_adj_3128));
    defparam i1_2_lut_3_lut_adj_918.LUT_INIT = 16'he0e0;
    SB_CARRY add_41_26 (.CI(n36953), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n36954));
    SB_LUT4 i1_2_lut_3_lut_adj_919 (.I0(n2_adj_3124), .I1(n42), .I2(\FRAME_MATCHER.state_c [26]), 
            .I3(GND_net), .O(n42661));
    defparam i1_2_lut_3_lut_adj_919.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43352));
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_921 (.I0(\data_in_frame[9] [6]), .I1(n43352), .I2(n23242), 
            .I3(n22928), .O(n39443));
    defparam i3_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_922 (.I0(n2_adj_3124), .I1(n42), .I2(\FRAME_MATCHER.state_c [27]), 
            .I3(GND_net), .O(n42663));
    defparam i1_2_lut_3_lut_adj_922.LUT_INIT = 16'he0e0;
    SB_LUT4 i3_4_lut_adj_923 (.I0(n39500), .I1(n43635), .I2(n43308), .I3(n39443), 
            .O(n39570));
    defparam i3_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i14892_2_lut_3_lut (.I0(n2_adj_3124), .I1(n42), .I2(\FRAME_MATCHER.state_c [28]), 
            .I3(GND_net), .O(n28289));
    defparam i14892_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_924 (.I0(n22454), .I1(n20125), .I2(n2_adj_3124), 
            .I3(n37), .O(n44497));   // verilog/coms.v(112[11:12])
    defparam i2_3_lut_4_lut_adj_924.LUT_INIT = 16'hfff4;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_925 (.I0(n22454), .I1(n20125), .I2(n37), 
            .I3(n54), .O(n44479));   // verilog/coms.v(112[11:12])
    defparam i2_2_lut_3_lut_4_lut_adj_925.LUT_INIT = 16'hfff4;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_in_frame[14][0] ), .I1(n39570), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3214));
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i10607_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n24022));
    defparam i10607_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15295_3_lut_4_lut (.I0(n54), .I1(n37), .I2(n59), .I3(\FRAME_MATCHER.state_c [7]), 
            .O(n28698));
    defparam i15295_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i4_4_lut_adj_927 (.I0(n43596), .I1(n40198), .I2(n40137), .I3(n6_adj_3214), 
            .O(n39479));
    defparam i4_4_lut_adj_927.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_928 (.I0(n39479), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43718));
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_929 (.I0(\data_in_frame[16] [4]), .I1(n39561), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3215));
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_930 (.I0(n43855), .I1(n43751), .I2(n43888), .I3(n6_adj_3215), 
            .O(n43471));
    defparam i4_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter_c[5]), .C(clk32MHz), 
           .D(n23834));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter_c[6]), .C(clk32MHz), 
           .D(n23837));   // verilog/coms.v(125[12] 284[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter_c[7]), .C(clk32MHz), 
           .D(n23840));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n24289));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10608_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n24023));
    defparam i10608_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_931 (.I0(n43471), .I1(\data_in_frame[18] [5]), 
            .I2(n43718), .I3(\data_in_frame[18] [4]), .O(n43453));   // verilog/coms.v(82[17:63])
    defparam i2_4_lut_adj_931.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_932 (.I0(n39570), .I1(n39561), .I2(\data_in_frame[16] [3]), 
            .I3(GND_net), .O(n22605));
    defparam i2_3_lut_adj_932.LUT_INIT = 16'h9696;
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n24288));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_4_lut_adj_933 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(n43477), .I3(n23251), .O(n39281));
    defparam i2_3_lut_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43441));
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n24287));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1][6] ), .C(clk32MHz), .D(n24240));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34518 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter_c[1]), .O(n50023));
    defparam byte_transmit_counter_0__bdd_4_lut_34518.LUT_INIT = 16'he4aa;
    SB_LUT4 n50023_bdd_4_lut (.I0(n50023), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter_c[1]), 
            .O(n50026));
    defparam n50023_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n24239));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSR tx_transmit_3220 (.Q(r_SM_Main_2__N_2747[0]), .C(clk32MHz), 
            .D(n2416[0]), .R(n44089));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 add_41_25_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n36952), .O(n2_adj_3161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_935 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n43703));
    defparam i1_2_lut_3_lut_adj_935.LUT_INIT = 16'h9696;
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n24286));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_4_lut_adj_936 (.I0(n23254), .I1(n10_adj_3216), .I2(\data_out_frame[16] [2]), 
            .I3(\data_out_frame[20] [4]), .O(n39470));
    defparam i1_2_lut_4_lut_adj_936.LUT_INIT = 16'h9669;
    SB_DFF data_in_0___i17 (.Q(\data_in[2]_c [0]), .C(clk32MHz), .D(n24238));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_2_lut_4_lut (.I0(n23254), .I1(n10_adj_3216), .I2(\data_out_frame[16] [2]), 
            .I3(n43397), .O(n10_adj_3217));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_937 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[12] [5]), 
            .I2(n22721), .I3(GND_net), .O(n43724));   // verilog/coms.v(82[17:28])
    defparam i2_3_lut_adj_937.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i18 (.Q(\data_in[2][1] ), .C(clk32MHz), .D(n27276));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n24285));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_adj_938 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43462));
    defparam i1_2_lut_adj_938.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_939 (.I0(\data_in_frame[10] [5]), .I1(n43724), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[15] [1]), .O(n43512));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n24320));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n24319));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n24318));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n24317));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_adj_940 (.I0(\data_in_frame[4] [5]), .I1(n5_adj_3218), 
            .I2(n4_adj_3219), .I3(GND_net), .O(n23183));   // verilog/coms.v(225[9:81])
    defparam i2_3_lut_adj_940.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_941 (.I0(n23183), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43684));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_942 (.I0(\data_in_frame[8] [5]), .I1(\data_in_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43557));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_adj_942.LUT_INIT = 16'h6666;
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n24284));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i5_4_lut_adj_943 (.I0(n43557), .I1(n43684), .I2(n23176), .I3(\data_in_frame[9] [1]), 
            .O(n12_adj_3220));   // verilog/coms.v(71[16:43])
    defparam i5_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i10609_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n24024));
    defparam i10609_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Kd_i1 (.Q(\Kd[1] ), .C(clk32MHz), .D(n24283));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_4_lut_adj_944 (.I0(\data_out_frame[11] [0]), .I1(n43837), 
            .I2(n22771), .I3(\data_out_frame[12] [6]), .O(n43767));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_DFF Kd_i2 (.Q(\Kd[2] ), .C(clk32MHz), .D(n24282));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i3 (.Q(\Kd[3] ), .C(clk32MHz), .D(n24281));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_3_lut_adj_945 (.I0(\data_out_frame[11] [0]), .I1(n43837), 
            .I2(\data_out_frame[6] [6]), .I3(GND_net), .O(n6_adj_3221));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_945.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n24306));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i6_4_lut_adj_946 (.I0(\data_in_frame[13] [3]), .I1(n12_adj_3220), 
            .I2(n43830), .I3(\data_in_frame[10] [7]), .O(n43343));   // verilog/coms.v(71[16:43])
    defparam i6_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_947 (.I0(\data_in_frame[14]_c [1]), .I1(\data_in_frame[12] [0]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n43308));
    defparam i2_3_lut_adj_947.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_948 (.I0(\data_in_frame[14][0] ), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43287));
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_949 (.I0(\data_in_frame[10][6] ), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43821));   // verilog/coms.v(69[16:41])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_950 (.I0(\data_in_frame[14]_c [6]), .I1(\data_in_frame[12] [6]), 
            .I2(\data_in_frame[14]_c [7]), .I3(\data_in_frame[15] [0]), 
            .O(n43508));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_951 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(n43566), .I3(GND_net), .O(n22928));
    defparam i1_3_lut_adj_951.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_952 (.I0(n22928), .I1(n23385), .I2(GND_net), 
            .I3(GND_net), .O(n40131));
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_in_frame[9] [6]), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43894));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_954 (.I0(n22953), .I1(\data_in_frame[7] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n43748));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_16__7__I_0_3242_2_lut (.I0(\data_in_frame[16] [7]), 
            .I1(\data_in_frame[16] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_804));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_16__7__I_0_3242_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i18_4_lut (.I0(\data_in_frame[13] [0]), .I1(n43748), .I2(n43459), 
            .I3(\data_in_frame[10] [2]), .O(n52));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10610_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n24025));
    defparam i10610_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_955 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n6_adj_3222));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_955.LUT_INIT = 16'h9696;
    SB_LUT4 i25_4_lut (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[9] [5]), 
            .I2(n22953), .I3(\data_in_frame[12] [1]), .O(n59_adj_3223));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(\data_in_frame[14]_c [3]), .I1(n43858), .I2(n43894), 
            .I3(n43770), .O(n56));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_956 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[7] [7]), .O(n43375));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_in_frame[15] [5]), .I1(n43678), .I2(n43804), 
            .I3(n43508), .O(n54_adj_3224));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n43343), .I1(\data_in_frame[11] [6]), .I2(\data_in_frame[8] [4]), 
            .I3(\data_in_frame[10] [0]), .O(n55));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n43870), .I1(n43299), .I2(n43596), .I3(\data_in_frame[7] [6]), 
            .O(n53));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n43388), .I1(n43287), .I2(n43308), .I3(\data_in_frame[14] [4]), 
            .O(n58));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n59_adj_3223), .I1(\data_in_frame[14]_c [2]), 
            .I2(n52), .I3(\data_in_frame[15] [3]), .O(n64));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n43727), .I1(n43512), .I2(n43626), .I3(n43462), 
            .O(n57));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n53), .I1(n55), .I2(n54_adj_3224), .I3(n56), 
            .O(n65));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut (.I0(n65), .I1(n57), .I2(n64), .I3(n58), .O(n40127));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_in_frame[14]_c [3]), .I1(\data_in_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43888));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\data_in_frame[7] [3]), .I1(n39466), .I2(GND_net), 
            .I3(GND_net), .O(n43538));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_4_lut_adj_959 (.I0(n22771), .I1(n43783), .I2(\data_out_frame[12] [6]), 
            .I3(n10_adj_3225), .O(n23436));
    defparam i5_3_lut_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i10611_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n24026));
    defparam i10611_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_960 (.I0(\data_in_frame[5] [5]), .I1(n43742), .I2(n43525), 
            .I3(\data_in_frame[1] [3]), .O(n22721));   // verilog/coms.v(70[16:34])
    defparam i3_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_961 (.I0(n43541), .I1(\data_in_frame[3] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3226));   // verilog/coms.v(82[17:28])
    defparam i2_2_lut_adj_961.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_962 (.I0(\data_in_frame[5] [3]), .I1(n21061), .I2(n6_adj_3226), 
            .I3(\data_in_frame[3] [2]), .O(n22953));
    defparam i1_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_DFF Kd_i4 (.Q(\Kd[4] ), .C(clk32MHz), .D(n24280));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i2_3_lut_adj_963 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[10] [1]), 
            .I2(n22953), .I3(GND_net), .O(n43867));
    defparam i2_3_lut_adj_963.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_964 (.I0(\data_in_frame[1] [3]), .I1(n43429), .I2(\data_in_frame[3] [6]), 
            .I3(\data_in_frame[5] [7]), .O(n8_adj_3117));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_965 (.I0(n43355), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[6] [1]), .O(n43861));
    defparam i1_2_lut_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_966 (.I0(n43355), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[5] [7]), .I3(n22746), .O(n43694));
    defparam i1_2_lut_4_lut_adj_966.LUT_INIT = 16'h6996;
    SB_LUT4 i10542_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n23957));
    defparam i10542_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_41_25 (.CI(n36952), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n36953));
    SB_LUT4 add_41_9_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n36936), .O(n2_adj_3186)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10612_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n24027));
    defparam i10612_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_967 (.I0(n8_adj_3117), .I1(n43867), .I2(\data_in_frame[8] [1]), 
            .I3(GND_net), .O(n43641));
    defparam i2_3_lut_adj_967.LUT_INIT = 16'h9696;
    SB_LUT4 add_41_24_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n36951), .O(n2_adj_3163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_24 (.CI(n36951), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n36952));
    SB_LUT4 add_41_23_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n36950), .O(n2_adj_3165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_23_lut.LUT_INIT = 16'h8228;
    SB_DFF Kd_i5 (.Q(\Kd[5] ), .C(clk32MHz), .D(n24279));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Kd_i6 (.Q(\Kd[6] ), .C(clk32MHz), .D(n24278));   // verilog/coms.v(125[12] 284[6])
    SB_CARRY add_41_23 (.CI(n36950), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n36951));
    SB_DFF Kd_i7 (.Q(\Kd[7] ), .C(clk32MHz), .D(n24277));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i1_2_lut_adj_968 (.I0(\data_in_frame[10] [2]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43882));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_969 (.I0(n40127), .I1(Kp_23__N_804), .I2(GND_net), 
            .I3(GND_net), .O(n43833));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_DFF deadband_i0_i0 (.Q(\deadband[0] ), .C(clk32MHz), .D(n23757));   // verilog/coms.v(125[12] 284[6])
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n23756));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n24203));   // verilog/coms.v(125[12] 284[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3227), .S(n3_adj_3228));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_34553 (.I0(byte_transmit_counter_c[1]), 
            .I1(n11), .I2(n12_adj_3229), .I3(byte_transmit_counter_c[2]), 
            .O(n50011));
    defparam byte_transmit_counter_1__bdd_4_lut_34553.LUT_INIT = 16'he4aa;
    SB_LUT4 i10543_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n23958));
    defparam i10543_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n24316));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n24315));   // verilog/coms.v(125[12] 284[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
           .D(n42561));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i10544_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n23959));
    defparam i10544_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n24314));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n24313));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i5_4_lut_adj_970 (.I0(n43754), .I1(n43846), .I2(\data_in_frame[7] [4]), 
            .I3(n43641), .O(n12_adj_3230));
    defparam i5_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i0 (.Q(\PWMLimit[0] ), .C(clk32MHz), .D(n23742));   // verilog/coms.v(125[12] 284[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n23741));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n23740));   // verilog/coms.v(125[12] 284[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0]_c [0]), .C(clk32MHz), .D(n23739));   // verilog/coms.v(125[12] 284[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n23738));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 i6_4_lut_adj_971 (.I0(\data_in_frame[7] [7]), .I1(n12_adj_3230), 
            .I2(n43882), .I3(\data_in_frame[10] [0]), .O(n40169));
    defparam i6_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_DFF Kd_i0 (.Q(\Kd[0] ), .C(clk32MHz), .D(n23737));   // verilog/coms.v(125[12] 284[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n23736));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 data_in_frame_18__7__I_0_3244_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_785));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_18__7__I_0_3244_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_972 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43349));   // verilog/coms.v(67[16:27])
    defparam i1_2_lut_adj_972.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_973 (.I0(n40169), .I1(n43691), .I2(\data_in_frame[17] [1]), 
            .I3(n43833), .O(n26));
    defparam i11_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n23735));   // verilog/coms.v(125[12] 284[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n23734));   // verilog/coms.v(125[12] 284[6])
    SB_LUT4 n50011_bdd_4_lut (.I0(n50011), .I1(n9), .I2(n8_adj_3231), 
            .I3(byte_transmit_counter_c[2]), .O(n50014));
    defparam n50011_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10613_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43247), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n24028));
    defparam i10613_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_974 (.I0(Kp_23__N_785), .I1(\data_in_frame[16] [0]), 
            .I2(\data_in_frame[18] [1]), .I3(n43349), .O(n24_adj_3232));
    defparam i9_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_975 (.I0(n43733), .I1(n43873), .I2(\data_in_frame[17] [0]), 
            .I3(n43593), .O(n25));
    defparam i10_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_LUT4 i10545_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n23960));
    defparam i10545_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut (.I0(\data_in_frame[18] [3]), .I1(n40163), .I2(n22605), 
            .I3(n43453), .O(n23));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_22_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n36949), .O(n2_adj_3167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_41_2_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2_adj_3227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_22 (.CI(n36949), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n36950));
    SB_CARRY add_41_9 (.CI(n36936), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n36937));
    SB_LUT4 add_41_21_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n36948), .O(n2_adj_3169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n36930));
    SB_LUT4 add_41_8_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n36935), .O(n2_adj_3188)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_41_21 (.CI(n36948), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n36949));
    SB_LUT4 i14_4_lut (.I0(n23), .I1(n25), .I2(n24_adj_3232), .I3(n26), 
            .O(n40194));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_41_20_lut (.I0(n1507), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n36947), .O(n2_adj_3171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_41_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_976 (.I0(n43706), .I1(n40234), .I2(\data_in_frame[18][0] ), 
            .I3(\data_in_frame[17] [5]), .O(n8_adj_3233));
    defparam i1_4_lut_adj_976.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_977 (.I0(n43671), .I1(n43824), .I2(\data_in_frame[15] [6]), 
            .I3(n43587), .O(n12_adj_3234));
    defparam i5_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_978 (.I0(\data_in_frame[19] [7]), .I1(n40194), 
            .I2(n12_adj_3234), .I3(n8_adj_3233), .O(n43278));
    defparam i1_4_lut_adj_978.LUT_INIT = 16'h9669;
    SB_LUT4 i10598_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n24013));
    defparam i10598_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_979 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[1] [0]), .O(n43541));   // verilog/coms.v(68[16:69])
    defparam i3_4_lut_adj_979.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_980 (.I0(n43541), .I1(\data_in_frame[5] [1]), .I2(n43415), 
            .I3(GND_net), .O(n39466));
    defparam i2_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i10546_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n23961));
    defparam i10546_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\data_in_frame[9] [3]), .I1(\data_in_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43626));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_982 (.I0(\data_in_frame[6] [7]), .I1(n43626), .I2(n39466), 
            .I3(\data_in_frame[7] [0]), .O(n12_adj_3236));
    defparam i5_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_983 (.I0(n23385), .I1(n12_adj_3236), .I2(n43795), 
            .I3(\data_in_frame[7] [2]), .O(n40137));
    defparam i6_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_984 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[6] [0]), .I3(GND_net), .O(n43371));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_984.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_985 (.I0(\data_in_frame[8] [2]), .I1(n23367), .I2(\data_in_frame[6] [1]), 
            .I3(GND_net), .O(n43644));   // verilog/coms.v(225[9:81])
    defparam i2_3_lut_adj_985.LUT_INIT = 16'h9696;
    SB_LUT4 i10547_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n23962));
    defparam i10547_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_986 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1][4] ), .O(Kp_23__N_458));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i10599_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n24014));
    defparam i10599_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_987 (.I0(Kp_23__N_458), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43804));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_987.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_988 (.I0(n22801), .I1(n43544), .I2(\data_in_frame[13] [1]), 
            .I3(GND_net), .O(n43824));
    defparam i2_3_lut_adj_988.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_989 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[11] [0]), 
            .I2(n43644), .I3(GND_net), .O(n14_adj_3237));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_989.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_990 (.I0(n43824), .I1(n43804), .I2(n22), .I3(\data_in_frame[12] [6]), 
            .O(n15_adj_3239));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_991 (.I0(n15_adj_3239), .I1(\data_in_frame[10] [5]), 
            .I2(n14_adj_3237), .I3(n43371), .O(n23346));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_992 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43593));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_993 (.I0(\data_in_frame[1] [6]), .I1(n43423), .I2(\data_in_frame[4] [2]), 
            .I3(GND_net), .O(n23176));   // verilog/coms.v(67[16:27])
    defparam i2_3_lut_adj_993.LUT_INIT = 16'h9696;
    SB_LUT4 i10548_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[1]), 
            .I3(\data_in_frame[16][1] ), .O(n23963));
    defparam i10548_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_994 (.I0(\data_in_frame[4] [6]), .I1(\data_in_frame[7] [0]), 
            .I2(\data_in_frame[11] [2]), .I3(n6_adj_3240), .O(n43830));   // verilog/coms.v(71[16:43])
    defparam i4_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43758));   // verilog/coms.v(75[16:50])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_996 (.I0(n23358), .I1(n43415), .I2(n23468), .I3(GND_net), 
            .O(Kp_23__N_328));
    defparam i2_3_lut_adj_996.LUT_INIT = 16'h9696;
    SB_LUT4 i10549_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43235), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n23964));
    defparam i10549_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_997 (.I0(n22796), .I1(\data_in_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43858));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_998 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43429));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_998.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_999 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43525));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1000 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43742));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43495));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h6666;
    SB_LUT4 i10534_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n23949));
    defparam i10534_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1002 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n43423));   // verilog/coms.v(67[16:27])
    defparam i2_3_lut_adj_1002.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1003 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [5]), .I3(GND_net), .O(n23358));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1003.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1004 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n5_adj_3218));   // verilog/coms.v(161[9:87])
    defparam i2_3_lut_adj_1004.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(n5_adj_3218), .I1(n23358), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_325));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1006 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(GND_net), .O(n43381));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1006.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43480));   // verilog/coms.v(68[16:69])
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i10535_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n23950));
    defparam i10535_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1008 (.I0(n23468), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[0] [4]), .O(n43566));   // verilog/coms.v(73[16:27])
    defparam i3_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(Kp_23__N_325), .I1(n43480), .I2(\data_in_frame[2] [6]), 
            .I3(n18_adj_3241), .O(n30));   // verilog/coms.v(75[16:27])
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10536_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n23951));
    defparam i10536_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i11_4_lut_adj_1009 (.I0(n43378), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[0] [3]), .I3(n43495), .O(n28));   // verilog/coms.v(75[16:27])
    defparam i11_4_lut_adj_1009.LUT_INIT = 16'h6996;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(148[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut_adj_1010 (.I0(\data_in_frame[0] [5]), .I1(n43655), 
            .I2(n43780), .I3(n43423), .O(n29));   // verilog/coms.v(75[16:27])
    defparam i12_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1011 (.I0(n43394), .I1(\data_in_frame[3] [1]), 
            .I2(n43525), .I3(n43429), .O(n27));   // verilog/coms.v(75[16:27])
    defparam i10_4_lut_adj_1011.LUT_INIT = 16'h6996;
    SB_LUT4 i10537_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n23952));
    defparam i10537_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10538_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n23953));
    defparam i10538_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30), .O(n43415));   // verilog/coms.v(75[16:27])
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10600_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n24015));
    defparam i10600_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34513 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter_c[1]), .O(n50005));
    defparam byte_transmit_counter_0__bdd_4_lut_34513.LUT_INIT = 16'he4aa;
    SB_LUT4 i10539_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n23954));
    defparam i10539_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(\data_in_frame[7] [1]), .I1(\data_in_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43563));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1013 (.I0(n43415), .I1(n43566), .I2(\data_in_frame[5] [0]), 
            .I3(GND_net), .O(n23385));
    defparam i2_3_lut_adj_1013.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1014 (.I0(n43858), .I1(\data_in_frame[9] [2]), 
            .I2(Kp_23__N_328), .I3(n43758), .O(n15_adj_3242));
    defparam i6_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1015 (.I0(n15_adj_3242), .I1(\data_in_frame[4] [7]), 
            .I2(n14_adj_3243), .I3(\data_in_frame[6] [5]), .O(n23202));
    defparam i8_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1016 (.I0(\data_in_frame[9] [0]), .I1(n43830), 
            .I2(n43758), .I3(n43544), .O(n22833));   // verilog/coms.v(75[16:50])
    defparam i3_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(n22833), .I1(n23202), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_865));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1018 (.I0(n23202), .I1(n40137), .I2(\data_in_frame[11] [4]), 
            .I3(GND_net), .O(n40155));
    defparam i2_3_lut_adj_1018.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1019 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[2] [3]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n4_adj_3219));   // verilog/coms.v(161[9:87])
    defparam i2_3_lut_adj_1019.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43318));   // verilog/coms.v(161[9:87])
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1021 (.I0(\data_in_frame[0] [0]), .I1(n43318), 
            .I2(n4_adj_3219), .I3(\data_in_frame[4] [4]), .O(n22801));   // verilog/coms.v(71[16:43])
    defparam i3_4_lut_adj_1021.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(\data_in_frame[6] [6]), .I1(n22801), 
            .I2(GND_net), .I3(GND_net), .O(n43795));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43394));   // verilog/coms.v(82[17:28])
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43584));   // verilog/coms.v(225[9:81])
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1025 (.I0(\data_in_frame[3] [7]), .I1(n43584), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[4] [1]), .O(n10_adj_3116));   // verilog/coms.v(225[9:81])
    defparam i3_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i10601_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n24016));
    defparam i10601_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1026 (.I0(\data_in_frame[4] [0]), .I1(n43394), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[1][4] ), .O(n23367));   // verilog/coms.v(82[17:28])
    defparam i3_4_lut_adj_1026.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[15] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43671));   // verilog/coms.v(69[16:41])
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1028 (.I0(n43388), .I1(n43367), .I2(n43870), 
            .I3(\data_in_frame[8] [5]), .O(n12_adj_3244));   // verilog/coms.v(68[16:27])
    defparam i5_4_lut_adj_1028.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1029 (.I0(n43684), .I1(n12_adj_3244), .I2(n43821), 
            .I3(n23209), .O(n23078));   // verilog/coms.v(68[16:27])
    defparam i6_4_lut_adj_1029.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1030 (.I0(n23078), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[17] [6]), .I3(GND_net), .O(n7_adj_3245));   // verilog/coms.v(67[16:27])
    defparam i2_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1031 (.I0(n40161), .I1(n43278), .I2(n40194), 
            .I3(\data_in_frame[17] [6]), .O(n12_adj_3246));
    defparam i5_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1032 (.I0(\data_in_frame[20] [0]), .I1(n12_adj_3246), 
            .I2(n43528), .I3(n44311), .O(n44324));
    defparam i6_4_lut_adj_1032.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1033 (.I0(n23169), .I1(\data_in_frame[20] [7]), 
            .I2(n23212), .I3(GND_net), .O(n8_adj_3247));
    defparam i1_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1034 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[16] [5]), 
            .I2(n40169), .I3(n22605), .O(n12_adj_3248));
    defparam i5_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1035 (.I0(n23078), .I1(n43789), .I2(n43528), 
            .I3(\data_in_frame[21] [7]), .O(n44580));
    defparam i2_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1036 (.I0(n43426), .I1(n43691), .I2(\data_in_frame[20] [3]), 
            .I3(GND_net), .O(n45075));
    defparam i2_3_lut_adj_1036.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1037 (.I0(n40149), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[21] [4]), .I3(n43730), .O(n44856));
    defparam i2_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 n50005_bdd_4_lut (.I0(n50005), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter_c[1]), 
            .O(n50008));
    defparam n50005_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(n20432), .I1(Kp_23__N_1179), .I2(GND_net), 
            .I3(GND_net), .O(n107));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_4_lut_adj_1039 (.I0(\data_in_frame[19] [3]), .I1(n43614), 
            .I2(n40149), .I3(\data_in_frame[21] [5]), .O(n44965));
    defparam i3_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1040 (.I0(\data_in_frame[20] [4]), .I1(\data_in_frame[18] [3]), 
            .I2(n40234), .I3(GND_net), .O(n14_adj_3249));
    defparam i5_3_lut_adj_1040.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1041 (.I0(n43718), .I1(\data_in_frame[13] [6]), 
            .I2(n40129), .I3(n43709), .O(n15_adj_3250));
    defparam i6_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1042 (.I0(n15_adj_3250), .I1(\data_in_frame[15] [7]), 
            .I2(n14_adj_3249), .I3(\data_in_frame[18][2] ), .O(n44172));
    defparam i8_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[20] [1]), .I1(n40194), .I2(n43278), 
            .I3(GND_net), .O(n8_adj_3251));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1043 (.I0(\data_in_frame[21] [6]), .I1(n44172), 
            .I2(n43614), .I3(n43789), .O(n18_adj_3252));
    defparam i1_4_lut_adj_1043.LUT_INIT = 16'h8448;
    SB_LUT4 i2_4_lut_adj_1044 (.I0(\data_in_frame[21] [0]), .I1(n23169), 
            .I2(Kp_23__N_785), .I3(n23212), .O(n44367));   // verilog/coms.v(73[16:43])
    defparam i2_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1045 (.I0(\data_in_frame[17] [7]), .I1(n18_adj_3252), 
            .I2(n8_adj_3251), .I3(n40161), .O(n26_adj_3253));
    defparam i9_4_lut_adj_1045.LUT_INIT = 16'h4884;
    SB_LUT4 i10602_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n24017));
    defparam i10602_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1046 (.I0(n7_adj_3245), .I1(n44311), .I2(\data_in_frame[20] [2]), 
            .I3(n43426), .O(n44888));   // verilog/coms.v(67[16:27])
    defparam i4_4_lut_adj_1046.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1047 (.I0(n43501), .I1(n44324), .I2(n43730), 
            .I3(\data_in_frame[21] [3]), .O(n24_adj_3254));
    defparam i7_4_lut_adj_1047.LUT_INIT = 16'h4884;
    SB_LUT4 i13_4_lut_adj_1048 (.I0(\data_in_frame[21] [1]), .I1(n26_adj_3253), 
            .I2(n44367), .I3(n23212), .O(n30_adj_3255));
    defparam i13_4_lut_adj_1048.LUT_INIT = 16'h4080;
    SB_LUT4 i3_4_lut_adj_1049 (.I0(\data_in_frame[21] [2]), .I1(n43501), 
            .I2(n23169), .I3(Kp_23__N_785), .O(n44977));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1050 (.I0(\data_in_frame[20] [5]), .I1(n45002), 
            .I2(\data_in_frame[18] [3]), .I3(n22605), .O(n8_adj_3256));
    defparam i3_4_lut_adj_1050.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1051 (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[16][1] ), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3257));
    defparam i2_2_lut_adj_1051.LUT_INIT = 16'h6666;
    SB_LUT4 i10603_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n24018));
    defparam i10603_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10540_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n23955));
    defparam i10540_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1052 (.I0(\data_in_frame[18] [5]), .I1(n44580), 
            .I2(n12_adj_3248), .I3(n8_adj_3247), .O(n20_adj_3258));
    defparam i3_4_lut_adj_1052.LUT_INIT = 16'h4884;
    SB_LUT4 i11_4_lut_adj_1053 (.I0(n44965), .I1(n107), .I2(n44856), .I3(n45075), 
            .O(n28_adj_3259));
    defparam i11_4_lut_adj_1053.LUT_INIT = 16'h4000;
    SB_LUT4 i15_4_lut (.I0(n44977), .I1(n30_adj_3255), .I2(n24_adj_3254), 
            .I3(n44888), .O(n32));
    defparam i15_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_4_lut_adj_1054 (.I0(\data_in_frame[20] [6]), .I1(n7_adj_3257), 
            .I2(n43453), .I3(n8_adj_3256), .O(n19_adj_3260));
    defparam i2_4_lut_adj_1054.LUT_INIT = 16'h2184;
    SB_LUT4 i16_4_lut_adj_1055 (.I0(n19_adj_3260), .I1(n32), .I2(n28_adj_3259), 
            .I3(n20_adj_3258), .O(n29738));
    defparam i16_4_lut_adj_1055.LUT_INIT = 16'h8000;
    SB_LUT4 i10541_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43235), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n23956));
    defparam i10541_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10526_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n23941));
    defparam i10526_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10604_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n24019));
    defparam i10604_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10527_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n23942));
    defparam i10527_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10528_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n23943));
    defparam i10528_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10529_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n23944));
    defparam i10529_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10530_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n23945));
    defparam i10530_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10531_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[2]), 
            .I3(\data_in_frame[18][2] ), .O(n23946));
    defparam i10531_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10605_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43247), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n24020));
    defparam i10605_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10532_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n23947));
    defparam i10532_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10533_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43235), .I2(rx_data[0]), 
            .I3(\data_in_frame[18][0] ), .O(n23948));
    defparam i10533_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10510_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n23925));
    defparam i10510_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10511_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n23926));
    defparam i10511_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_955_i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[16] [0]), .O(n3799));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i1_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10512_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n23927));
    defparam i10512_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32395_3_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(n29738), .I3(GND_net), .O(n47239));   // verilog/coms.v(125[12] 284[6])
    defparam i32395_3_lut_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 mux_955_i2_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [1]), .I3(\data_in_frame[16][1] ), .O(n3800));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i2_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10513_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n23928));
    defparam i10513_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10514_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n23929));
    defparam i10514_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3262));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32003_4_lut (.I0(byte_transmit_counter[0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter_c[2]), 
            .O(n47504));   // verilog/coms.v(103[34:55])
    defparam i32003_4_lut.LUT_INIT = 16'h880a;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3263));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29801_4_lut (.I0(n19_adj_3262), .I1(\data_out_frame[22] [0]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n45301));
    defparam i29801_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_955_i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[16] [2]), .O(n3801));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i3_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i29802_3_lut (.I0(n50026), .I1(n45301), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45302));
    defparam i29802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29773_4_lut (.I0(n5_adj_3263), .I1(n47504), .I2(byte_transmit_counter_c[2]), 
            .I3(byte_transmit_counter_c[1]), .O(n45273));
    defparam i29773_4_lut.LUT_INIT = 16'haccc;
    SB_LUT4 i29775_4_lut (.I0(n45273), .I1(n45302), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n45275));
    defparam i29775_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29774_3_lut (.I0(n50062), .I1(n50068), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45274));
    defparam i29774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_955_i4_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[16] [3]), .O(n3802));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i4_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_955_i5_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [4]), .I3(\data_in_frame[16] [4]), .O(n3803));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i5_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10515_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n23930));
    defparam i10515_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10516_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n23931));
    defparam i10516_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10517_3_lut_4_lut (.I0(n8), .I1(n43235), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n23932));
    defparam i10517_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_955_i6_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[16] [5]), .O(n3804));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i6_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_955_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[16] [6]), .O(n3805));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i7_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34500 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter_c[1]), .O(n49999));
    defparam byte_transmit_counter_0__bdd_4_lut_34500.LUT_INIT = 16'he4aa;
    SB_LUT4 n49999_bdd_4_lut (.I0(n49999), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter_c[1]), 
            .O(n50002));
    defparam n49999_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1056 (.I0(\FRAME_MATCHER.state_c [9]), .I1(\FRAME_MATCHER.state_c [11]), 
            .I2(\FRAME_MATCHER.state_c [8]), .I3(\FRAME_MATCHER.state_c [15]), 
            .O(n43132));
    defparam i3_4_lut_adj_1056.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1057 (.I0(\FRAME_MATCHER.state_c [4]), .I1(\FRAME_MATCHER.state_c [5]), 
            .I2(\FRAME_MATCHER.state_c [7]), .I3(\FRAME_MATCHER.state_c [6]), 
            .O(n43271));
    defparam i3_4_lut_adj_1057.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1058 (.I0(\FRAME_MATCHER.state_c [13]), .I1(\FRAME_MATCHER.state_c [12]), 
            .I2(\FRAME_MATCHER.state_c [10]), .I3(\FRAME_MATCHER.state_c [14]), 
            .O(n43273));   // verilog/coms.v(125[12] 284[6])
    defparam i3_4_lut_adj_1058.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1059 (.I0(\FRAME_MATCHER.state_c [25]), .I1(\FRAME_MATCHER.state_c [29]), 
            .I2(\FRAME_MATCHER.state_c [18]), .I3(\FRAME_MATCHER.state_c [16]), 
            .O(n18_adj_3264));   // verilog/coms.v(147[5:27])
    defparam i7_4_lut_adj_1059.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(\FRAME_MATCHER.state_c [19]), .I1(\FRAME_MATCHER.state_c [26]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3265));   // verilog/coms.v(147[5:27])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1060 (.I0(\FRAME_MATCHER.state_c [21]), .I1(n18_adj_3264), 
            .I2(\FRAME_MATCHER.state_c [28]), .I3(\FRAME_MATCHER.state_c [17]), 
            .O(n20_adj_3266));   // verilog/coms.v(147[5:27])
    defparam i9_4_lut_adj_1060.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i8_3_lut (.I0(\data_out_frame[8] [4]), 
            .I1(\data_out_frame[9] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n8_adj_3231));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i9_3_lut (.I0(\data_out_frame[10] [4]), 
            .I1(\data_out_frame[11] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n9));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1061 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n20_adj_3266), 
            .I2(n16_adj_3265), .I3(\FRAME_MATCHER.state_c [22]), .O(n43127));   // verilog/coms.v(147[5:27])
    defparam i10_4_lut_adj_1061.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\FRAME_MATCHER.state_c [24]), .I1(\FRAME_MATCHER.state_c [27]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3267));   // verilog/coms.v(125[12] 284[6])
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1063 (.I0(\FRAME_MATCHER.state_c [23]), .I1(\FRAME_MATCHER.state_c [31]), 
            .I2(\FRAME_MATCHER.state_c [20]), .I3(n6_adj_3267), .O(n43245));   // verilog/coms.v(125[12] 284[6])
    defparam i4_4_lut_adj_1063.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(n43271), .I1(n43132), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3268));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'heeee;
    SB_LUT4 i17692_3_lut (.I0(\data_in[0]_c [0]), .I1(\data_in[1] [0]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n23739));   // verilog/coms.v(87[7:20])
    defparam i17692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1065 (.I0(n43245), .I1(n43127), .I2(n43273), 
            .I3(n4_adj_3268), .O(n28723));
    defparam i2_4_lut_adj_1065.LUT_INIT = 16'hfffe;
    SB_LUT4 i28509_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n28723), .I2(GND_net), 
            .I3(GND_net), .O(n44005));
    defparam i28509_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10787_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[9]), .I3(\data_out_frame[7] [1]), .O(n24202));
    defparam i10787_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i29752_4_lut (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[2] [5]), .O(n45252));
    defparam i29752_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1066 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [6]), .O(n38));
    defparam i14_4_lut_adj_1066.LUT_INIT = 16'h8000;
    SB_LUT4 i15_4_lut_adj_1067 (.I0(\data_in_frame[1][4] ), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[2] [4]), .O(n39));
    defparam i15_4_lut_adj_1067.LUT_INIT = 16'h0002;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i12_3_lut (.I0(\data_out_frame[14] [4]), 
            .I1(\data_out_frame[15] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n12_adj_3229));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i11_3_lut (.I0(\data_out_frame[12] [4]), 
            .I1(\data_out_frame[13] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n11));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_277_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3228));
    defparam select_277_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1068 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [2]), .O(n37_adj_3269));
    defparam i13_4_lut_adj_1068.LUT_INIT = 16'h2000;
    SB_LUT4 i29748_4_lut (.I0(\data_in_frame[2] [2]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [3]), .O(n45248));
    defparam i29748_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1069 (.I0(n37_adj_3269), .I1(n39), .I2(n38), 
            .I3(n45252), .O(n46));
    defparam i22_4_lut_adj_1069.LUT_INIT = 16'h0080;
    SB_LUT4 mux_955_i8_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[16] [7]), .O(n3806));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i8_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i29750_4_lut (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[0] [1]), .O(n45250));
    defparam i29750_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_3_lut (.I0(n45250), .I1(n46), .I2(n45248), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_1924 [3]));
    defparam i23_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i10786_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[10]), .I3(\data_out_frame[7] [2]), .O(n24201));
    defparam i10786_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i22971_3_lut (.I0(n23530), .I1(r_SM_Main[1]), .I2(tx_active), 
            .I3(GND_net), .O(n25425));   // verilog/uart_tx.v(31[16:25])
    defparam i22971_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(n5024), .I1(\FRAME_MATCHER.state_31__N_1924 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n22429));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h8888;
    SB_LUT4 i10788_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[8]), .I3(\data_out_frame[7] [0]), .O(n24203));
    defparam i10788_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i9_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [0]), .I3(\data_in_frame[15] [0]), .O(n3807));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i9_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10678_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[6]), .I3(\data_out_frame[20] [6]), .O(n24093));
    defparam i10678_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i10_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[15] [1]), .O(n3808));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i10_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10769_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[19]), .I3(\data_out_frame[9] [3]), .O(n24184));
    defparam i10769_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10797_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(control_mode[7]), .I3(\data_out_frame[5] [7]), .O(n24212));
    defparam i10797_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10799_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(control_mode[5]), .I3(\data_out_frame[5] [5]), .O(n24214));
    defparam i10799_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10743_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[21]), .I3(\data_out_frame[12] [5]), .O(n24158));
    defparam i10743_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10740_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[8]), .I3(\data_out_frame[13] [0]), .O(n24155));
    defparam i10740_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10742_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[22]), .I3(\data_out_frame[12] [6]), .O(n24157));
    defparam i10742_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i11_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[15] [2]), .O(n3809));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i11_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_955_i12_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [3]), .I3(\data_in_frame[15] [3]), .O(n3810));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i12_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_955_i13_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [4]), .I3(\data_in_frame[15] [4]), .O(n3811));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i13_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10741_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[23]), .I3(\data_out_frame[12] [7]), .O(n24156));
    defparam i10741_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10744_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[20]), .I3(\data_out_frame[12] [4]), .O(n24159));
    defparam i10744_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10745_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[19]), .I3(\data_out_frame[12] [3]), .O(n24160));
    defparam i10745_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10746_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[18]), .I3(\data_out_frame[12] [2]), .O(n24161));
    defparam i10746_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10747_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[17]), .I3(\data_out_frame[12] [1]), .O(n24162));
    defparam i10747_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3270));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_955_i14_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[15] [5]), .O(n3812));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i14_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i29771_4_lut (.I0(n19_adj_3270), .I1(\data_out_frame[22] [7]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n45271));
    defparam i29771_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32175_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n47677));   // verilog/coms.v(103[34:55])
    defparam i32175_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3271));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29772_3_lut (.I0(n50002), .I1(n45271), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45272));
    defparam i29772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29797_4_lut (.I0(n5_adj_3271), .I1(n47677), .I2(n47022), 
            .I3(byte_transmit_counter[0]), .O(n45297));
    defparam i29797_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29799_4_lut (.I0(n45297), .I1(n45272), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n45299));
    defparam i29799_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i17130_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[15]), .I3(\data_out_frame[19] [7]), .O(n24100));
    defparam i17130_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3272));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29768_4_lut (.I0(n19_adj_3272), .I1(\data_out_frame[22] [6]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n45268));
    defparam i29768_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32168_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n47670));   // verilog/coms.v(103[34:55])
    defparam i32168_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3273));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29769_3_lut (.I0(n49996), .I1(n45268), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45269));
    defparam i29769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29794_4_lut (.I0(n5_adj_3273), .I1(n47670), .I2(n47022), 
            .I3(byte_transmit_counter[0]), .O(n45294));
    defparam i29794_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29796_4_lut (.I0(n45294), .I1(n45269), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n45296));
    defparam i29796_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_955_i15_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[15] [6]), .O(n3813));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i15_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10721_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[19]), .I3(\data_out_frame[15] [3]), .O(n24136));
    defparam i10721_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10789_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[23]), .I3(\data_out_frame[6] [7]), .O(n24204));
    defparam i10789_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10790_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[22]), .I3(\data_out_frame[6] [6]), .O(n24205));
    defparam i10790_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3274));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10749_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[7]), .I3(\data_out_frame[11] [7]), .O(n24164));
    defparam i10749_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter_c[1]), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n47665));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3275));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29765_4_lut (.I0(n19_adj_3274), .I1(\data_out_frame[22] [5]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n45265));
    defparam i29765_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29766_3_lut (.I0(n49990), .I1(n45265), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45266));
    defparam i29766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29791_4_lut (.I0(n5_adj_3275), .I1(byte_transmit_counter[0]), 
            .I2(n47022), .I3(n47665), .O(n45291));
    defparam i29791_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29793_4_lut (.I0(n45291), .I1(n45266), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n45293));
    defparam i29793_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29792_3_lut (.I0(n49966), .I1(n50098), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45292));
    defparam i29792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17693_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2]_c [0]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n24246));   // verilog/coms.v(87[7:20])
    defparam i17693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10750_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[6]), .I3(\data_out_frame[11] [6]), .O(n24165));
    defparam i10750_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13870_3_lut (.I0(\data_in[0]_c [7]), .I1(\data_in[1] [7]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n24247));   // verilog/coms.v(87[7:20])
    defparam i13870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10791_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[21]), .I3(\data_out_frame[6] [5]), .O(n24206));
    defparam i10791_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3276));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29762_4_lut (.I0(n19_adj_3276), .I1(\data_out_frame[22] [4]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n45262));
    defparam i29762_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29763_3_lut (.I0(n49984), .I1(n45262), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45263));
    defparam i29763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33377_3_lut (.I0(n50086), .I1(n50014), .I2(byte_transmit_counter_c[3]), 
            .I3(GND_net), .O(n48879));   // verilog/coms.v(103[34:55])
    defparam i33377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33378_4_lut (.I0(n48879), .I1(n45263), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(tx_data[4]));   // verilog/coms.v(103[34:55])
    defparam i33378_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10792_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[20]), .I3(\data_out_frame[6] [4]), .O(n24207));
    defparam i10792_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10793_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[19]), .I3(\data_out_frame[6] [3]), .O(n24208));
    defparam i10793_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10794_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[18]), .I3(\data_out_frame[6] [2]), .O(n24209));
    defparam i10794_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i32151_2_lut (.I0(\data_out_frame[0][3] ), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n47202));   // verilog/coms.v(103[34:55])
    defparam i32151_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n47202), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3277));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3278));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29782_3_lut (.I0(n5_adj_3278), .I1(n6_adj_3277), .I2(n47022), 
            .I3(GND_net), .O(n45282));
    defparam i29782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29784_4_lut (.I0(n45282), .I1(n50092), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n45284));
    defparam i29784_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29783_3_lut (.I0(n49978), .I1(n49972), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45283));
    defparam i29783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10796_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[16]), .I3(\data_out_frame[6] [0]), .O(n24211));
    defparam i10796_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10751_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[5]), .I3(\data_out_frame[11] [5]), .O(n24166));
    defparam i10751_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i32394_2_lut (.I0(\data_out_frame[0][2] ), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n47199));   // verilog/coms.v(103[34:55])
    defparam i32394_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3279));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5][2] ), 
            .I1(n47199), .I2(byte_transmit_counter_c[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_3280));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'ha00c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3281));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29807_4_lut (.I0(n19_adj_3279), .I1(\data_out_frame[22] [2]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n45307));
    defparam i29807_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29808_3_lut (.I0(n50038), .I1(n45307), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45308));
    defparam i29808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29779_3_lut (.I0(n5_adj_3281), .I1(n6_adj_3280), .I2(n47022), 
            .I3(GND_net), .O(n45279));
    defparam i29779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29781_4_lut (.I0(n45279), .I1(n45308), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n45281));
    defparam i29781_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29780_3_lut (.I0(n50044), .I1(n50008), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45280));
    defparam i29780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10752_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[4]), .I3(\data_out_frame[11] [4]), .O(n24167));
    defparam i10752_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10753_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[3]), .I3(\data_out_frame[11] [3]), .O(n24168));
    defparam i10753_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10754_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[2]), .I3(\data_out_frame[11] [2]), .O(n24169));
    defparam i10754_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10798_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(control_mode[6]), .I3(\data_out_frame[5] [6]), .O(n24213));
    defparam i10798_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_3282));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32144_2_lut (.I0(byte_transmit_counter_c[2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n47645));   // verilog/coms.v(103[34:55])
    defparam i32144_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_3283));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29804_4_lut (.I0(n19_adj_3282), .I1(\data_out_frame[22] [1]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter[0]), 
            .O(n45304));
    defparam i29804_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29805_3_lut (.I0(n50032), .I1(n45304), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45305));
    defparam i29805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29776_4_lut (.I0(n5_adj_3283), .I1(n47645), .I2(n47022), 
            .I3(byte_transmit_counter[0]), .O(n45276));
    defparam i29776_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i29778_4_lut (.I0(n45276), .I1(n45305), .I2(byte_transmit_counter_c[4]), 
            .I3(byte_transmit_counter_c[3]), .O(n45278));
    defparam i29778_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i29777_3_lut (.I0(n50056), .I1(n50050), .I2(byte_transmit_counter_c[2]), 
            .I3(GND_net), .O(n45277));
    defparam i29777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10801_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(control_mode[3]), .I3(\data_out_frame[5] [3]), .O(n24216));
    defparam i10801_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10760_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[12]), .I3(\data_out_frame[10] [4]), .O(n24175));
    defparam i10760_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10756_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[0]), .I3(\data_out_frame[11] [0]), .O(n24171));
    defparam i10756_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i16_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[2] [7]), .I3(\data_in_frame[15] [7]), .O(n3814));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i16_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17701_3_lut (.I0(\data_in[2][1] ), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n27276));   // verilog/coms.v(87[7:20])
    defparam i17701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17700_3_lut (.I0(\data_in[2]_c [0]), .I1(\data_in[3] [0]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n24238));   // verilog/coms.v(87[7:20])
    defparam i17700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10757_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[15]), .I3(\data_out_frame[10] [7]), .O(n24172));
    defparam i10757_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i28591_3_lut (.I0(n28723), .I1(\FRAME_MATCHER.state [3]), .I2(n44238), 
            .I3(GND_net), .O(n44089));
    defparam i28591_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i31875_4_lut (.I0(n47), .I1(\FRAME_MATCHER.state [2]), .I2(tx_transmit_N_2639), 
            .I3(\FRAME_MATCHER.state [0]), .O(n47095));   // verilog/coms.v(109[11:16])
    defparam i31875_4_lut.LUT_INIT = 16'hc044;
    SB_LUT4 i16394_4_lut (.I0(n28723), .I1(n29738), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n23_adj_3284));   // verilog/coms.v(109[11:16])
    defparam i16394_4_lut.LUT_INIT = 16'hc5c0;
    SB_LUT4 i16398_4_lut (.I0(n23_adj_3284), .I1(n47095), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [0]), .O(n2416[0]));   // verilog/coms.v(109[11:16])
    defparam i16398_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i13871_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2]_c [7]), 
            .I2(rx_data_ready), .I3(GND_net), .O(n24239));   // verilog/coms.v(87[7:20])
    defparam i13871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_955_i17_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[14][0] ), .O(n3815));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i17_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10758_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[14]), .I3(\data_out_frame[10] [6]), .O(n24173));
    defparam i10758_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_4_lut_adj_1071 (.I0(n5024), .I1(n47239), .I2(\FRAME_MATCHER.state_31__N_1924 [3]), 
            .I3(n5022), .O(n23563));
    defparam i1_4_lut_adj_1071.LUT_INIT = 16'ha088;
    SB_LUT4 i10759_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[13]), .I3(\data_out_frame[10] [5]), .O(n24174));
    defparam i10759_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i19_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[14]_c [2]), .O(n3817));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i19_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_955_i20_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[14]_c [3]), .O(n3818));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i20_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_4_lut_adj_1072 (.I0(\FRAME_MATCHER.state [3]), .I1(n44005), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n5022));
    defparam i2_4_lut_adj_1072.LUT_INIT = 16'h0102;
    SB_LUT4 i10761_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[11]), .I3(\data_out_frame[10] [3]), .O(n24176));
    defparam i10761_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10766_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[22]), .I3(\data_out_frame[9] [6]), .O(n24181));
    defparam i10766_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i24_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[14]_c [7]), .O(n3822));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i24_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 mux_955_i18_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[14]_c [1]), .O(n3816));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i18_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17696_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24224));   // verilog/coms.v(87[7:20])
    defparam i17696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10762_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[10]), .I3(\data_out_frame[10] [2]), .O(n24177));
    defparam i10762_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i22_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[14]_c [5]), .O(n3820));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i22_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10763_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[9]), .I3(\data_out_frame[10] [1]), .O(n24178));
    defparam i10763_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 mux_955_i23_3_lut_4_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n47), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[14]_c [6]), .O(n3821));   // verilog/coms.v(125[12] 284[6])
    defparam mux_955_i23_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10764_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[8]), .I3(\data_out_frame[10] [0]), .O(n24179));
    defparam i10764_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10767_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[21]), .I3(\data_out_frame[9] [5]), .O(n24182));
    defparam i10767_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10771_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[17]), .I3(\data_out_frame[9] [1]), .O(n24186));
    defparam i10771_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i17695_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24229));   // verilog/coms.v(87[7:20])
    defparam i17695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10772_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[16]), .I3(\data_out_frame[9] [0]), .O(n24187));
    defparam i10772_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10590_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n24005));
    defparam i10590_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10776_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[4]), .I3(\data_out_frame[8] [4]), .O(n24191));
    defparam i10776_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i17694_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24230));   // verilog/coms.v(87[7:20])
    defparam i17694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10773_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[7]), .I3(\data_out_frame[8] [7]), .O(n24188));
    defparam i10773_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13869_3_lut (.I0(\data_in[2]_c [7]), .I1(\data_in[3][7] ), 
            .I2(rx_data_ready), .I3(GND_net), .O(n24231));   // verilog/coms.v(87[7:20])
    defparam i13869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10774_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[6]), .I3(\data_out_frame[8] [6]), .O(n24189));
    defparam i10774_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i17697_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n24232));   // verilog/coms.v(87[7:20])
    defparam i17697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10775_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[5]), .I3(\data_out_frame[8] [5]), .O(n24190));
    defparam i10775_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10777_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[3]), .I3(\data_out_frame[8] [3]), .O(n24192));
    defparam i10777_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10778_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[2]), .I3(\data_out_frame[8] [2]), .O(n24193));
    defparam i10778_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10779_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[1]), .I3(\data_out_frame[8] [1]), .O(n24194));
    defparam i10779_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10781_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[15]), .I3(\data_out_frame[7] [7]), .O(n24196));
    defparam i10781_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10782_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[14]), .I3(\data_out_frame[7] [6]), .O(n24197));
    defparam i10782_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i17702_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3][3] ), .I2(rx_data_ready), 
            .I3(GND_net), .O(n27275));   // verilog/coms.v(87[7:20])
    defparam i17702_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10677_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[7]), .I3(\data_out_frame[20] [7]), .O(n24092));
    defparam i10677_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10679_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[5]), .I3(\data_out_frame[20] [5]), .O(n24094));
    defparam i10679_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10680_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[4]), .I3(\data_out_frame[20] [4]), .O(n24095));
    defparam i10680_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10681_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[3]), .I3(\data_out_frame[20] [3]), .O(n24096));
    defparam i10681_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10682_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[2]), .I3(\data_out_frame[20] [2]), .O(n24097));
    defparam i10682_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10683_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[1]), .I3(\data_out_frame[20] [1]), .O(n24098));
    defparam i10683_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10684_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[0]), .I3(\data_out_frame[20] [0]), .O(n24099));
    defparam i10684_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i69_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n31), .I2(n63), 
            .I3(GND_net), .O(n122));   // verilog/coms.v(109[11:16])
    defparam i69_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_312_Select_2_i7_4_lut (.I0(n103), .I1(n22442), .I2(n3758), 
            .I3(n122), .O(n7));
    defparam select_312_Select_2_i7_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i10686_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[14]), .I3(\data_out_frame[19] [6]), .O(n24101));
    defparam i10686_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_312_Select_2_i5_4_lut (.I0(n2854), .I1(n22454), .I2(n103), 
            .I3(n122), .O(n5));
    defparam select_312_Select_2_i5_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i10691_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[9]), .I3(\data_out_frame[19] [1]), .O(n24106));
    defparam i10691_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10687_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[13]), .I3(\data_out_frame[19] [5]), .O(n24102));
    defparam i10687_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10688_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[12]), .I3(\data_out_frame[19] [4]), .O(n24103));
    defparam i10688_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10689_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[11]), .I3(\data_out_frame[19] [3]), .O(n24104));
    defparam i10689_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10690_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[10]), .I3(\data_out_frame[19] [2]), .O(n24105));
    defparam i10690_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10692_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[8]), .I3(\data_out_frame[19] [0]), .O(n24107));
    defparam i10692_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10693_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[23]), .I3(\data_out_frame[18] [7]), .O(n24108));
    defparam i10693_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10695_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[21]), .I3(\data_out_frame[18] [5]), .O(n24110));
    defparam i10695_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10696_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[20]), .I3(\data_out_frame[18] [4]), .O(n24111));
    defparam i10696_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10591_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[6]), 
            .I3(\data_in_frame[10][6] ), .O(n24006));
    defparam i10591_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10697_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[19]), .I3(\data_out_frame[18] [3]), .O(n24112));
    defparam i10697_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10698_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[18]), .I3(\data_out_frame[18] [2]), .O(n24113));
    defparam i10698_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10699_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[17]), .I3(\data_out_frame[18] [1]), .O(n24114));
    defparam i10699_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10703_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[5]), .I3(\data_out_frame[17] [5]), .O(n24118));
    defparam i10703_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10700_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[16]), .I3(\data_out_frame[18] [0]), .O(n24115));
    defparam i10700_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10702_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[6]), .I3(\data_out_frame[17] [6]), .O(n24117));
    defparam i10702_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10704_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[4]), .I3(\data_out_frame[17] [4]), .O(n24119));
    defparam i10704_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10706_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[2]), .I3(\data_out_frame[17] [2]), .O(n24121));
    defparam i10706_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10707_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[1]), .I3(\data_out_frame[17] [1]), .O(n24122));
    defparam i10707_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10708_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[0]), .I3(\data_out_frame[17] [0]), .O(n24123));
    defparam i10708_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10709_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[15]), .I3(\data_out_frame[16] [7]), .O(n24124));
    defparam i10709_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10710_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[14]), .I3(\data_out_frame[16] [6]), .O(n24125));
    defparam i10710_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10713_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[11]), .I3(\data_out_frame[16] [3]), .O(n24128));
    defparam i10713_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10714_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[10]), .I3(\data_out_frame[16] [2]), .O(n24129));
    defparam i10714_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10715_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[9]), .I3(\data_out_frame[16] [1]), .O(n24130));
    defparam i10715_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10716_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[8]), .I3(\data_out_frame[16] [0]), .O(n24131));
    defparam i10716_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10717_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[23]), .I3(\data_out_frame[15] [7]), .O(n24132));
    defparam i10717_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10718_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[22]), .I3(\data_out_frame[15] [6]), .O(n24133));
    defparam i10718_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10719_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[21]), .I3(\data_out_frame[15] [5]), .O(n24134));
    defparam i10719_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10720_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[20]), .I3(\data_out_frame[15] [4]), .O(n24135));
    defparam i10720_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10722_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[18]), .I3(\data_out_frame[15] [2]), .O(n24137));
    defparam i10722_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10723_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[17]), .I3(\data_out_frame[15] [1]), .O(n24138));
    defparam i10723_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10724_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[16]), .I3(\data_out_frame[15] [0]), .O(n24139));
    defparam i10724_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10725_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[7]), .I3(\data_out_frame[14] [7]), .O(n24140));
    defparam i10725_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10592_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n24007));
    defparam i10592_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10726_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[6]), .I3(\data_out_frame[14] [6]), .O(n24141));
    defparam i10726_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3196));
    defparam select_277_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10727_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[5]), .I3(\data_out_frame[14] [5]), .O(n24142));
    defparam i10727_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3194));
    defparam select_277_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3192));
    defparam select_277_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10728_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[4]), .I3(\data_out_frame[14] [4]), .O(n24143));
    defparam i10728_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3191));
    defparam select_277_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3190));
    defparam select_277_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3189));
    defparam select_277_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3187));
    defparam select_277_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10729_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[3]), .I3(\data_out_frame[14] [3]), .O(n24144));
    defparam i10729_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3185));
    defparam select_277_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3183));
    defparam select_277_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3181));
    defparam select_277_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3179));
    defparam select_277_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3178));
    defparam select_277_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10730_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[2]), .I3(\data_out_frame[14] [2]), .O(n24145));
    defparam i10730_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3177));
    defparam select_277_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3176));
    defparam select_277_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3175));
    defparam select_277_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3174));
    defparam select_277_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3173));
    defparam select_277_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3172));
    defparam select_277_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3170));
    defparam select_277_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3168));
    defparam select_277_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3166));
    defparam select_277_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3164));
    defparam select_277_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10731_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[1]), .I3(\data_out_frame[14] [1]), .O(n24146));
    defparam i10731_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10732_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[0]), .I3(\data_out_frame[14] [0]), .O(n24147));
    defparam i10732_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3162));
    defparam select_277_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3160));
    defparam select_277_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10733_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[15]), .I3(\data_out_frame[13] [7]), .O(n24148));
    defparam i10733_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3158));
    defparam select_277_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10734_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[14]), .I3(\data_out_frame[13] [6]), .O(n24149));
    defparam i10734_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 select_277_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3156));
    defparam select_277_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3154));
    defparam select_277_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3152));
    defparam select_277_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3150));
    defparam select_277_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3148));
    defparam select_277_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_277_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2123), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_277_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i10735_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[13]), .I3(\data_out_frame[13] [5]), .O(n24150));
    defparam i10735_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10736_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[12]), .I3(\data_out_frame[13] [4]), .O(n24151));
    defparam i10736_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10737_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[11]), .I3(\data_out_frame[13] [3]), .O(n24152));
    defparam i10737_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10738_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[10]), .I3(\data_out_frame[13] [2]), .O(n24153));
    defparam i10738_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_3_lut_adj_1073 (.I0(n22133), .I1(\data_out_frame[20] [7]), 
            .I2(n43450), .I3(GND_net), .O(n8_adj_3287));   // verilog/coms.v(68[16:27])
    defparam i3_3_lut_adj_1073.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1074 (.I0(n22984), .I1(n8_adj_3287), .I2(\data_out_frame[20] [6]), 
            .I3(n23259), .O(n44821));   // verilog/coms.v(68[16:27])
    defparam i4_4_lut_adj_1074.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1075 (.I0(n39498), .I1(n43284), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_3288));
    defparam i2_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1076 (.I0(n7_adj_3288), .I1(\data_out_frame[20] [7]), 
            .I2(n44835), .I3(n43608), .O(n44955));
    defparam i4_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i10783_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[13]), .I3(\data_out_frame[7] [5]), .O(n24198));
    defparam i10783_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\data_out_frame[18] [6]), .I1(n43652), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3289));
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i10780_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[0]), .I3(\data_out_frame[8] [0]), .O(n24195));
    defparam i10780_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(\data_out_frame[19] [1]), .I1(n1713), 
            .I2(n43314), .I3(n6_adj_3289), .O(n45043));
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(n39866), .I1(n23282), .I2(GND_net), 
            .I3(GND_net), .O(n43608));
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1080 (.I0(n23436), .I1(n43620), .I2(n43608), 
            .I3(\data_out_frame[19] [1]), .O(n44983));
    defparam i3_4_lut_adj_1080.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[17] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43620));
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34495 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter_c[1]), .O(n49993));
    defparam byte_transmit_counter_0__bdd_4_lut_34495.LUT_INIT = 16'he4aa;
    SB_LUT4 n49993_bdd_4_lut (.I0(n49993), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter_c[1]), 
            .O(n49996));
    defparam n49993_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10770_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[18]), .I3(\data_out_frame[9] [2]), .O(n24185));
    defparam i10770_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10768_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[20]), .I3(\data_out_frame[9] [4]), .O(n24183));
    defparam i10768_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_1082 (.I0(\data_out_frame[16] [7]), .I1(n43786), 
            .I2(n43611), .I3(n43605), .O(n43284));
    defparam i3_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34490 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n49987));
    defparam byte_transmit_counter_0__bdd_4_lut_34490.LUT_INIT = 16'he4aa;
    SB_LUT4 n49987_bdd_4_lut (.I0(n49987), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n49990));
    defparam n49987_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1083 (.I0(n22809), .I1(n43284), .I2(n23436), 
            .I3(\data_out_frame[19] [3]), .O(n44887));
    defparam i3_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34485 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter_c[1]), .O(n49981));
    defparam byte_transmit_counter_0__bdd_4_lut_34485.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1084 (.I0(n43581), .I1(n43777), .I2(n44887), 
            .I3(GND_net), .O(n44383));
    defparam i2_3_lut_adj_1084.LUT_INIT = 16'h9696;
    SB_LUT4 i10765_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[23]), .I3(\data_out_frame[9] [7]), .O(n24180));
    defparam i10765_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10804_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(control_mode[0]), .I3(\data_out_frame[5] [0]), .O(n24219));
    defparam i10804_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1085 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43777));
    defparam i1_2_lut_adj_1085.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1086 (.I0(n43590), .I1(n1692), .I2(\data_out_frame[15] [0]), 
            .I3(n43694), .O(n10_adj_3225));
    defparam i4_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1087 (.I0(n43688), .I1(n23436), .I2(n39462), 
            .I3(n43777), .O(n10_adj_3290));
    defparam i4_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1088 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3291));
    defparam i2_2_lut_adj_1088.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1089 (.I0(\data_out_frame[8] [5]), .I1(n40119), 
            .I2(n43697), .I3(\data_out_frame[13] [0]), .O(n14_adj_3292));
    defparam i6_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i10803_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(control_mode[1]), .I3(\data_out_frame[5] [1]), .O(n24218));
    defparam i10803_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i7_4_lut_adj_1090 (.I0(\data_out_frame[15] [1]), .I1(n14_adj_3292), 
            .I2(n10_adj_3291), .I3(n43837), .O(n43605));
    defparam i7_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i10800_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(control_mode[4]), .I3(\data_out_frame[5] [4]), .O(n24215));
    defparam i10800_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_adj_1091 (.I0(n39990), .I1(n43605), .I2(\data_out_frame[14] [7]), 
            .I3(GND_net), .O(n39462));
    defparam i2_3_lut_adj_1091.LUT_INIT = 16'h9696;
    SB_LUT4 i10755_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder1_position[1]), .I3(\data_out_frame[11] [1]), .O(n24170));
    defparam i10755_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_out_frame[17] [3]), .I1(n23405), 
            .I2(GND_net), .I3(GND_net), .O(n43581));
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 i10795_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[17]), .I3(\data_out_frame[6] [1]), .O(n24210));
    defparam i10795_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10785_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[11]), .I3(\data_out_frame[7] [3]), .O(n24200));
    defparam i10785_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10712_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[12]), .I3(\data_out_frame[16] [4]), .O(n24127));
    defparam i10712_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_1093 (.I0(n44835), .I1(n44973), .I2(n43581), 
            .I3(n6_adj_3293), .O(n45019));
    defparam i4_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i10748_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[16]), .I3(\data_out_frame[12] [0]), .O(n24163));
    defparam i10748_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1094 (.I0(\data_out_frame[17] [5]), .I1(n1784), 
            .I2(GND_net), .I3(GND_net), .O(n43599));
    defparam i1_2_lut_adj_1094.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_out_frame[16] [3]), .I1(\data_out_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n23259));
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1096 (.I0(\data_out_frame[16] [6]), .I1(n43326), 
            .I2(\data_out_frame[14] [6]), .I3(n39781), .O(n12_adj_3294));
    defparam i5_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1097 (.I0(n23259), .I1(n12_adj_3294), .I2(n43813), 
            .I3(\data_out_frame[18] [7]), .O(n39866));
    defparam i6_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1098 (.I0(\data_out_frame[18] [7]), .I1(n39866), 
            .I2(\data_out_frame[16] [4]), .I3(\data_out_frame[19] [0]), 
            .O(n43652));
    defparam i3_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43385));   // verilog/coms.v(94[12:26])
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1100 (.I0(n39404), .I1(n43807), .I2(\data_out_frame[16] [5]), 
            .I3(n43465), .O(n20_adj_3295));
    defparam i8_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1101 (.I0(n43450), .I1(n23381), .I2(\data_out_frame[18] [4]), 
            .I3(n43647), .O(n19_adj_3296));
    defparam i7_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1102 (.I0(n22146), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[18] [3]), .I3(\data_out_frame[18] [7]), 
            .O(n21));
    defparam i9_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut (.I0(n21), .I1(n19_adj_3296), .I2(n20_adj_3295), 
            .I3(GND_net), .O(n44765));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1103 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[19] [7]), 
            .I2(n44765), .I3(\data_out_frame[19] [4]), .O(n12_adj_3297));   // verilog/coms.v(94[12:26])
    defparam i5_4_lut_adj_1103.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1104 (.I0(\data_out_frame[19] [2]), .I1(n12_adj_3297), 
            .I2(n43385), .I3(\data_out_frame[19] [3]), .O(n39498));   // verilog/coms.v(94[12:26])
    defparam i6_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1105 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [4]), 
            .I2(n43409), .I3(\data_out_frame[20] [1]), .O(n14_adj_3298));
    defparam i6_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1106 (.I0(n43295), .I1(n14_adj_3298), .I2(n10_adj_3217), 
            .I3(n22166), .O(n43638));
    defparam i7_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1107 (.I0(n43810), .I1(\data_out_frame[14] [4]), 
            .I2(n43599), .I3(\data_out_frame[14] [6]), .O(n24_adj_3299));
    defparam i10_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut (.I0(n43652), .I1(n22190), .I2(GND_net), .I3(GND_net), 
            .O(n17_adj_3300));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i10711_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[13]), .I3(\data_out_frame[16] [5]), .O(n24126));
    defparam i10711_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i8_4_lut_adj_1108 (.I0(n43864), .I1(n43329), .I2(n22771), 
            .I3(n39498), .O(n22_adj_3301));
    defparam i8_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i10593_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n24008));
    defparam i10593_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_4_lut_adj_1109 (.I0(n17_adj_3300), .I1(n24_adj_3299), .I2(n40167), 
            .I3(n43891), .O(n26_adj_3302));
    defparam i12_4_lut_adj_1109.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut_adj_1110 (.I0(\data_out_frame[17] [0]), .I1(n26_adj_3302), 
            .I2(n22_adj_3301), .I3(\data_out_frame[16] [5]), .O(n22126));
    defparam i13_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(n22126), .I1(n43638), .I2(GND_net), 
            .I3(GND_net), .O(n43282));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h9999;
    SB_LUT4 i2_2_lut_adj_1112 (.I0(n43767), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3303));   // verilog/coms.v(72[16:27])
    defparam i2_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i10705_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[3]), .I3(\data_out_frame[17] [3]), .O(n24120));
    defparam i10705_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10594_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n24009));
    defparam i10594_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1113 (.I0(n43861), .I1(\data_out_frame[10] [7]), 
            .I2(n43554), .I3(\data_out_frame[13] [1]), .O(n14_adj_3304));   // verilog/coms.v(72[16:27])
    defparam i6_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1114 (.I0(\data_out_frame[15] [2]), .I1(n14_adj_3304), 
            .I2(n10_adj_3303), .I3(\data_out_frame[8] [6]), .O(n23405));   // verilog/coms.v(72[16:27])
    defparam i7_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(n23405), .I1(\data_out_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43617));
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1116 (.I0(n1592), .I1(n43403), .I2(\data_out_frame[13] [1]), 
            .I3(n22596), .O(n1784));   // verilog/coms.v(70[16:42])
    defparam i3_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1117 (.I0(n39504), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[20] [0]), .I3(n1784), .O(n12_adj_3305));
    defparam i5_4_lut_adj_1117.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1118 (.I0(\data_out_frame[17] [6]), .I1(n12_adj_3305), 
            .I2(n43617), .I3(\data_out_frame[19] [6]), .O(n44973));
    defparam i6_4_lut_adj_1118.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1119 (.I0(n44973), .I1(\data_out_frame[20] [1]), 
            .I2(n39844), .I3(GND_net), .O(n44772));
    defparam i2_3_lut_adj_1119.LUT_INIT = 16'h9696;
    SB_LUT4 i10784_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(encoder0_position[12]), .I3(\data_out_frame[7] [4]), .O(n24199));
    defparam i10784_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_out_frame[12] [7]), .I1(n43861), 
            .I2(GND_net), .I3(GND_net), .O(n43697));
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1121 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[10] [7]), 
            .I2(n43292), .I3(n6_adj_3306), .O(n1592));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1122 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[17] [5]), .I3(GND_net), .O(n43647));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1122.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1123 (.I0(\data_out_frame[15] [3]), .I1(n43419), 
            .I2(n1503), .I3(n1592), .O(n43688));   // verilog/coms.v(70[16:42])
    defparam i3_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1124 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43403));   // verilog/coms.v(70[16:42])
    defparam i1_2_lut_adj_1124.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43419));   // verilog/coms.v(70[16:42])
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43864));
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43554));
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43355));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1129 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22746));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1129.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1130 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n23337));   // verilog/coms.v(68[16:62])
    defparam i1_2_lut_adj_1130.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1131 (.I0(\data_out_frame[10] [4]), .I1(n43447), 
            .I2(n23337), .I3(\data_out_frame[8] [3]), .O(n22771));   // verilog/coms.v(70[16:34])
    defparam i3_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i10701_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(pwm[7]), .I3(\data_out_frame[17] [7]), .O(n24116));
    defparam i10701_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10595_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n24010));
    defparam i10595_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10739_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(setpoint[9]), .I3(\data_out_frame[13] [1]), .O(n24154));
    defparam i10739_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i18_4_lut_adj_1132 (.I0(\data_out_frame[11] [7]), .I1(n43767), 
            .I2(n43412), .I3(n23331), .O(n52_adj_3307));   // verilog/coms.v(71[16:27])
    defparam i18_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i10694_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n22429), 
            .I2(displacement[22]), .I3(\data_out_frame[18] [6]), .O(n24109));
    defparam i10694_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i22_4_lut_adj_1133 (.I0(\data_out_frame[12] [7]), .I1(n43375), 
            .I2(n43694), .I3(n43703), .O(n56_adj_3308));   // verilog/coms.v(71[16:27])
    defparam i22_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1134 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[6] [7]), 
            .I2(n22746), .I3(n43554), .O(n58_adj_3309));   // verilog/coms.v(71[16:27])
    defparam i24_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1135 (.I0(n23337), .I1(\data_out_frame[6] [6]), 
            .I2(n43764), .I3(\data_out_frame[5] [4]), .O(n59_adj_3310));   // verilog/coms.v(71[16:27])
    defparam i25_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1136 (.I0(\data_out_frame[8] [0]), .I1(n43438), 
            .I2(\data_out_frame[8] [2]), .I3(n43355), .O(n57_adj_3311));   // verilog/coms.v(71[16:27])
    defparam i23_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1137 (.I0(n23110), .I1(n43681), .I2(n43864), 
            .I3(n43456), .O(n54_adj_3312));   // verilog/coms.v(71[16:27])
    defparam i20_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n7_adj_3313), .I1(n56_adj_3308), .I2(\data_out_frame[10] [3]), 
            .I3(\data_out_frame[11] [3]), .O(n62));   // verilog/coms.v(71[16:27])
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i32_4_lut (.I0(n57_adj_3311), .I1(n59_adj_3310), .I2(n58_adj_3309), 
            .I3(n60), .O(n66));   // verilog/coms.v(71[16:27])
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1138 (.I0(n43876), .I1(n43340), .I2(n43484), 
            .I3(n22142), .O(n53_adj_3314));   // verilog/coms.v(71[16:27])
    defparam i19_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut_adj_1139 (.I0(n53_adj_3314), .I1(n66), .I2(n62), 
            .I3(n54_adj_3312), .O(n39990));   // verilog/coms.v(71[16:27])
    defparam i33_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(n39990), .I1(n43325), .I2(GND_net), 
            .I3(GND_net), .O(n40119));
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 i936_2_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1692));   // verilog/coms.v(68[16:27])
    defparam i936_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1141 (.I0(n22190), .I1(\data_out_frame[12] [3]), 
            .I2(\data_out_frame[12] [2]), .I3(n23081), .O(n43891));
    defparam i3_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(\data_out_frame[10] [2]), .I1(n43891), 
            .I2(GND_net), .I3(GND_net), .O(n43484));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n43681));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1144 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n43456));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23119));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1146 (.I0(\data_out_frame[6] [0]), .I1(n23119), 
            .I2(n43456), .I3(n6_adj_3222), .O(n22190));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1147 (.I0(\data_out_frame[8] [1]), .I1(n43447), 
            .I2(n23327), .I3(\data_out_frame[6] [1]), .O(n22142));   // verilog/coms.v(70[16:34])
    defparam i3_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_out_frame[10] [3]), .I1(n22142), 
            .I2(GND_net), .I3(GND_net), .O(n43783));
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1149 (.I0(\data_out_frame[12] [4]), .I1(n22190), 
            .I2(\data_out_frame[10] [2]), .I3(GND_net), .O(n43590));
    defparam i2_3_lut_adj_1149.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_1150 (.I0(n43375), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_3315));
    defparam i2_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1151 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(n43681), .I3(\data_out_frame[6] [0]), .O(n14_adj_3316));
    defparam i6_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1152 (.I0(\data_out_frame[14] [5]), .I1(n14_adj_3316), 
            .I2(n10_adj_3315), .I3(\data_out_frame[12] [3]), .O(n43611));
    defparam i7_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1153 (.I0(\data_out_frame[16] [6]), .I1(n22599), 
            .I2(GND_net), .I3(GND_net), .O(n43314));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1153.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1154 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43810));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1154.LUT_INIT = 16'h6666;
    SB_LUT4 i3_2_lut_adj_1155 (.I0(\data_out_frame[13] [3]), .I1(n22599), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3317));   // verilog/coms.v(70[16:42])
    defparam i3_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1156 (.I0(n43786), .I1(n43332), .I2(n43572), 
            .I3(n1713), .O(n22_adj_3318));   // verilog/coms.v(70[16:42])
    defparam i9_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1157 (.I0(n43487), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3319));   // verilog/coms.v(70[16:42])
    defparam i1_2_lut_adj_1157.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1158 (.I0(n49269), .I1(n22_adj_3318), .I2(n16_adj_3317), 
            .I3(n43773), .O(n24_adj_3320));   // verilog/coms.v(70[16:42])
    defparam i11_4_lut_adj_1158.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1159 (.I0(\data_out_frame[14] [0]), .I1(n43419), 
            .I2(n43326), .I3(n14_adj_3319), .O(n23_adj_3321));   // verilog/coms.v(70[16:42])
    defparam i10_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_adj_1160 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_3322));
    defparam i3_2_lut_adj_1160.LUT_INIT = 16'h6666;
    SB_LUT4 i10596_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n24011));
    defparam i10596_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1161 (.I0(n40167), .I1(n1512), .I2(\data_out_frame[15] [1]), 
            .I3(n43400), .O(n22_adj_3323));
    defparam i9_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1162 (.I0(n23_adj_3321), .I1(n43363), .I2(n24_adj_3320), 
            .I3(\data_out_frame[15] [0]), .O(n20_adj_3324));
    defparam i7_4_lut_adj_1162.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_1163 (.I0(\data_out_frame[16] [0]), .I1(n22_adj_3323), 
            .I2(n16_adj_3322), .I3(n43403), .O(n24_adj_3325));
    defparam i11_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1164 (.I0(\data_out_frame[15] [5]), .I1(n24_adj_3325), 
            .I2(n20_adj_3324), .I3(\data_out_frame[13] [5]), .O(n43813));
    defparam i12_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1165 (.I0(n23381), .I1(n43813), .I2(n43810), 
            .I3(n23282), .O(n39781));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1165.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n22809));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1167 (.I0(\data_out_frame[17] [3]), .I1(n22809), 
            .I2(n39781), .I3(\data_out_frame[17] [4]), .O(n43305));
    defparam i3_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1168 (.I0(n43305), .I1(n43688), .I2(n43647), 
            .I3(GND_net), .O(n39404));   // verilog/coms.v(70[16:42])
    defparam i1_3_lut_adj_1168.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1169 (.I0(n39404), .I1(n43623), .I2(n43305), 
            .I3(\data_out_frame[19] [7]), .O(n39844));
    defparam i3_4_lut_adj_1169.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(n39844), .I1(n40144), .I2(GND_net), 
            .I3(GND_net), .O(n43295));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1171 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n43837));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1171.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1172 (.I0(n23085), .I1(\data_out_frame[11] [1]), 
            .I2(\data_out_frame[9] [0]), .I3(n6_adj_3221), .O(n1503));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1173 (.I0(n43522), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[17] [6]), .I3(n43667), .O(n20_adj_3326));   // verilog/coms.v(71[16:27])
    defparam i8_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1174 (.I0(\data_out_frame[18] [0]), .I1(n43818), 
            .I2(\data_out_frame[13] [2]), .I3(\data_out_frame[13] [5]), 
            .O(n19_adj_3327));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1175 (.I0(n43477), .I1(\data_out_frame[15] [6]), 
            .I2(n1503), .I3(\data_out_frame[17] [7]), .O(n21_adj_3328));   // verilog/coms.v(71[16:27])
    defparam i9_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1176 (.I0(n21_adj_3328), .I1(n19_adj_3327), .I2(n20_adj_3326), 
            .I3(GND_net), .O(n43807));   // verilog/coms.v(71[16:27])
    defparam i11_3_lut_adj_1176.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1177 (.I0(\data_out_frame[20] [2]), .I1(n39476), 
            .I2(GND_net), .I3(GND_net), .O(n43409));
    defparam i1_2_lut_adj_1177.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1178 (.I0(\data_out_frame[16] [0]), .I1(n43792), 
            .I2(n43623), .I3(n22146), .O(n40144));
    defparam i3_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43292));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1180 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[11] [2]), .I3(GND_net), .O(n44734));
    defparam i2_3_lut_adj_1180.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1181 (.I0(n23085), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[6] [3]), .I3(n44734), .O(n7_adj_3313));   // verilog/coms.v(68[16:27])
    defparam i2_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1182 (.I0(n7_adj_3313), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[13] [3]), .I3(\data_out_frame[7] [0]), .O(n22596));   // verilog/coms.v(68[16:27])
    defparam i4_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1183 (.I0(\data_out_frame[13] [4]), .I1(n22596), 
            .I2(GND_net), .I3(GND_net), .O(n43522));
    defparam i1_2_lut_adj_1183.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n45299), .I3(n50074), 
            .O(tx_data[7]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i2_3_lut_adj_1184 (.I0(n39281), .I1(n43522), .I2(\data_out_frame[15] [5]), 
            .I3(GND_net), .O(n39504));
    defparam i2_3_lut_adj_1184.LUT_INIT = 16'h9696;
    SB_LUT4 i10597_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43247), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n24012));
    defparam i10597_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_out_frame[17] [7]), .I1(n39504), 
            .I2(GND_net), .I3(GND_net), .O(n40117));
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1186 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3329));
    defparam i1_2_lut_adj_1186.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n45296), .I3(n50080), 
            .O(tx_data[6]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i4_4_lut_adj_1187 (.I0(n40117), .I1(n22972), .I2(n43465), 
            .I3(n6_adj_3329), .O(n39476));
    defparam i4_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1188 (.I0(n39476), .I1(n39470), .I2(GND_net), 
            .I3(GND_net), .O(n22915));
    defparam i1_2_lut_adj_1188.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n23331));
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3330));
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n45293), .I3(n45292), 
            .O(tx_data[5]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i4_4_lut_adj_1191 (.I0(\data_out_frame[5] [0]), .I1(n23331), 
            .I2(\data_out_frame[11] [2]), .I3(n6_adj_3330), .O(n43477));
    defparam i4_4_lut_adj_1191.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1192 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43572));   // verilog/coms.v(94[12:26])
    defparam i1_2_lut_adj_1192.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43400));   // verilog/coms.v(82[17:63])
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1194 (.I0(\data_out_frame[18] [2]), .I1(n23323), 
            .I2(n49269), .I3(n43660), .O(n16_adj_3331));
    defparam i6_4_lut_adj_1194.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1195 (.I0(\data_out_frame[13] [7]), .I1(n43400), 
            .I2(n43572), .I3(n39281), .O(n17_adj_3332));
    defparam i7_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1196 (.I0(n17_adj_3332), .I1(\data_out_frame[11] [5]), 
            .I2(n16_adj_3331), .I3(n43340), .O(n43798));
    defparam i9_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n45284), .I3(n45283), 
            .O(tx_data[3]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n45278), .I3(n45277), 
            .O(tx_data[1]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n45275), .I3(n45274), 
            .O(tx_data[0]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(byte_transmit_counter_c[4]), 
            .I1(byte_transmit_counter_c[3]), .I2(n45281), .I3(n45280), 
            .O(tx_data[2]));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(n22133), .I1(n43498), .I2(GND_net), 
            .I3(GND_net), .O(n22994));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1198 (.I0(n43629), .I1(n22994), .I2(\data_out_frame[16] [0]), 
            .I3(n43798), .O(n10_adj_3216));
    defparam i4_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1199 (.I0(\data_out_frame[20] [5]), .I1(n40171), 
            .I2(n39470), .I3(GND_net), .O(n44472));
    defparam i2_3_lut_adj_1199.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1200 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n43505));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1200.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1201 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23327));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1201.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1202 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[12] [1]), 
            .I2(n43700), .I3(GND_net), .O(n14_adj_3333));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_adj_1202.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1203 (.I0(n43876), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[8] [0]), .I3(n43840), .O(n15_adj_3334));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1204 (.I0(n15_adj_3334), .I1(n43505), .I2(n14_adj_3333), 
            .I3(\data_out_frame[10] [1]), .O(n23381));   // verilog/coms.v(71[16:27])
    defparam i8_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1205 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43363));
    defparam i1_2_lut_adj_1205.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(\data_out_frame[18] [5]), .I1(n23254), 
            .I2(GND_net), .I3(GND_net), .O(n43329));
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1207 (.I0(n23381), .I1(n43346), .I2(GND_net), 
            .I3(GND_net), .O(n1713));
    defparam i1_2_lut_adj_1207.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1208 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n43438));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1208.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1209 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[5][2] ), .I3(GND_net), .O(n43700));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1209.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1210 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[5] [3]), .I3(GND_net), .O(n43764));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1210.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1211 (.I0(\data_out_frame[7] [2]), .I1(n43764), 
            .I2(n43663), .I3(n43468), .O(n23323));
    defparam i3_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1212 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[7] [6]), 
            .I2(n43438), .I3(n6_adj_3335), .O(n23081));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n23110));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n43840));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut_adj_1215 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[12] [0]), 
            .I2(\data_out_frame[11] [5]), .I3(GND_net), .O(n14_adj_3336));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_adj_1215.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1216 (.I0(n43840), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[14] [1]), .O(n15_adj_3337));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1217 (.I0(n15_adj_3337), .I1(\data_out_frame[5] [3]), 
            .I2(n14_adj_3336), .I3(\data_out_frame[7] [5]), .O(n43487));   // verilog/coms.v(70[16:27])
    defparam i8_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1218 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [1]), .I3(GND_net), .O(n43721));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1218.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1219 (.I0(\data_out_frame[13] [7]), .I1(n43721), 
            .I2(n43487), .I3(\data_out_frame[9] [3]), .O(n23254));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1220 (.I0(\data_out_frame[11] [5]), .I1(n43358), 
            .I2(n43703), .I3(n6_adj_3338), .O(n22146));
    defparam i4_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43358));
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_out_frame[5][2] ), .I1(\data_out_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n43663));
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1223 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[7] [4]), .I3(GND_net), .O(n43468));
    defparam i2_3_lut_adj_1223.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n43773));
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1225 (.I0(n43773), .I1(\data_out_frame[7] [0]), 
            .I2(n43412), .I3(\data_out_frame[13] [6]), .O(n14_adj_3339));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1226 (.I0(\data_out_frame[5] [3]), .I1(n14_adj_3339), 
            .I2(n10_adj_3340), .I3(\data_out_frame[13] [7]), .O(n22133));   // verilog/coms.v(70[16:27])
    defparam i7_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1227 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n43818));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_adj_1227.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1228 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23251));
    defparam i1_2_lut_adj_1228.LUT_INIT = 16'h6666;
    SB_LUT4 i33767_2_lut (.I0(n22133), .I1(\data_out_frame[13] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n49269));   // verilog/coms.v(94[12:26])
    defparam i33767_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1229 (.I0(\data_out_frame[7] [1]), .I1(n43667), 
            .I2(n43332), .I3(\data_out_frame[7] [0]), .O(n1512));   // verilog/coms.v(68[16:27])
    defparam i3_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1230 (.I0(n1512), .I1(n49269), .I2(\data_out_frame[15] [7]), 
            .I3(\data_out_frame[13] [5]), .O(n43498));   // verilog/coms.v(94[12:26])
    defparam i3_4_lut_adj_1230.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_out_frame[14] [0]), .I1(n43498), 
            .I2(GND_net), .I3(GND_net), .O(n22972));
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1232 (.I0(n23110), .I1(n23081), .I2(n23323), 
            .I3(\data_out_frame[14] [2]), .O(n43346));
    defparam i3_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1233 (.I0(n22146), .I1(n23254), .I2(\data_out_frame[18] [4]), 
            .I3(\data_out_frame[16] [1]), .O(n12_adj_3341));
    defparam i5_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 n49981_bdd_4_lut (.I0(n49981), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter_c[1]), 
            .O(n49984));
    defparam n49981_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1234 (.I0(n43346), .I1(n12_adj_3341), .I2(\data_out_frame[16] [3]), 
            .I3(n43629), .O(n40171));
    defparam i6_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1235 (.I0(n40171), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [6]), .I3(GND_net), .O(n43397));
    defparam i2_3_lut_adj_1235.LUT_INIT = 16'h6969;
    SB_LUT4 i10319_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10] [0]), 
            .I3(IntegralLimit[0]), .O(n23734));   // verilog/coms.v(248[5:27])
    defparam i10319_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_1236 (.I0(n1713), .I1(n43329), .I2(n22133), .I3(n22984), 
            .O(n22166));
    defparam i3_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i33774_2_lut (.I0(n5024), .I1(n5022), .I2(GND_net), .I3(GND_net), 
            .O(n23557));
    defparam i33774_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1237 (.I0(n22166), .I1(n43397), .I2(GND_net), 
            .I3(GND_net), .O(n43398));
    defparam i1_2_lut_adj_1237.LUT_INIT = 16'h6666;
    SB_LUT4 i10320_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[0] ), .O(n23735));   // verilog/coms.v(248[5:27])
    defparam i10320_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10321_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [0]), 
            .I3(\Ki[0] ), .O(n23736));   // verilog/coms.v(248[5:27])
    defparam i10321_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10322_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [0]), 
            .I3(\Kd[0] ), .O(n23737));   // verilog/coms.v(248[5:27])
    defparam i10322_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10323_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [0]), 
            .I3(gearBoxRatio[0]), .O(n23738));   // verilog/coms.v(248[5:27])
    defparam i10323_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_3_lut_adj_1238 (.I0(n2119), .I1(n744), .I2(n22448), .I3(GND_net), 
            .O(n5_adj_3));
    defparam i1_3_lut_adj_1238.LUT_INIT = 16'haeae;
    SB_LUT4 i10326_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n23741));   // verilog/coms.v(248[5:27])
    defparam i10326_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10327_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [0]), 
            .I3(\PWMLimit[0] ), .O(n23742));   // verilog/coms.v(248[5:27])
    defparam i10327_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34480 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n49975));
    defparam byte_transmit_counter_0__bdd_4_lut_34480.LUT_INIT = 16'he4aa;
    SB_LUT4 i10898_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [0]), 
            .I3(IntegralLimit[8]), .O(n24313));   // verilog/coms.v(248[5:27])
    defparam i10898_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n49975_bdd_4_lut (.I0(n49975), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n49978));
    defparam n49975_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_adj_1239 (.I0(\data_in[0] [3]), .I1(\data_in[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3344));
    defparam i2_2_lut_adj_1239.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1240 (.I0(n7_adj_3344), .I1(n4_c), .I2(n8_adj_3205), 
            .I3(\FRAME_MATCHER.state [1]), .O(\FRAME_MATCHER.state_31__N_1860 [1]));   // verilog/coms.v(92[12:19])
    defparam i1_4_lut_adj_1240.LUT_INIT = 16'hb3a0;
    SB_LUT4 i1_2_lut_adj_1241 (.I0(n737), .I1(\FRAME_MATCHER.state_31__N_1860 [1]), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_1892 [1]));   // verilog/coms.v(92[12:19])
    defparam i1_2_lut_adj_1241.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1242 (.I0(\FRAME_MATCHER.state_31__N_1860 [1]), .I1(n2854), 
            .I2(n44019), .I3(n22454), .O(n6_adj_3345));
    defparam i2_4_lut_adj_1242.LUT_INIT = 16'h0aee;
    SB_LUT4 i3_4_lut_adj_1243 (.I0(n22458), .I1(n6_adj_3345), .I2(\FRAME_MATCHER.state_31__N_1892 [1]), 
            .I3(n22443), .O(n50100));
    defparam i3_4_lut_adj_1243.LUT_INIT = 16'hddfd;
    SB_LUT4 i10899_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10] [7]), 
            .I3(IntegralLimit[7]), .O(n24314));   // verilog/coms.v(248[5:27])
    defparam i10899_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10900_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10][6] ), 
            .I3(IntegralLimit[6]), .O(n24315));   // verilog/coms.v(248[5:27])
    defparam i10900_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10901_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10] [5]), 
            .I3(IntegralLimit[5]), .O(n24316));   // verilog/coms.v(248[5:27])
    defparam i10901_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1244 (.I0(\FRAME_MATCHER.state_31__N_1860 [1]), .I1(n5_adj_3), 
            .I2(GND_net), .I3(GND_net), .O(n42487));
    defparam i1_2_lut_adj_1244.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1245 (.I0(n22451), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state_31__N_1924 [3]), .I3(n44497), .O(n42727));
    defparam i1_4_lut_adj_1245.LUT_INIT = 16'hdc50;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n7_adj_3346), 
            .I2(GND_net), .I3(GND_net), .O(n42493));
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42581));
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1248 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42579));
    defparam i1_2_lut_adj_1248.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\FRAME_MATCHER.state_c [8]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42577));
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1250 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42575));
    defparam i1_2_lut_adj_1250.LUT_INIT = 16'h8888;
    SB_LUT4 i10342_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [0]), 
            .I3(\deadband[0] ), .O(n23757));   // verilog/coms.v(248[5:27])
    defparam i10342_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42573));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42571));
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\FRAME_MATCHER.state_c [12]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42569));
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\FRAME_MATCHER.state_c [13]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42567));
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42565));
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\FRAME_MATCHER.state_c [15]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42563));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1257 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42501));
    defparam i1_2_lut_adj_1257.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\FRAME_MATCHER.state_c [17]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42511));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\FRAME_MATCHER.state_c [18]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42559));
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h8888;
    SB_LUT4 i10862_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [7]), 
            .I3(\Kd[7] ), .O(n24277));   // verilog/coms.v(248[5:27])
    defparam i10862_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10863_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [6]), 
            .I3(\Kd[6] ), .O(n24278));   // verilog/coms.v(248[5:27])
    defparam i10863_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n7_adj_3346), 
            .I2(GND_net), .I3(GND_net), .O(n42557));
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h8888;
    SB_LUT4 i10864_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [5]), 
            .I3(\Kd[5] ), .O(n24279));   // verilog/coms.v(248[5:27])
    defparam i10864_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n7_adj_3346), 
            .I2(GND_net), .I3(GND_net), .O(n42509));
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\FRAME_MATCHER.state_c [21]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42589));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h8888;
    SB_LUT4 i10865_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [4]), 
            .I3(\Kd[4] ), .O(n24280));   // verilog/coms.v(248[5:27])
    defparam i10865_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\FRAME_MATCHER.state_c [22]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42553));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1264 (.I0(n20099), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3348));
    defparam i1_2_lut_adj_1264.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1265 (.I0(\FRAME_MATCHER.state_c [22]), .I1(n2_adj_3124), 
            .I2(n22441), .I3(n4_adj_3348), .O(n42593));
    defparam i1_4_lut_adj_1265.LUT_INIT = 16'h8a88;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42427));
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1267 (.I0(n54), .I1(n37), .I2(n20098), .I3(n43218), 
            .O(n7_adj_3347));
    defparam i1_4_lut_adj_1267.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\FRAME_MATCHER.state_c [24]), .I1(n7_adj_3347), 
            .I2(GND_net), .I3(GND_net), .O(n42555));
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1269 (.I0(\data_in_frame[9] [5]), .I1(n43299), 
            .I2(n22953), .I3(\data_in_frame[7] [4]), .O(n39500));
    defparam i1_2_lut_3_lut_4_lut_adj_1269.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1270 (.I0(\FRAME_MATCHER.state_c [25]), .I1(n44479), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3129));
    defparam i1_2_lut_adj_1270.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1271 (.I0(\FRAME_MATCHER.state_c [26]), .I1(n7_adj_3346), 
            .I2(GND_net), .I3(GND_net), .O(n42507));
    defparam i1_2_lut_adj_1271.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1272 (.I0(n22453), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n43218));
    defparam i2_3_lut_adj_1272.LUT_INIT = 16'h4040;
    SB_LUT4 i2_4_lut_adj_1273 (.I0(n37), .I1(n20125), .I2(n54), .I3(n43218), 
            .O(n7_adj_3346));
    defparam i2_4_lut_adj_1273.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_adj_1274 (.I0(\FRAME_MATCHER.state_c [27]), .I1(n7_adj_3346), 
            .I2(GND_net), .I3(GND_net), .O(n42519));
    defparam i1_2_lut_adj_1274.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(n20136), .I1(n2854), .I2(GND_net), 
            .I3(GND_net), .O(n20125));
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h2222;
    SB_LUT4 i5_2_lut_3_lut_4_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[14] [4]), 
            .I2(\data_in_frame[14]_c [3]), .I3(\data_in_frame[11] [7]), 
            .O(n15_adj_3139));
    defparam i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(\FRAME_MATCHER.state_c [28]), .I1(n44479), 
            .I2(GND_net), .I3(GND_net), .O(n42481));
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1277 (.I0(n20098), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n22453), .O(n44728));
    defparam i3_4_lut_adj_1277.LUT_INIT = 16'h0080;
    SB_LUT4 i1_4_lut_adj_1278 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n44574), 
            .I2(n44728), .I3(n54), .O(n42551));
    defparam i1_4_lut_adj_1278.LUT_INIT = 16'haaa8;
    SB_LUT4 i10891_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [7]), 
            .I3(IntegralLimit[15]), .O(n24306));   // verilog/coms.v(248[5:27])
    defparam i10891_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1279 (.I0(n22343), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_3349));
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'heeee;
    SB_LUT4 i15033_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_3349), .I3(\FRAME_MATCHER.i [1]), .O(n737));   // verilog/coms.v(152[9:60])
    defparam i15033_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(\FRAME_MATCHER.state [1]), .I1(n22441), 
            .I2(GND_net), .I3(GND_net), .O(n22443));   // verilog/coms.v(147[5:27])
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1281 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[3] [3]), .O(n6_adj_3213));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i10866_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [3]), 
            .I3(\Kd[3] ), .O(n24281));   // verilog/coms.v(248[5:27])
    defparam i10866_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_1282 (.I0(n22456), .I1(n44009), .I2(\FRAME_MATCHER.state [0]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n22458));   // verilog/coms.v(190[5:24])
    defparam i3_4_lut_adj_1282.LUT_INIT = 16'hfeff;
    SB_LUT4 i10867_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [2]), 
            .I3(\Kd[2] ), .O(n24282));   // verilog/coms.v(248[5:27])
    defparam i10867_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10868_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[4] [1]), 
            .I3(\Kd[1] ), .O(n24283));   // verilog/coms.v(248[5:27])
    defparam i10868_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i4_4_lut_adj_1283 (.I0(n22448), .I1(n28434), .I2(n22458), 
            .I3(n22451), .O(n10_adj_3350));
    defparam i4_4_lut_adj_1283.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1284 (.I0(\FRAME_MATCHER.state [0]), .I1(n10_adj_3350), 
            .I2(n63_adj_3342), .I3(n22447), .O(n2119));
    defparam i5_4_lut_adj_1284.LUT_INIT = 16'hc080;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(n20136), .I1(n2119), .I2(GND_net), 
            .I3(GND_net), .O(n54));   // verilog/coms.v(244[6] 246[9])
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'h8888;
    SB_LUT4 i77_2_lut (.I0(n22454), .I1(n20098), .I2(GND_net), .I3(GND_net), 
            .O(n59));   // verilog/coms.v(112[11:12])
    defparam i77_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i5_4_lut_adj_1286 (.I0(\data_in[2] [3]), .I1(\data_in[3][5] ), 
            .I2(n27228), .I3(\data_in[0] [2]), .O(n12_adj_3351));
    defparam i5_4_lut_adj_1286.LUT_INIT = 16'h0800;
    SB_LUT4 i1_4_lut_adj_1287 (.I0(\data_in[0]_c [7]), .I1(n31), .I2(n12_adj_3351), 
            .I3(n8_adj_3352), .O(n4_c));
    defparam i1_4_lut_adj_1287.LUT_INIT = 16'h7333;
    SB_LUT4 i4_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [14]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3353));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1288 (.I0(\FRAME_MATCHER.i [16]), .I1(\FRAME_MATCHER.i [9]), 
            .I2(\FRAME_MATCHER.i [19]), .I3(\FRAME_MATCHER.i [13]), .O(n36));
    defparam i14_4_lut_adj_1288.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1289 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [10]), .O(n44869));
    defparam i3_4_lut_adj_1289.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1290 (.I0(\FRAME_MATCHER.i [18]), .I1(\FRAME_MATCHER.i [7]), 
            .I2(n44869), .I3(\FRAME_MATCHER.i [22]), .O(n34));
    defparam i12_4_lut_adj_1290.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1291 (.I0(\FRAME_MATCHER.i [20]), .I1(n36), .I2(n26_adj_3353), 
            .I3(\FRAME_MATCHER.i [15]), .O(n40));
    defparam i18_4_lut_adj_1291.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1292 (.I0(\FRAME_MATCHER.i [25]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(\FRAME_MATCHER.i [28]), .I3(\FRAME_MATCHER.i [6]), .O(n38_adj_3354));
    defparam i16_4_lut_adj_1292.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n34), .I2(\FRAME_MATCHER.i [29]), 
            .I3(GND_net), .O(n39_adj_3355));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1293 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [23]), .O(n37_adj_3356));
    defparam i15_4_lut_adj_1293.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1294 (.I0(n37_adj_3356), .I1(n39_adj_3355), .I2(n38_adj_3354), 
            .I3(n40), .O(n22501));
    defparam i21_4_lut_adj_1294.LUT_INIT = 16'hfffe;
    SB_LUT4 i15041_4_lut (.I0(n10_adj_3121), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n22501), .O(n3758));   // verilog/coms.v(244[9:58])
    defparam i15041_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i10869_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [7]), 
            .I3(\Ki[7] ), .O(n24284));   // verilog/coms.v(248[5:27])
    defparam i10869_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1295 (.I0(\data_in[3] [1]), .I1(\data_in[3][3] ), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_3357));   // verilog/coms.v(125[12] 284[6])
    defparam i1_2_lut_adj_1295.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1296 (.I0(\data_in[0] [6]), .I1(\data_in[0] [3]), 
            .I2(\data_in[1] [0]), .I3(\data_in[3] [0]), .O(n10_adj_3208));
    defparam i3_4_lut_adj_1296.LUT_INIT = 16'hbfff;
    SB_LUT4 i4_4_lut_adj_1297 (.I0(\data_in[2] [2]), .I1(\data_in[1][5] ), 
            .I2(\data_in[1][4] ), .I3(n6_adj_3358), .O(n139));
    defparam i4_4_lut_adj_1297.LUT_INIT = 16'hfff7;
    SB_LUT4 i2_2_lut_adj_1298 (.I0(\data_in[0] [2]), .I1(\data_in[0]_c [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3359));
    defparam i2_2_lut_adj_1298.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_1299 (.I0(\data_in[3][5] ), .I1(\data_in[3] [1]), 
            .I2(\data_in[2][1] ), .I3(\data_in[3][3] ), .O(n44946));   // verilog/coms.v(137[7:80])
    defparam i3_4_lut_adj_1299.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1300 (.I0(n44946), .I1(\data_in[2] [3]), .I2(n6_adj_3359), 
            .I3(\data_in[3] [6]), .O(n22475));   // verilog/coms.v(137[7:80])
    defparam i7_4_lut_adj_1300.LUT_INIT = 16'hfeff;
    SB_LUT4 i4_4_lut_adj_1301 (.I0(\data_in[1] [7]), .I1(\data_in[0]_c [0]), 
            .I2(\data_in[1][1] ), .I3(\data_in[0] [4]), .O(n10_adj_3360));
    defparam i4_4_lut_adj_1301.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1302 (.I0(\data_in[3][4] ), .I1(n10_adj_3360), 
            .I2(\data_in[2]_c [7]), .I3(GND_net), .O(n22564));
    defparam i5_3_lut_adj_1302.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_1303 (.I0(\data_in[1][3] ), .I1(\data_in[0] [1]), 
            .I2(\data_in[3][2] ), .I3(\data_in[0] [5]), .O(n16_adj_3361));
    defparam i6_4_lut_adj_1303.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1304 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2]_c [0]), .I3(\data_in[1][2] ), .O(n17_adj_3362));
    defparam i7_4_lut_adj_1304.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1305 (.I0(n17_adj_3362), .I1(\data_in[1][6] ), 
            .I2(n16_adj_3361), .I3(\data_in[3][7] ), .O(n22432));
    defparam i9_4_lut_adj_1305.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_2_lut_adj_1306 (.I0(n22432), .I1(\data_in[2] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3363));
    defparam i2_2_lut_adj_1306.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1307 (.I0(n22564), .I1(\data_in[0] [3]), .I2(\data_in[0] [6]), 
            .I3(\data_in[2] [4]), .O(n14_adj_3364));
    defparam i6_4_lut_adj_1307.LUT_INIT = 16'hefff;
    SB_LUT4 i7_4_lut_adj_1308 (.I0(\data_in[1][4] ), .I1(n14_adj_3364), 
            .I2(n10_adj_3363), .I3(\data_in[1][5] ), .O(n45152));
    defparam i7_4_lut_adj_1308.LUT_INIT = 16'hfffd;
    SB_LUT4 i3_4_lut_adj_1309 (.I0(\data_in[1] [0]), .I1(n22475), .I2(n45152), 
            .I3(\data_in[3] [0]), .O(n31));   // verilog/coms.v(125[12] 284[6])
    defparam i3_4_lut_adj_1309.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(n22475), .I1(\data_in[3][7] ), .I2(GND_net), 
            .I3(GND_net), .O(n12_adj_3365));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1311 (.I0(\data_in[2] [6]), .I1(\data_in[1][6] ), 
            .I2(\data_in[0] [1]), .I3(\data_in[1][3] ), .O(n18_adj_3366));
    defparam i7_4_lut_adj_1311.LUT_INIT = 16'hefff;
    SB_LUT4 i29754_4_lut (.I0(\data_in[2]_c [0]), .I1(\data_in[2] [5]), 
            .I2(\data_in[1][2] ), .I3(\data_in[3][2] ), .O(n45254));
    defparam i29754_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut_adj_1312 (.I0(n45254), .I1(\data_in[0] [5]), .I2(n18_adj_3366), 
            .I3(n12_adj_3365), .O(n43263));
    defparam i10_4_lut_adj_1312.LUT_INIT = 16'hfff7;
    SB_LUT4 i5_4_lut_adj_1313 (.I0(\data_in[0]_c [7]), .I1(n15_adj_3357), 
            .I2(\data_in[2][1] ), .I3(\data_in[2] [3]), .O(n12_adj_3367));
    defparam i5_4_lut_adj_1313.LUT_INIT = 16'hbfff;
    SB_LUT4 i6_4_lut_adj_1314 (.I0(\data_in[3][5] ), .I1(n12_adj_3367), 
            .I2(\data_in[0] [2]), .I3(n27228), .O(n63));
    defparam i6_4_lut_adj_1314.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_adj_1315 (.I0(n139), .I1(n10_adj_3208), .I2(GND_net), 
            .I3(GND_net), .O(n25797));   // verilog/coms.v(125[12] 284[6])
    defparam i1_2_lut_adj_1315.LUT_INIT = 16'heeee;
    SB_LUT4 i31518_2_lut (.I0(byte_transmit_counter_c[2]), .I1(byte_transmit_counter_c[1]), 
            .I2(GND_net), .I3(GND_net), .O(n47022));
    defparam i31518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_1316 (.I0(byte_transmit_counter_c[5]), .I1(byte_transmit_counter_c[6]), 
            .I2(byte_transmit_counter_c[7]), .I3(n21_adj_3368), .O(n7_adj_3203));   // verilog/coms.v(99[12:33])
    defparam i3_4_lut_adj_1316.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1317 (.I0(n25797), .I1(n63), .I2(n43263), .I3(n31), 
            .O(n20136));
    defparam i2_4_lut_adj_1317.LUT_INIT = 16'hc800;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\FRAME_MATCHER.state [0]), .I1(n22447), 
            .I2(GND_net), .I3(GND_net), .O(n22448));   // verilog/coms.v(201[5:16])
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'hdddd;
    SB_LUT4 i10902_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10] [4]), 
            .I3(IntegralLimit[4]), .O(n24317));   // verilog/coms.v(248[5:27])
    defparam i10902_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(\FRAME_MATCHER.state [1]), .I1(n22441), 
            .I2(GND_net), .I3(GND_net), .O(n22442));   // verilog/coms.v(239[5:25])
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'hdddd;
    SB_LUT4 i10903_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10] [3]), 
            .I3(IntegralLimit[3]), .O(n24318));   // verilog/coms.v(248[5:27])
    defparam i10903_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10904_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10] [2]), 
            .I3(IntegralLimit[2]), .O(n24319));   // verilog/coms.v(248[5:27])
    defparam i10904_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10905_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[10] [1]), 
            .I3(IntegralLimit[1]), .O(n24320));   // verilog/coms.v(248[5:27])
    defparam i10905_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10870_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [6]), 
            .I3(\Ki[6] ), .O(n24285));   // verilog/coms.v(248[5:27])
    defparam i10870_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10871_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [5]), 
            .I3(\Ki[5] ), .O(n24286));   // verilog/coms.v(248[5:27])
    defparam i10871_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10872_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [4]), 
            .I3(\Ki[4] ), .O(n24287));   // verilog/coms.v(248[5:27])
    defparam i10872_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10873_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [3]), 
            .I3(\Ki[3] ), .O(n24288));   // verilog/coms.v(248[5:27])
    defparam i10873_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(n29726), .I1(n23829), .I2(GND_net), 
            .I3(GND_net), .O(n75));   // verilog/coms.v(109[11:16])
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h8888;
    SB_LUT4 i10874_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [2]), 
            .I3(\Ki[2] ), .O(n24289));   // verilog/coms.v(248[5:27])
    defparam i10874_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10486_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[6] [1]), 
            .I3(\PWMLimit[9] ), .O(n23901));   // verilog/coms.v(248[5:27])
    defparam i10486_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10487_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[6] [0]), 
            .I3(\PWMLimit[8] ), .O(n23902));   // verilog/coms.v(248[5:27])
    defparam i10487_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14699_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [7]), 
            .I3(\PWMLimit[7] ), .O(n23903));   // verilog/coms.v(248[5:27])
    defparam i14699_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14661_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [6]), 
            .I3(\PWMLimit[6] ), .O(n28060));   // verilog/coms.v(248[5:27])
    defparam i14661_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14606_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [5]), 
            .I3(\PWMLimit[5] ), .O(n23905));   // verilog/coms.v(248[5:27])
    defparam i14606_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10491_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [4]), 
            .I3(\PWMLimit[4] ), .O(n23906));   // verilog/coms.v(248[5:27])
    defparam i10491_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10492_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [3]), 
            .I3(\PWMLimit[3] ), .O(n23907));   // verilog/coms.v(248[5:27])
    defparam i10492_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10493_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [2]), 
            .I3(\PWMLimit[2] ), .O(n23908));   // verilog/coms.v(248[5:27])
    defparam i10493_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10494_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[7] [1]), 
            .I3(\PWMLimit[1] ), .O(n23909));   // verilog/coms.v(248[5:27])
    defparam i10494_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10495_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n23910));   // verilog/coms.v(248[5:27])
    defparam i10495_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10892_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [6]), 
            .I3(IntegralLimit[14]), .O(n24307));   // verilog/coms.v(248[5:27])
    defparam i10892_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10893_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [5]), 
            .I3(IntegralLimit[13]), .O(n24308));   // verilog/coms.v(248[5:27])
    defparam i10893_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10501_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n23916));   // verilog/coms.v(248[5:27])
    defparam i10501_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10500_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n23915));   // verilog/coms.v(248[5:27])
    defparam i10500_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i29845_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45345));
    defparam i29845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29846_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45346));
    defparam i29846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29849_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45349));
    defparam i29849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29848_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45348));
    defparam i29848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29839_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45339));
    defparam i29839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29840_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45340));
    defparam i29840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29843_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45343));
    defparam i29843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29842_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45342));
    defparam i29842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32165_2_lut (.I0(\data_out_frame[5] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n47217));
    defparam i32165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_3122));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32158_2_lut (.I0(\data_out_frame[22] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n47245));
    defparam i32158_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19));   // verilog/coms.v(103[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n22447), 
            .I2(n20136), .I3(n744), .O(n2_adj_3124));   // verilog/coms.v(201[5:16])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h2000;
    SB_LUT4 i1_3_lut_4_lut_adj_1321 (.I0(byte_transmit_counter_c[4]), .I1(byte_transmit_counter_c[2]), 
            .I2(byte_transmit_counter_c[1]), .I3(byte_transmit_counter_c[3]), 
            .O(n21_adj_3368));   // verilog/coms.v(99[12:33])
    defparam i1_3_lut_4_lut_adj_1321.LUT_INIT = 16'haa80;
    SB_LUT4 i10499_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n23914));   // verilog/coms.v(248[5:27])
    defparam i10499_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10498_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1][4] ), 
            .I3(control_mode[4]), .O(n23913));   // verilog/coms.v(248[5:27])
    defparam i10498_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10497_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n23912));   // verilog/coms.v(248[5:27])
    defparam i10497_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10496_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n23911));   // verilog/coms.v(248[5:27])
    defparam i10496_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_4_lut_adj_1322 (.I0(\data_in[3][4] ), .I1(n10_adj_3360), 
            .I2(\data_in[2]_c [7]), .I3(\data_in[2] [4]), .O(n6_adj_3358));
    defparam i1_2_lut_4_lut_adj_1322.LUT_INIT = 16'hffdf;
    SB_LUT4 i2_3_lut_4_lut_adj_1323 (.I0(\data_in[3] [6]), .I1(n139), .I2(n10_adj_3208), 
            .I3(n22432), .O(n27228));
    defparam i2_3_lut_4_lut_adj_1323.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1324 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n22456), .O(n22447));
    defparam i2_3_lut_4_lut_adj_1324.LUT_INIT = 16'hfff7;
    SB_LUT4 i10849_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18] [5]), 
            .I3(gearBoxRatio[13]), .O(n24264));   // verilog/coms.v(248[5:27])
    defparam i10849_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_adj_1325 (.I0(n29726), .I1(n23826), .I2(GND_net), 
            .I3(GND_net), .O(n23828));   // verilog/coms.v(109[11:16])
    defparam i1_2_lut_adj_1325.LUT_INIT = 16'h8888;
    SB_LUT4 i10850_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18] [4]), 
            .I3(gearBoxRatio[12]), .O(n24265));   // verilog/coms.v(248[5:27])
    defparam i10850_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10851_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18] [3]), 
            .I3(gearBoxRatio[11]), .O(n24266));   // verilog/coms.v(248[5:27])
    defparam i10851_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10852_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18][2] ), 
            .I3(gearBoxRatio[10]), .O(n24267));   // verilog/coms.v(248[5:27])
    defparam i10852_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10853_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18] [1]), 
            .I3(gearBoxRatio[9]), .O(n24268));   // verilog/coms.v(248[5:27])
    defparam i10853_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10854_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18][0] ), 
            .I3(gearBoxRatio[8]), .O(n24269));   // verilog/coms.v(248[5:27])
    defparam i10854_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10855_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [7]), 
            .I3(gearBoxRatio[7]), .O(n24270));   // verilog/coms.v(248[5:27])
    defparam i10855_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10856_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [6]), 
            .I3(gearBoxRatio[6]), .O(n24271));   // verilog/coms.v(248[5:27])
    defparam i10856_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10857_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [5]), 
            .I3(gearBoxRatio[5]), .O(n24272));   // verilog/coms.v(248[5:27])
    defparam i10857_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34475 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter_c[1]), .O(n49969));
    defparam byte_transmit_counter_0__bdd_4_lut_34475.LUT_INIT = 16'he4aa;
    SB_LUT4 i10847_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18] [7]), 
            .I3(gearBoxRatio[15]), .O(n24262));   // verilog/coms.v(248[5:27])
    defparam i10847_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10848_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[18] [6]), 
            .I3(gearBoxRatio[14]), .O(n24263));   // verilog/coms.v(248[5:27])
    defparam i10848_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10846_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [0]), 
            .I3(gearBoxRatio[16]), .O(n24261));   // verilog/coms.v(248[5:27])
    defparam i10846_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10861_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [1]), 
            .I3(gearBoxRatio[1]), .O(n24276));   // verilog/coms.v(248[5:27])
    defparam i10861_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10860_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [2]), 
            .I3(gearBoxRatio[2]), .O(n24275));   // verilog/coms.v(248[5:27])
    defparam i10860_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10859_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [3]), 
            .I3(gearBoxRatio[3]), .O(n24274));   // verilog/coms.v(248[5:27])
    defparam i10859_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1326 (.I0(\data_in[2][1] ), .I1(\data_in[3] [1]), 
            .I2(\data_in[3][3] ), .I3(GND_net), .O(n8_adj_3352));
    defparam i1_2_lut_3_lut_adj_1326.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_1327 (.I0(\FRAME_MATCHER.state [1]), .I1(n22441), 
            .I2(n20136), .I3(n3758), .O(n42));   // verilog/coms.v(112[11:12])
    defparam i1_3_lut_4_lut_adj_1327.LUT_INIT = 16'h0020;
    SB_LUT4 i1_3_lut_4_lut_adj_1328 (.I0(n20136), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n22441), .I3(n737), .O(n37));   // verilog/coms.v(147[5:27])
    defparam i1_3_lut_4_lut_adj_1328.LUT_INIT = 16'h0002;
    SB_LUT4 i1_3_lut_4_lut_adj_1329 (.I0(\FRAME_MATCHER.state [3]), .I1(n20136), 
            .I2(n2119), .I3(n42), .O(n42491));
    defparam i1_3_lut_4_lut_adj_1329.LUT_INIT = 16'haa80;
    SB_LUT4 i10858_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[19] [4]), 
            .I3(gearBoxRatio[4]), .O(n24273));   // verilog/coms.v(248[5:27])
    defparam i10858_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i28523_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(n22441), 
            .I2(n3758), .I3(GND_net), .O(n44019));
    defparam i28523_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1330 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[14] [0]), 
            .I2(n43498), .I3(GND_net), .O(n43629));
    defparam i1_2_lut_3_lut_adj_1330.LUT_INIT = 16'h9696;
    SB_LUT4 i10999_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [2]), 
            .I3(\deadband[2] ), .O(n24414));   // verilog/coms.v(248[5:27])
    defparam i10999_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11000_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [3]), 
            .I3(\deadband[3] ), .O(n24415));   // verilog/coms.v(248[5:27])
    defparam i11000_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11001_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [4]), 
            .I3(\deadband[4] ), .O(n24416));   // verilog/coms.v(248[5:27])
    defparam i11001_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14607_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [5]), 
            .I3(\deadband[5] ), .O(n24417));   // verilog/coms.v(248[5:27])
    defparam i14607_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14656_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [6]), 
            .I3(\deadband[6] ), .O(n24418));   // verilog/coms.v(248[5:27])
    defparam i14656_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14704_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [7]), 
            .I3(\deadband[7] ), .O(n24419));   // verilog/coms.v(248[5:27])
    defparam i14704_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11005_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[12] [0]), 
            .I3(\deadband[8] ), .O(n24420));   // verilog/coms.v(248[5:27])
    defparam i11005_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i11006_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[12] [1]), 
            .I3(\deadband[9] ), .O(n24421));   // verilog/coms.v(248[5:27])
    defparam i11006_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10839_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [7]), 
            .I3(gearBoxRatio[23]), .O(n24254));   // verilog/coms.v(248[5:27])
    defparam i10839_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n43667));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1332 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(n43818), .I3(GND_net), .O(n43332));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1332.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1333 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[5][2] ), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[6] [7]), .O(n10_adj_3340));   // verilog/coms.v(70[16:27])
    defparam i2_2_lut_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1334 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[9] [5]), .I3(\data_out_frame[7] [4]), .O(n43412));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1335 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[5][2] ), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n43660));
    defparam i1_2_lut_3_lut_adj_1335.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1336 (.I0(\data_out_frame[5][2] ), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[6] [6]), .I3(\data_out_frame[9] [2]), .O(n6_adj_3338));
    defparam i1_2_lut_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1337 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[5][2] ), .O(n6_adj_3335));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1338 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[16] [2]), .I3(\data_out_frame[18] [4]), 
            .O(n22984));
    defparam i2_3_lut_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n43876));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(n43721), .I3(GND_net), .O(n43340));
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1341 (.I0(n22133), .I1(n43498), .I2(\data_out_frame[18] [1]), 
            .I3(n43798), .O(n43465));
    defparam i1_2_lut_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(n22133), .I1(n43498), .I2(\data_out_frame[18] [1]), 
            .I3(GND_net), .O(n43792));
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n23085));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1344 (.I0(n40144), .I1(\data_out_frame[20] [2]), 
            .I2(n39476), .I3(GND_net), .O(n43410));
    defparam i1_2_lut_3_lut_adj_1344.LUT_INIT = 16'h9696;
    SB_LUT4 i10840_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [6]), 
            .I3(gearBoxRatio[22]), .O(n24255));   // verilog/coms.v(248[5:27])
    defparam i10840_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1345 (.I0(\data_out_frame[17] [7]), .I1(n39504), 
            .I2(n43807), .I3(GND_net), .O(n43623));
    defparam i1_2_lut_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i10841_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [5]), 
            .I3(gearBoxRatio[21]), .O(n24256));   // verilog/coms.v(248[5:27])
    defparam i10841_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10842_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [4]), 
            .I3(gearBoxRatio[20]), .O(n24257));   // verilog/coms.v(248[5:27])
    defparam i10842_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_4_lut_adj_1346 (.I0(\data_out_frame[20] [2]), .I1(n39844), 
            .I2(n40144), .I3(\data_out_frame[20] [1]), .O(n44636));
    defparam i2_3_lut_4_lut_adj_1346.LUT_INIT = 16'h9669;
    SB_LUT4 i10843_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [3]), 
            .I3(gearBoxRatio[19]), .O(n24258));   // verilog/coms.v(248[5:27])
    defparam i10843_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10844_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [2]), 
            .I3(gearBoxRatio[18]), .O(n24259));   // verilog/coms.v(248[5:27])
    defparam i10844_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n49969_bdd_4_lut (.I0(n49969), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter_c[1]), 
            .O(n49972));
    defparam n49969_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10845_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[17] [1]), 
            .I3(gearBoxRatio[17]), .O(n24260));   // verilog/coms.v(248[5:27])
    defparam i10845_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_34470 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter_c[1]), .O(n49963));
    defparam byte_transmit_counter_0__bdd_4_lut_34470.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[16] [6]), 
            .I2(n22599), .I3(GND_net), .O(n23282));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n43447));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1349 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[14] [6]), 
            .I2(n39990), .I3(n43325), .O(n43786));
    defparam i1_2_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i26_3_lut_4_lut (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [7]), 
            .I2(n52_adj_3307), .I3(\data_out_frame[5][2] ), .O(n60));   // verilog/coms.v(71[16:27])
    defparam i26_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1350 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[12] [7]), 
            .I2(n43861), .I3(GND_net), .O(n6_adj_3306));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1350.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(n44973), .I1(n22126), .I2(n43638), 
            .I3(GND_net), .O(n43283));
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(\data_out_frame[19] [6]), .I1(\data_out_frame[19] [5]), 
            .I2(n43638), .I3(GND_net), .O(n6_adj_3293));
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 i10883_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [7]), 
            .I3(IntegralLimit[23]), .O(n24298));   // verilog/coms.v(248[5:27])
    defparam i10883_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_3_lut_4_lut_adj_1353 (.I0(n23405), .I1(\data_out_frame[17] [4]), 
            .I2(n10_adj_3290), .I3(\data_out_frame[19] [5]), .O(n44400));
    defparam i5_3_lut_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i10884_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [6]), 
            .I3(IntegralLimit[22]), .O(n24299));   // verilog/coms.v(248[5:27])
    defparam i10884_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 n49963_bdd_4_lut (.I0(n49963), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter_c[1]), 
            .O(n49966));
    defparam n49963_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n44238));   // verilog/coms.v(109[11:16])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i10885_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [5]), 
            .I3(IntegralLimit[21]), .O(n24300));   // verilog/coms.v(248[5:27])
    defparam i10885_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10886_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [4]), 
            .I3(IntegralLimit[20]), .O(n24301));   // verilog/coms.v(248[5:27])
    defparam i10886_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10887_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [3]), 
            .I3(IntegralLimit[19]), .O(n24302));   // verilog/coms.v(248[5:27])
    defparam i10887_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10888_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [2]), 
            .I3(IntegralLimit[18]), .O(n24303));   // verilog/coms.v(248[5:27])
    defparam i10888_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10998_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[13] [1]), 
            .I3(\deadband[1] ), .O(n24413));   // verilog/coms.v(248[5:27])
    defparam i10998_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10878_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[5] ), .O(n24293));   // verilog/coms.v(248[5:27])
    defparam i10878_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10879_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[4] ), .O(n24294));   // verilog/coms.v(248[5:27])
    defparam i10879_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10880_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[3] ), .O(n24295));   // verilog/coms.v(248[5:27])
    defparam i10880_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_4_lut_adj_1354 (.I0(\FRAME_MATCHER.state [0]), .I1(n28723), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n44009), .O(n5024));
    defparam i2_3_lut_4_lut_adj_1354.LUT_INIT = 16'h0100;
    SB_LUT4 i10890_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [0]), 
            .I3(IntegralLimit[16]), .O(n24305));   // verilog/coms.v(248[5:27])
    defparam i10890_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10895_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [3]), 
            .I3(IntegralLimit[11]), .O(n24310));   // verilog/coms.v(248[5:27])
    defparam i10895_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10896_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [2]), 
            .I3(IntegralLimit[10]), .O(n24311));   // verilog/coms.v(248[5:27])
    defparam i10896_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10897_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [1]), 
            .I3(IntegralLimit[9]), .O(n24312));   // verilog/coms.v(248[5:27])
    defparam i10897_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10881_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[2] ), .O(n24296));   // verilog/coms.v(248[5:27])
    defparam i10881_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10882_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[1] ), .O(n24297));   // verilog/coms.v(248[5:27])
    defparam i10882_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10894_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[9] [4]), 
            .I3(IntegralLimit[12]), .O(n24309));   // verilog/coms.v(248[5:27])
    defparam i10894_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10875_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[3] [1]), 
            .I3(\Ki[1] ), .O(n24290));   // verilog/coms.v(248[5:27])
    defparam i10875_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10876_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[7] ), .O(n24291));   // verilog/coms.v(248[5:27])
    defparam i10876_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i10877_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[6] ), .O(n24292));   // verilog/coms.v(248[5:27])
    defparam i10877_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i1_2_lut_3_lut_adj_1355 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[6] [6]), 
            .I2(n22801), .I3(GND_net), .O(n43388));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_3_lut_adj_1355.LUT_INIT = 16'h9696;
    SB_LUT4 i10889_3_lut_4_lut (.I0(n63_adj_3342), .I1(n29738), .I2(\data_in_frame[8] [1]), 
            .I3(IntegralLimit[17]), .O(n24304));   // verilog/coms.v(248[5:27])
    defparam i10889_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_3_lut_4_lut_adj_1356 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[15] [4]), .O(n43870));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1357 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [4]), 
            .I2(\data_in_frame[19] [6]), .I3(n23346), .O(n43528));
    defparam i2_3_lut_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1358 (.I0(\data_in_frame[8] [7]), .I1(n23385), 
            .I2(\data_in_frame[7] [1]), .I3(\data_in_frame[6] [7]), .O(n14_adj_3243));
    defparam i5_3_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1359 (.I0(\data_in_frame[1][4] ), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[1] [2]), .O(n43780));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(n10_adj_3116), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[8] [3]), .I3(GND_net), .O(n43490));   // verilog/coms.v(69[16:41])
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1361 (.I0(n10_adj_3116), .I1(\data_in_frame[6] [2]), 
            .I2(n23367), .I3(\data_in_frame[8] [4]), .O(n43367));   // verilog/coms.v(69[16:41])
    defparam i2_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i10325_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n23740));
    defparam i10325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10670_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n24085));
    defparam i10670_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10671_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n24086));
    defparam i10671_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10672_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n24087));
    defparam i10672_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10673_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n24088));
    defparam i10673_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10674_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n24089));
    defparam i10674_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10675_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n24090));
    defparam i10675_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1362 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[1] [0]), .O(n18_adj_3241));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 i10676_3_lut_4_lut (.I0(n8_adj_3212), .I1(n43226), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n24091));
    defparam i10676_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1363 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n28284), .O(n43247));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_1363.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n21061));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1365 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n28284), .O(n43226));   // verilog/coms.v(149[7:23])
    defparam i2_3_lut_4_lut_adj_1365.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_59_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3235));   // verilog/coms.v(149[7:23])
    defparam equal_59_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_3_lut_4_lut_adj_1366 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [0]), .O(n23468));   // verilog/coms.v(68[16:69])
    defparam i2_3_lut_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 equal_60_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3212));   // verilog/coms.v(149[7:23])
    defparam equal_60_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[13] [1]), .I3(n43821), .O(n43678));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n43655));   // verilog/coms.v(225[9:81])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n43378));   // verilog/coms.v(70[16:34])
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1370 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[1] [7]), 
            .I2(n43318), .I3(\data_in_frame[4] [3]), .O(n22796));   // verilog/coms.v(225[9:81])
    defparam i2_3_lut_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1371 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(n23176), .I3(\data_in_frame[8] [6]), .O(n43544));   // verilog/coms.v(71[16:43])
    defparam i2_3_lut_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1372 (.I0(\data_in_frame[6] [7]), .I1(n5_adj_3218), 
            .I2(n23358), .I3(GND_net), .O(n6_adj_3240));   // verilog/coms.v(71[16:43])
    defparam i1_2_lut_3_lut_adj_1372.LUT_INIT = 16'h9696;
    SB_LUT4 i10662_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n24077));
    defparam i10662_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1373 (.I0(\data_in_frame[15] [5]), .I1(n43873), 
            .I2(n43879), .I3(\data_in_frame[16] [5]), .O(n40161));
    defparam i1_2_lut_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[14]_c [3]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n43846));
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1375 (.I0(n16), .I1(\data_in_frame[7] [3]), 
            .I2(n39466), .I3(GND_net), .O(n43299));
    defparam i1_2_lut_3_lut_adj_1375.LUT_INIT = 16'h6969;
    SB_LUT4 equal_1044_i16_2_lut_4_lut (.I0(n23358), .I1(n43415), .I2(n23468), 
            .I3(\data_in_frame[4] [7]), .O(n16));   // verilog/coms.v(225[9:81])
    defparam equal_1044_i16_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1376 (.I0(n22771), .I1(\data_out_frame[10] [3]), 
            .I2(n22142), .I3(\data_out_frame[12] [5]), .O(n43325));
    defparam i1_2_lut_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i10663_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n24078));
    defparam i10663_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1377 (.I0(n43590), .I1(\data_out_frame[10] [3]), 
            .I2(n22142), .I3(n43611), .O(n40167));
    defparam i1_2_lut_3_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i10664_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n24079));
    defparam i10664_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10665_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[4]), 
            .I3(\data_in_frame[1][4] ), .O(n24080));
    defparam i10665_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10666_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n24081));
    defparam i10666_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10667_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n24082));
    defparam i10667_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10668_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n24083));
    defparam i10668_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10669_3_lut_4_lut (.I0(n8_adj_3235), .I1(n43226), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n24084));
    defparam i10669_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10654_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n24069));
    defparam i10654_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(\data_in_frame[11] [5]), .I1(n22928), 
            .I2(n23385), .I3(GND_net), .O(n43770));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1379 (.I0(n43590), .I1(\data_out_frame[10] [3]), 
            .I2(n22142), .I3(n43325), .O(n43326));
    defparam i1_2_lut_3_lut_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1380 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[10] [2]), 
            .I2(n43891), .I3(n40167), .O(n22599));
    defparam i1_2_lut_3_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1381 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[10] [2]), 
            .I2(n43891), .I3(\data_out_frame[18] [6]), .O(n43450));
    defparam i1_2_lut_3_lut_4_lut_adj_1381.LUT_INIT = 16'h9669;
    SB_LUT4 i10655_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n24070));
    defparam i10655_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1382 (.I0(\data_in_frame[10] [4]), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[6] [0]), .I3(n43490), .O(n43727));   // verilog/coms.v(82[17:28])
    defparam i1_2_lut_4_lut_adj_1382.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1383 (.I0(\data_in_frame[13] [7]), .I1(n23183), 
            .I2(n10_adj_3211), .I3(\data_in_frame[9] [3]), .O(n43635));
    defparam i1_2_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1384 (.I0(n23126), .I1(\data_in_frame[9] [7]), 
            .I2(n43754), .I3(\data_in_frame[7] [6]), .O(n43391));
    defparam i1_2_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1385 (.I0(\data_in_frame[10] [0]), .I1(\data_in_frame[7] [4]), 
            .I2(\data_in_frame[7] [5]), .I3(GND_net), .O(n23126));
    defparam i1_2_lut_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1386 (.I0(\data_in_frame[9] [5]), .I1(n43299), 
            .I2(n43748), .I3(n43474), .O(n40198));
    defparam i1_2_lut_4_lut_adj_1386.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1387 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[7] [7]), 
            .I2(\data_in_frame[10] [2]), .I3(\data_in_frame[6] [0]), .O(n43301));
    defparam i1_2_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1388 (.I0(n8_adj_3117), .I1(n43867), .I2(\data_in_frame[8] [1]), 
            .I3(n43801), .O(n43802));
    defparam i1_2_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1389 (.I0(\data_in_frame[7] [5]), .I1(Kp_23__N_515), 
            .I2(n43882), .I3(\data_in_frame[9] [7]), .O(n43801));
    defparam i2_3_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1390 (.I0(\data_in_frame[13] [5]), .I1(n23202), 
            .I2(n40137), .I3(\data_in_frame[11] [4]), .O(n40234));
    defparam i1_2_lut_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_4_lut (.I0(n43490), .I1(Kp_23__N_865), .I2(n43441), 
            .I3(n23209), .O(n16_adj_3199));   // verilog/coms.v(82[17:28])
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_in_frame[12] [7]), .I1(n22827), .I2(\data_in_frame[16] [7]), 
            .I3(GND_net), .O(n16_adj_3146));
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i10656_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n24071));
    defparam i10656_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(\data_in_frame[10][6] ), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[8] [1]), .I3(\data_in_frame[14]_c [7]), .O(n43739));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i10657_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n24072));
    defparam i10657_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10658_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n24073));
    defparam i10658_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10659_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n24074));
    defparam i10659_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1392 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n22456), .I3(GND_net), .O(n22453));   // verilog/coms.v(211[5:21])
    defparam i1_2_lut_3_lut_adj_1392.LUT_INIT = 16'hfefe;
    SB_LUT4 i10660_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n24075));
    defparam i10660_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10661_3_lut_4_lut (.I0(n8_adj_3261), .I1(n43226), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n24076));
    defparam i10661_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1393 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(\FRAME_MATCHER.state [3]), .I2(n22456), .I3(\FRAME_MATCHER.state [0]), 
            .O(n22441));   // verilog/coms.v(156[5:29])
    defparam i1_2_lut_3_lut_4_lut_adj_1393.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_3_lut_4_lut_adj_1394 (.I0(n22721), .I1(n5_adj_3218), .I2(n23358), 
            .I3(\data_in_frame[4] [6]), .O(n6_adj_3115));
    defparam i1_3_lut_4_lut_adj_1394.LUT_INIT = 16'hd77d;
    SB_LUT4 i29696_3_lut_4_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n22334), .I3(\FRAME_MATCHER.state [0]), 
            .O(n28434));
    defparam i29696_3_lut_4_lut_4_lut_4_lut.LUT_INIT = 16'hf8ff;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1395 (.I0(\FRAME_MATCHER.state [2]), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n22334), .I3(\FRAME_MATCHER.state [0]), 
            .O(n22454));
    defparam i2_2_lut_3_lut_4_lut_adj_1395.LUT_INIT = 16'hfdff;
    SB_LUT4 equal_66_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3261));   // verilog/coms.v(149[7:23])
    defparam equal_66_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1396 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43226), .I3(\FRAME_MATCHER.i [0]), .O(n43229));   // verilog/coms.v(149[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1396.LUT_INIT = 16'hfdff;
    SB_LUT4 i14888_2_lut_2_lut_3_lut (.I0(n28434), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n28284));
    defparam i14888_2_lut_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1397 (.I0(\FRAME_MATCHER.state [0]), 
            .I1(\FRAME_MATCHER.state [1]), .I2(n22334), .I3(\FRAME_MATCHER.state [2]), 
            .O(n63_adj_3342));   // verilog/coms.v(248[5:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1397.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1398 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43235), .I3(\FRAME_MATCHER.i [0]), .O(n43236));   // verilog/coms.v(149[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1398.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_3_lut_4_lut_adj_1399 (.I0(n22126), .I1(\data_out_frame[17] [5]), 
            .I2(n1784), .I3(n39462), .O(n44835));
    defparam i2_3_lut_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1400 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n43247), .I3(\FRAME_MATCHER.i [0]), .O(n43251));   // verilog/coms.v(149[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1400.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_3_lut_4_lut_adj_1401 (.I0(\data_in_frame[9] [5]), .I1(n43299), 
            .I2(\data_in_frame[12] [1]), .I3(n22721), .O(n43754));
    defparam i2_3_lut_4_lut_adj_1401.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1402 (.I0(n23282), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[17] [1]), .I3(n44887), .O(n44979));
    defparam i2_3_lut_4_lut_adj_1402.LUT_INIT = 16'h6996;
    uart_tx tx (.n23776(n23776), .n23779(n23779), .n23778(n23778), .clk32MHz(clk32MHz), 
            .n23781(n23781), .n23784(n23784), .n23787(n23787), .n23790(n23790), 
            .n23793(n23793), .n23796(n23796), .n23799(n23799), .n23803(n23803), 
            .r_Bit_Index({r_Bit_Index}), .n23806(n23806), .\r_SM_Main[1] (r_SM_Main[1]), 
            .n23782(n23782), .tx_data({tx_data}), .n23785(n23785), .n23788(n23788), 
            .GND_net(GND_net), .n23602(n23602), .n23716(n23716), .n4037(n4037), 
            .n23845(n23845), .n23791(n23791), .n23794(n23794), .n23797(n23797), 
            .n23844(n23844), .VCC_net(VCC_net), .n23846(n23846), .n23849(n23849), 
            .n25425(n25425), .tx_active(tx_active), .tx_o(tx_o), .\r_SM_Main_2__N_2747[0] (r_SM_Main_2__N_2747[0]), 
            .n23530(n23530), .tx_enable(tx_enable)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(104[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n23809(n23809), .r_Bit_Index({r_Bit_Index_adj_9}), 
            .n23812(n23812), .n28794(n28794), .r_SM_Main({\r_SM_Main[2] , 
            \r_SM_Main[1] , Open_47}), .n24357(n24357), .rx_data({rx_data}), 
            .VCC_net(VCC_net), .rx_data_ready(rx_data_ready), .r_Rx_Data(r_Rx_Data), 
            .LED_c(LED_c), .GND_net(GND_net), .n23596(n23596), .n23714(n23714), 
            .n4015(n4015), .n23819(n23819), .n23818(n23818), .n23817(n23817), 
            .n23816(n23816), .n23853(n23853), .n23815(n23815), .n23814(n23814), 
            .n23813(n23813), .n23751(n23751), .n28760(n28760), .n1(n1), 
            .n28350(n28350), .n4(n4), .n4_adj_1(n4_adj_7), .n22470(n22470), 
            .n22462(n22462), .n4_adj_2(n4_adj_8), .n47207(n47207), .n47206(n47206)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(90[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n23776, n23779, n23778, clk32MHz, n23781, n23784, 
            n23787, n23790, n23793, n23796, n23799, n23803, r_Bit_Index, 
            n23806, \r_SM_Main[1] , n23782, tx_data, n23785, n23788, 
            GND_net, n23602, n23716, n4037, n23845, n23791, n23794, 
            n23797, n23844, VCC_net, n23846, n23849, n25425, tx_active, 
            tx_o, \r_SM_Main_2__N_2747[0] , n23530, tx_enable) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output n23776;
    output n23779;
    input n23778;
    input clk32MHz;
    input n23781;
    input n23784;
    input n23787;
    input n23790;
    input n23793;
    input n23796;
    input n23799;
    input n23803;
    output [2:0]r_Bit_Index;
    input n23806;
    output \r_SM_Main[1] ;
    output n23782;
    input [7:0]tx_data;
    output n23785;
    output n23788;
    input GND_net;
    output n23602;
    output n23716;
    output n4037;
    output n23845;
    output n23791;
    output n23794;
    output n23797;
    output n23844;
    input VCC_net;
    input n23846;
    input n23849;
    input n25425;
    output tx_active;
    output tx_o;
    input \r_SM_Main_2__N_2747[0] ;
    output n23530;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n36982, n36981, n43041, n36980, n20331;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n36979, n36978;
    wire [2:0]r_SM_Main_2__N_2744;
    
    wire n28703, n28574, n39058, n10, n45246, n9, n45244, n36977, 
        n36976, n36975, n45354, n45355, n50017, n45286, n45285, 
        o_Tx_Serial_N_2775, n44263, n23755, n10_adj_3109, n5, n12, 
        n19647;
    
    SB_LUT4 add_59_10_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[8]), 
            .I2(r_SM_Main[2]), .I3(n36982), .O(n23776)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_59_9_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[7]), 
            .I2(r_SM_Main[2]), .I3(n36981), .O(n23779)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hA3AC;
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n23778));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23781));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23784));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n23787));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23790));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23793));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n23796));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n23799));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23803));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23806));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(\r_SM_Main[1] ), .C(clk32MHz), .D(n43041));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_9 (.CI(n36981), .I0(r_Clock_Count[7]), .I1(r_SM_Main[2]), 
            .CO(n36982));
    SB_LUT4 add_59_8_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[6]), 
            .I2(r_SM_Main[2]), .I3(n36980), .O(n23782)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hA3AC;
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY add_59_8 (.CI(n36980), .I0(r_Clock_Count[6]), .I1(r_SM_Main[2]), 
            .CO(n36981));
    SB_LUT4 add_59_7_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[5]), 
            .I2(r_SM_Main[2]), .I3(n36979), .O(n23785)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_7 (.CI(n36979), .I0(r_Clock_Count[5]), .I1(r_SM_Main[2]), 
            .CO(n36980));
    SB_LUT4 add_59_6_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[4]), 
            .I2(r_SM_Main[2]), .I3(n36978), .O(n23788)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_6 (.CI(n36978), .I0(r_Clock_Count[4]), .I1(r_SM_Main[2]), 
            .CO(n36979));
    SB_LUT4 i15300_2_lut (.I0(r_SM_Main_2__N_2744[1]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n28703));
    defparam i15300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n28574));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n39058), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(r_SM_Main_2__N_2744[1]));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_2744[1]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main[1] ), .O(n23602));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i10301_3_lut (.I0(n23602), .I1(n28574), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n23716));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i10301_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1122_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4037));   // verilog/uart_tx.v(98[36:51])
    defparam i1122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n39058));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i29746_2_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[4]), 
            .I2(GND_net), .I3(GND_net), .O(n45246));
    defparam i29746_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_825 (.I0(r_Clock_Count[6]), .I1(\r_SM_Main[1] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n9));
    defparam i2_3_lut_adj_825.LUT_INIT = 16'h5454;
    SB_LUT4 i29744_3_lut (.I0(r_Clock_Count[7]), .I1(n39058), .I2(r_Clock_Count[5]), 
            .I3(GND_net), .O(n45244));
    defparam i29744_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n45244), .I2(n9), .I3(n45246), 
            .O(n23845));   // verilog/uart_tx.v(31[16:25])
    defparam i1_4_lut.LUT_INIT = 16'haaba;
    SB_LUT4 add_59_5_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[3]), 
            .I2(r_SM_Main[2]), .I3(n36977), .O(n23791)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_5 (.CI(n36977), .I0(r_Clock_Count[3]), .I1(r_SM_Main[2]), 
            .CO(n36978));
    SB_LUT4 add_59_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[2]), 
            .I2(r_SM_Main[2]), .I3(n36976), .O(n23794)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_4 (.CI(n36976), .I0(r_Clock_Count[2]), .I1(r_SM_Main[2]), 
            .CO(n36977));
    SB_LUT4 add_59_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[1]), 
            .I2(r_SM_Main[2]), .I3(n36975), .O(n23797)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_3 (.CI(n36975), .I0(r_Clock_Count[1]), .I1(r_SM_Main[2]), 
            .CO(n36976));
    SB_LUT4 add_59_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[0]), 
            .I2(r_SM_Main[2]), .I3(VCC_net), .O(n23844)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(r_SM_Main[2]), 
            .CO(n36975));
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n23846));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n20331), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n45354), 
            .I2(n45355), .I3(r_Bit_Index[2]), .O(n50017));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n23849));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 n50017_bdd_4_lut (.I0(n50017), .I1(n45286), .I2(n45285), .I3(r_Bit_Index[2]), 
            .O(o_Tx_Serial_N_2775));
    defparam n50017_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n44263));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n23755));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n25425));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n10_adj_3109));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2747[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n5));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i26_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_2775), .I2(\r_SM_Main[1] ), 
            .I3(GND_net), .O(n12));
    defparam i26_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i25_3_lut (.I0(n12), .I1(tx_o), .I2(r_SM_Main[2]), .I3(GND_net), 
            .O(n10_adj_3109));
    defparam i25_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i2_4_lut_adj_826 (.I0(n5), .I1(r_SM_Main[2]), .I2(\r_SM_Main[1] ), 
            .I3(n28703), .O(n23530));
    defparam i2_4_lut_adj_826.LUT_INIT = 16'h3202;
    SB_LUT4 i6341_4_lut (.I0(\r_SM_Main_2__N_2747[0] ), .I1(n28574), .I2(\r_SM_Main[1] ), 
            .I3(r_SM_Main_2__N_2744[1]), .O(n19647));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i6341_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i1_4_lut_adj_827 (.I0(r_SM_Main[2]), .I1(n19647), .I2(r_SM_Main_2__N_2744[1]), 
            .I3(r_SM_Main[0]), .O(n23755));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut_adj_827.LUT_INIT = 16'h0544;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29785_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45285));
    defparam i29785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29786_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45286));
    defparam i29786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29855_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45355));
    defparam i29855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29854_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45354));
    defparam i29854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main_2__N_2744[1]), .I1(r_SM_Main[0]), 
            .I2(\r_SM_Main[1] ), .I3(r_SM_Main[2]), .O(n44263));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i3_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_2747[0] ), 
            .I2(r_SM_Main[2]), .I3(\r_SM_Main[1] ), .O(n20331));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_2744[1]), 
            .I2(r_SM_Main[0]), .I3(\r_SM_Main[1] ), .O(n43041));   // verilog/uart_tx.v(31[16:25])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1540;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n23809, r_Bit_Index, n23812, n28794, r_SM_Main, 
            n24357, rx_data, VCC_net, rx_data_ready, r_Rx_Data, LED_c, 
            GND_net, n23596, n23714, n4015, n23819, n23818, n23817, 
            n23816, n23853, n23815, n23814, n23813, n23751, n28760, 
            n1, n28350, n4, n4_adj_1, n22470, n22462, n4_adj_2, 
            n47207, n47206) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n23809;
    output [2:0]r_Bit_Index;
    input n23812;
    input n28794;
    output [2:0]r_SM_Main;
    input n24357;
    output [7:0]rx_data;
    input VCC_net;
    output rx_data_ready;
    output r_Rx_Data;
    input LED_c;
    input GND_net;
    output n23596;
    output n23714;
    output n4015;
    input n23819;
    input n23818;
    input n23817;
    input n23816;
    input n23853;
    input n23815;
    input n23814;
    input n23813;
    input n23751;
    output n28760;
    output n1;
    output n28350;
    output n4;
    output n4_adj_1;
    output n22470;
    output n22462;
    output n4_adj_2;
    output n47207;
    output n47206;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[8:16])
    
    wire n23749;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n23760, n42679, n23766, n23769, n23772, n23775, n42673, 
        r_Rx_Data_R, n28551;
    wire [2:0]r_SM_Main_2__N_2673;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    
    wire n43189, n47082, n43901, n47088, n47085, n47083, n47246, 
        n47086, n4_c, n30515, n14, n47251, n10, n47248, n38;
    wire [2:0]r_SM_Main_2__N_2679;
    
    wire n44886, n47087, n36974, n108, n36973, n36972, n36971, 
        n36970, n36969, n36968, n47084, n23843, n23517, n22317;
    
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n23749));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n23760));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n42679));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n23766));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n23769));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n23772));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n23775));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n23809));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n23812));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n28794));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n24357));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n42673));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(LED_c));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n28551));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_2673[2]), .I2(r_SM_Main_c[0]), 
            .I3(r_SM_Main[1]), .O(n23596));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i10299_3_lut (.I0(n23596), .I1(n28551), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n23714));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i10299_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1100_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4015));   // verilog/uart_rx.v(102[36:51])
    defparam i1100_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_2673[2]), 
            .R(n43189));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i17179_3_lut (.I0(r_Clock_Count[1]), .I1(n47082), .I2(n43901), 
            .I3(GND_net), .O(n23775));
    defparam i17179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17209_3_lut (.I0(r_Clock_Count[2]), .I1(n47088), .I2(n43901), 
            .I3(GND_net), .O(n23772));
    defparam i17209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17195_3_lut (.I0(r_Clock_Count[3]), .I1(n47085), .I2(n43901), 
            .I3(GND_net), .O(n23769));
    defparam i17195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17185_3_lut (.I0(r_Clock_Count[4]), .I1(n47083), .I2(n43901), 
            .I3(GND_net), .O(n23766));
    defparam i17185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_3_lut (.I0(r_Clock_Count[5]), .I1(n47246), .I2(n43901), 
            .I3(GND_net), .O(n42679));
    defparam i11_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i17199_3_lut (.I0(r_Clock_Count[6]), .I1(n47086), .I2(n43901), 
            .I3(GND_net), .O(n23760));
    defparam i17199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15169_3_lut (.I0(r_Clock_Count[3]), .I1(n4_c), .I2(n30515), 
            .I3(GND_net), .O(r_SM_Main_2__N_2673[2]));
    defparam i15169_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i6_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[6]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i32423_4_lut (.I0(n47251), .I1(r_SM_Main_c[0]), .I2(n14), 
            .I3(n10), .O(n47248));
    defparam i32423_4_lut.LUT_INIT = 16'hb333;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n47248), .I2(r_SM_Main_2__N_2673[2]), 
            .I3(r_SM_Main[1]), .O(n38));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_4_lut_adj_821 (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_Clock_Count[4]), .O(n4_c));
    defparam i1_4_lut_adj_821.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_2__N_2679[0]), .I2(r_Rx_Data), 
            .I3(r_SM_Main_c[0]), .O(n44886));
    defparam i3_4_lut.LUT_INIT = 16'h1000;
    SB_LUT4 i28410_3_lut (.I0(r_SM_Main[2]), .I1(n38), .I2(n44886), .I3(GND_net), 
            .O(n43901));
    defparam i28410_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i17203_3_lut (.I0(r_Clock_Count[7]), .I1(n47087), .I2(n43901), 
            .I3(GND_net), .O(n23749));
    defparam i17203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_62_9_lut (.I0(n108), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n36974), .O(n47087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n108), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n36973), .O(n47086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_8 (.CI(n36973), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n36974));
    SB_LUT4 add_62_7_lut (.I0(n108), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n36972), .O(n47246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n36972), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n36973));
    SB_LUT4 add_62_6_lut (.I0(n108), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n36971), .O(n47083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n36971), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n36972));
    SB_LUT4 add_62_5_lut (.I0(n108), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n36970), .O(n47085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n36970), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n36971));
    SB_LUT4 add_62_4_lut (.I0(n108), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n36969), .O(n47088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_4 (.CI(n36969), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n36970));
    SB_LUT4 add_62_3_lut (.I0(n108), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n36968), .O(n47082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n36968), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n36969));
    SB_LUT4 add_62_2_lut (.I0(n108), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n47084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n36968));
    SB_LUT4 i2_3_lut_4_lut (.I0(n4_c), .I1(n30515), .I2(r_Rx_Data), .I3(r_Clock_Count[5]), 
            .O(n10));   // verilog/uart_rx.v(68[17:52])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h00bf;
    SB_LUT4 i1_2_lut_3_lut (.I0(n4_c), .I1(n30515), .I2(r_Clock_Count[3]), 
            .I3(GND_net), .O(r_SM_Main_2__N_2679[0]));   // verilog/uart_rx.v(68[17:52])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i32401_2_lut_3_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[7]), .I3(GND_net), .O(n47251));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i32401_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i1_2_lut_3_lut_adj_822 (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[1]), 
            .I2(r_Clock_Count[0]), .I3(GND_net), .O(n30515));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_adj_822.LUT_INIT = 16'h8080;
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n23843));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n23819));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n23818));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n23817));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n23816));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n23853));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n23815));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n23814));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n23813));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n23751));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i34447_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_c[0]), 
            .I3(GND_net), .O(n43189));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34447_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_2673[2]), 
            .I3(r_SM_Main_c[0]), .O(n23517));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n23517), 
            .I3(rx_data_ready), .O(n42673));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n28551), .I1(r_SM_Main_2__N_2673[2]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n28760));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_2679[0]), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i14950_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n28350));
    defparam i14950_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_72_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_72_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_74_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_74_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(n22317), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n22470));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i17191_3_lut (.I0(r_Clock_Count[0]), .I1(n47084), .I2(n43901), 
            .I3(GND_net), .O(n23843));
    defparam i17191_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_823 (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main_2__N_2673[2]), .O(n22317));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut_adj_823.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_824 (.I0(r_Bit_Index[0]), .I1(n22317), .I2(GND_net), 
            .I3(GND_net), .O(n22462));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_824.LUT_INIT = 16'heeee;
    SB_LUT4 equal_76_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_76_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32408_2_lut (.I0(r_SM_Main_2__N_2673[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n47207));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i32408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32171_3_lut (.I0(r_SM_Main_c[0]), .I1(r_SM_Main_2__N_2679[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n47206));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i32171_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i39_1_lut_4_lut (.I0(r_SM_Main[2]), .I1(n47248), .I2(r_SM_Main_2__N_2673[2]), 
            .I3(r_SM_Main[1]), .O(n108));
    defparam i39_1_lut_4_lut.LUT_INIT = 16'hafbb;
    
endmodule
