// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Feb 17 14:18:35 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, CS_CLK_c, CS_c, CS_MISO_c, 
        INLC_c_0, INHC_c_0, INLB_c_0, INHB_c_0, INLA_c_0, INHA_c_0;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3, pwm_out, dir, GHA, GHB, GHC;
    wire [23:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[20:32])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire h1, h2, h3;
    wire [7:0]commutation_state;   // verilog/TinyFPGA_B.v(116[12:29])
    wire [7:0]commutation_state_prev;   // verilog/TinyFPGA_B.v(117[12:34])
    
    wire dti;
    wire [7:0]dti_counter;   // verilog/TinyFPGA_B.v(126[12:23])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(223[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(225[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(226[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(227[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(228[22:24])
    
    wire n38196, n15;
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(229[22:24])
    
    wire n37970;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(231[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(232[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(233[22:35])
    
    wire n14, n37798, n37969;
    wire [12:0]current;   // verilog/TinyFPGA_B.v(235[22:29])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(263[22:33])
    wire [7:0]data;   // verilog/TinyFPGA_B.v(326[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(350[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(358[15:20])
    
    wire pwm_setpoint_23__N_215;
    wire [23:0]pwm_setpoint_23__N_191;
    
    wire n38195, n33, n32, n31, n30, n29, n28, n27, n26, n25, 
        n24, n23, n22, n21, n38194;
    wire [7:0]commutation_state_7__N_216;
    
    wire commutation_state_7__N_224, n28304, n28303;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(222[11:28])
    
    wire n28302, n28301, n28300, n28299, n28298, n28297, GHA_N_367, 
        GLA_N_384, GHB_N_389, GLB_N_398, GHC_N_403, GLC_N_412, dti_N_416, 
        n28296, n28295, n28294, n28293, n28292, n28291, RX_N_10, 
        n48513, n1632;
    wire [31:0]motor_state_23__N_123;
    wire [32:0]encoder0_position_scaled_23__N_51;
    
    wire encoder1_position_scaled_23__N_279;
    wire [31:0]encoder1_position_scaled_23__N_75;
    wire [23:0]displacement_23__N_99;
    
    wire n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
        n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
        n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, 
        n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
        n37968, n731, n1195, n37967, n38193, n38192, n37966, n28290, 
        n47541, n37797, n38191, n43094, n43084, n1673;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(224[11:28])
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n28289, n37965, n37796, n43068, n28288, n26390, n37795, 
        n37964;
    wire [3:0]state_3__N_528;
    
    wire n38190, n37963, n37794, n37962, n37961, n37960, n37793, 
        n18934, n38189, n37792, n37959, n33280, n37791, n38188, 
        n28287, n28286, n28285, n28284, n28283, n28282, n28281, 
        n28280, n28279, n6, n37958, n37957, n38187, n38186, n23805, 
        n28278, n38185, n38184, n44848, n20, n652, n37956, n37955, 
        n37790, n37954, n43722, n38183, n38182, n37953, n38181, 
        n28277, n19, n18, n37952, n37951, n28276, n28275, n28274, 
        n37950, n38180, n37949, n28273, n37789, n37948, n28272, 
        n37947, n38179, n37946, n43011, n38178, n28271, n28270, 
        n38177, n38176, n38175, n37945, n38174, n28269, n42999, 
        n42997, n42995, n42993, n37788, n37787, n38173, n38172, 
        n625, n42988;
    wire [2:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n17, n37944, n623, n3, n4, n5, n6_adj_5138, n7, n8, 
        n9, n10, n11, n12, n13, n14_adj_5139, n15_adj_5140, n16, 
        n17_adj_5141, n18_adj_5142, n19_adj_5143, n20_adj_5144, n21_adj_5145, 
        n22_adj_5146, n23_adj_5147, n24_adj_5148, n25_adj_5149, n622, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n38171, n38170, n38169, n38168, n38167;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire n621, tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n38166, n38165, n122, n10_adj_5150, n37943, n37942;
    wire [31:0]\FRAME_MATCHER.state_31__N_2660 ;
    
    wire n38164, n38163, n37941, n38162, n38161, n16_adj_5151, n38160, 
        n37438, n37940, n38159, n37786, n38158, n38157, n37785, 
        n41451, n38156, n37784, n37783, n37782, n48548, n37781, 
        n38155, n38154, n8_adj_5152, n47540, n4_adj_5153, n38153, 
        n38152, n37939, n37938, n34196, n38151, n37937, n37936, 
        n37935, n37934, n37933, n47612, n7_adj_5154, n38150, n37422, 
        n37932, n38149, n38148, n4_adj_5155, n37931, n38147, n38146, 
        n37930, n38145, n37780, n37779, n38144, n37929, n37928, 
        n38143, n37778, n37927, n38142, n43273, n38141, n38140, 
        n37777, n38139, n38138, n38137, n37776, n38136, n37926, 
        n37775, n38135, n38134, n38133, n38132, n38131, n37774, 
        n38130, n38129, n38128, n38127, n37773, n38126, n38125, 
        n37772, n43352, n38124, n48486, n37925, n38123, n38122, 
        n38121, n38120, n43363, n37924, n37923, n37527, n38119, 
        n33250, n37922, n37921, n37526, n37771, n37770, n37920, 
        n48064, n38118, n37919, n37769, n37918, n37917, n37768, 
        n37767, n38117, n37766, n38116, n37916, n37915, n38115, 
        n38114, n38113, n38112, n37914, n37913, n38111, n37912, 
        n37911, n38110, n37525, n37910, n38109, n38108, n38107, 
        n37909, n38106, n38105, n33185, n38104, n34134, n33903, 
        n38103, n38102, n37908, n38101, n38100, n37907, n38099, 
        n37524, n38098, n34130, n38097, n38096, n38095, n38094, 
        n37906, n38093, n38092, n38091, n38090, n38089, n38088, 
        n38087, n37905, n37904, n34122, n34010, n37903, n37902, 
        n37523, n37522, n34118, n37901, n37900, n37521, n37899, 
        n38086, n34114, n38085, n37749, n37748, n33881, n38084, 
        n34084, n34106, n34102, n37520, n34100, n34096, n34022, 
        n37898, n34094, n37747, n34092, n34090, n38083, n37897, 
        n38082, n33332, n37896, n34070, n33328, n37519, n37518, 
        n2, n37517, n48457, n37895, n38081, n37894, n38080, n37893, 
        n3303, n37746, n37745;
    wire [31:0]\FRAME_MATCHER.state_31__N_2788 ;
    
    wire n37744, n38079, n37743, n37742, n37892, n37891, n37741, 
        n37890, n37740, n38078, n37516, n37739, n37515, n38077, 
        n37514, n37437, n37738, n37889, n38076, n37888, n37737, 
        n37887, n37886, n37513, n38075, n37736, n37735, n34066, 
        n37885, n34064, n37512, n38074, n37884, n38073, n37734, 
        n37511, n37510, n37733, n37509, n38072, n37732, n4452, 
        n37883, n37882, n37881, n38071, n37880, n37879, n37508, 
        n38070, n34062, n37878, n37731, n38069, n38068, n37507, 
        n38067, n37877, n37506, n37505, n37876, n37504, n37730, 
        n37503, n37502, n7_adj_5156, n38066, n37729, n37875, n37874, 
        n38065, n37873, n37728, n37501, n37727, n37872, n37871, 
        n38064, n37500, n37436, n38063, n37870, n38062, n37869, 
        n37435, n37868, n38061, n37867, n38060, n37421, n37420, 
        n38059, n37866, n5_adj_5157, n44019, n60, n62, n43381, 
        n45760, n48428, n42989, n15_adj_5158, n6_adj_5159, n25_adj_5160, 
        n24_adj_5161, n47600, n43289, n48395, n405, n44592, n23_adj_5162, 
        n22_adj_5163, n21_adj_5164, n20_adj_5165, n19_adj_5166, n18_adj_5167, 
        n17_adj_5168, n16_adj_5169, n15_adj_5170, n14_adj_5171, n13_adj_5172, 
        n12_adj_5173, n11_adj_5174, n10_adj_5175, n9_adj_5176, n8_adj_5177, 
        n7_adj_5178, n6_adj_5179, n5_adj_5180, n4_adj_5181, n3_adj_5182, 
        n48874, n8_adj_5183, n4_adj_5184, n44235, n48364, n5615, 
        n45757, n14_adj_5185, n48873, n38058, n47917, n37865, n34024, 
        n38057, n28783, n28782, n28781, n28780, n26277, n5_adj_5186, 
        n28779, n28778, n28777, n28776, n28775, n28774, n28773;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n28772, n28771, n28770, n15_adj_5187, n14_adj_5188, 
        n13_adj_5189, direction_N_3907, n10_adj_5190, n28746, n28745, 
        n28744, n28743, n28742, n28741, n28740, n28739, n48333, 
        n15_adj_5191, n28730, n28729, n28728, n4_adj_5192, n28727, 
        n28726, n28725, n28724, n28723, n28714, n28713;
    wire [1:0]a_new_adj_5325;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_5194, n1964, n28712, n28711, n28710, n28709, 
        n37864, n37434, n28708, n28707, direction_N_3907_adj_5195, 
        n28692, n28691, n28690, n28689, n28688, n5_adj_5196, n28687, 
        n28686, n28685, n11_adj_5197, n28684, n28683, n28682, n28681, 
        n9_adj_5198, n46900, n28669, n28668, n28667, n26409, n28666, 
        n28665, n37433, n28664, n28663, n28662, n4_adj_5199, n28652, 
        n28651, n28650, n28649, n4_adj_5200, rw;
    wire [7:0]state_adj_5349;   // verilog/eeprom.v(23[11:16])
    
    wire n28648, n28647, n28646, n28645, n28644, n28643, n28642, 
        n28641, n28640, n28639, n12_adj_5202, n11_adj_5203, n28638, 
        n28637, n28636, n28635, n10_adj_5204, n9_adj_5205, n28634, 
        n28633, n28632, n28631;
    wire [15:0]data_adj_5353;   // verilog/tli4970.v(27[14:18])
    
    wire n28630, n28629, n28628, n8_adj_5214, n7_adj_5215, n28268, 
        n28267, n28266, n28265, n28264, n28263, n28262, n28261, 
        n28260, n28259, n28258, n28257, n28256, n28255, n28254, 
        n28253, n28627, n28626, n28625, n27874, n46890, n28624, 
        n28623, n28622, n28621, n28620, n28619, n28618, n28617, 
        n28616, n28615, n28614, n28613, n28612, n28611, n28610, 
        n28609, n28608, n28607, n28606, n28605, n4_adj_5216, n28604, 
        n28603, n6_adj_5217, n28602, n28601, n28600, state_7__N_4293, 
        n7072, n28599, n28598, n28252, n28251, n28597, n28596, 
        n28595, n28594, n28593, n28592, n28591, n28590, n28589, 
        n28588, n28587, n28586, n28585, n28584, n45546, n4_adj_5218, 
        n28583, n38056, n28582, n28581, n28580, n27844, n28084, 
        n28579, n28578, n27840, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n28577, n28576, n28575, n28574, n28573, n28572, n28571, 
        n45538, n48038, n34018, n40583;
    wire [2:0]r_SM_Main_2__N_3542;
    
    wire n45534, n28250;
    wire [2:0]r_SM_Main_adj_5364;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5366;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main_2__N_3616;
    wire [2:0]r_SM_Main_2__N_3613;
    
    wire n43278, n28125, n48300, n28546, n28545, n28544, n28543, 
        n28542, n28541, n28540, n28539, n28249, n28123, n28248, 
        n28530, n28529, n28528, n28527, n28526, n28525, n45526, 
        n43298;
    wire [7:0]state_adj_5377;   // verilog/i2c_controller.v(33[12:17])
    
    wire n28524;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n28523, n28522, n28521, n28520, enable_slow_N_4190, n45520, 
        n7233, n42299, n28519;
    wire [7:0]state_7__N_4087;
    
    wire n28518, n28517, n28516, n28515, n28514, n28247, n6692, 
        n28510, n28509, n28508, n46883, n38055, n37863, n28507, 
        n28506, n28505;
    wire [7:0]state_7__N_4103;
    
    wire n45514, n38054, n28501, n28500, n28499, n28498, n28497, 
        n28496, n28495, n28494, n45510, n28493, n28492, n28491, 
        n27791, n28246, n28245, n28244, n28243, n28242, n28241, 
        n28240, n28239, n5_adj_5224, n7270, n28238, n28490, n28237, 
        n28236, n28489, n4_adj_5225, n3_adj_5226, n2_adj_5227, n45498, 
        n45494, n28488, n28235, n28234, n28233, n28232, n28229, 
        n28227, n28226, n28225, n28224, n28223, n28222, n28221, 
        n28219, n28218, n28217, n28215, n28214, n28213, n28212, 
        n28211, n28210, n28209, n28208, n28207, n28206, n28205, 
        n28204, n28203, n28202, n28487, n28201, n28200, n28486, 
        n28199, n28198, n28483, n38053, n45490, n28482, n28480, 
        n28479, n28478, n28197, n28196, n28195, n28477, n28476, 
        n44847, n28475, n28474, n45484, n28473, n828, n829, n830, 
        n831, n832, n833, n834, n861, n46878, n896, n897, n898, 
        n899, n900, n901, n45482, n927, n928, n929, n930, n931, 
        n932, n933, n934, n935, n936, n937, n938, n939, n940, 
        n941, n942, n943, n944, n945, n946, n947, n948, n949, 
        n950, n951, n952, n953, n954, n955, n956, n957, n960, 
        n43335, n995, n996, n997, n998, n999, n1000, n1001, 
        n45476, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
        n1033, n6_adj_5228, n1059, n1093_adj_5229, n1094_adj_5230, 
        n1095_adj_5231, n1096_adj_5232, n1097_adj_5233, n1098_adj_5234, 
        n1099_adj_5235, n1100_adj_5236, n1101_adj_5237, n1125, n1126, 
        n1127, n1128, n1129, n1130, n1131, n1132, n1133, n42087, 
        n45468, n1158, n1193, n1194, n1195_adj_5238, n1196, n1197, 
        n1198, n1199, n1200, n1201, n45462, n1224, n1225, n1226, 
        n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1257, 
        n28472, n28156, n45456, n37862, n1292, n1293, n1294, n1295, 
        n1296, n1297, n1298, n1299, n1300, n1301, n37861, n34058, 
        n45452, n37860, n1323, n1324, n1325, n1326, n1327, n1328, 
        n1329, n1330, n1331, n1332, n1333, n45450, n1356, n38052, 
        n28471, n38051, n38050, n1391, n1392, n1393, n1394, n1395, 
        n1396, n1397, n1398, n1399, n1400, n1401, n1422, n1423, 
        n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
        n1432, n1433, n45436, n1455, n45430, n1490, n1491, n1492, 
        n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, 
        n1501, n45424, n1521, n1522, n1523, n1524, n1525, n1526, 
        n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1554, 
        n48262, n45422, n1589, n1590, n1591, n1592, n1593, n1594, 
        n1595, n1596, n1597, n1598, n1599, n1600, n1601, n45416, 
        n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
        n1628, n1629, n1630, n1631, n1632_adj_5239, n1633, n1653, 
        n23516, n45414, n45412, n1688, n1689, n1690, n1691, n1692, 
        n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
        n1701, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
        n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, 
        n43320, n1752, n45796, n1787, n1788, n1789, n1790, n1791, 
        n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
        n1800, n1801, n1818, n1819, n1820, n1821, n1822, n1823, 
        n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, 
        n1832, n1833, n45392, n1851, n45386, n44824, n45384, n45382, 
        n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, 
        n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, 
        n45376, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
        n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, 
        n1932, n1933, n23622, n45374, n1950, n1985, n1986, n1987, 
        n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
        n1996, n1997, n1998, n1999, n2000, n2001, n2016, n2017, 
        n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, 
        n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, 
        n2049, n45360, n2084, n2085, n2086, n2087, n2088, n2089, 
        n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
        n2098, n2099, n2100, n2101, n2115, n2116, n2117, n2118, 
        n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, 
        n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2148, 
        n28469, n27716, n2183, n2184, n2185, n2186, n2187, n2188, 
        n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, 
        n2197, n2198, n2199, n2200, n2201, n5_adj_5240, n2214, 
        n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
        n2231, n2232, n2233, n45354, n26445, n45350, n26440, n2247, 
        n45344, n2282, n2283, n2284, n2285, n2286, n2287, n2288, 
        n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, 
        n2297, n2298, n2299, n2300, n2301, n8_adj_5241, n45342, 
        n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
        n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, 
        n2329, n2330, n2331, n2332, n2333, n2346, n28468, n42267, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n45330, n38049, n37859, n2445, n42266, 
        n41875, n38048, n2480, n2481, n2482, n2483, n2484, n2485, 
        n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, 
        n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, 
        n42277, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
        n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, 
        n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, 
        n42264, n2544, n45324, n12_adj_5242, n43114, n45318, n2579, 
        n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, 
        n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, 
        n2596, n2597, n2598, n2599, n2600, n2601, n41869, n2610, 
        n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, 
        n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, 
        n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2643, 
        n42289, n45312, n26429, n2678, n2679, n2680, n2681, n2682, 
        n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, 
        n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, 
        n2699, n2700, n2701, n2709, n2710, n2711, n2712, n2713, 
        n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, 
        n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
        n2730, n2731, n2732, n2733, n45308, n2742, n42288, n42255, 
        n42287, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
        n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, 
        n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
        n2800, n2801, n2808, n2809, n2810, n2811, n2812, n2813, 
        n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, 
        n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
        n2830, n2831, n2832, n2833, n2841, n42285, n2876, n2877, 
        n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
        n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
        n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, 
        n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, 
        n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, 
        n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
        n2931, n2932, n2933, n45294, n2940, n28467, n2975, n2976, 
        n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, 
        n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, 
        n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
        n3001, n3006, n3007, n3008, n3009, n3010, n3011, n3012, 
        n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
        n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, 
        n3029, n3030, n3031, n3032, n3033, n3039, n45288, n3073, 
        n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
        n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
        n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
        n3098, n3099, n3100, n3101, n3105, n3106, n3107, n3108, 
        n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, 
        n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, 
        n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, 
        n3133, n3138, n26435, n41973, n3173, n3174, n3175, n3176, 
        n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, 
        n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, 
        n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, 
        n3201, n3204, n3205, n3206, n3207, n3208, n3209, n3210, 
        n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, 
        n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
        n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3237, 
        n48205, n26494, n3271, n3272, n3273, n3274, n3275, n3276, 
        n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, 
        n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
        n3293, n3294, n3295, n3296, n3298, n3299, n3300, n3301, 
        n43421, n28466, n45282, n34054, n28465, n28193, n45278, 
        n24_adj_5243, n28464, n41203, n44392, n28463, n28462, n62_adj_5244, 
        n7651, n28461, n27647, n27644, n45272, n27973, n26299, 
        n28458, n26302, n28457, n44389, n28456, n28455, n28454, 
        n27620, n7650, n28453, n27617, n45746, n45262, n45256, 
        n28192, n46841, n46840, n37468, n45252, n7648, n45242, 
        n37858, n38047, n45236, n45230, n7647, n7646, n14_adj_5245, 
        n10_adj_5246, n48191, n46839, n45220, n46838, n46837, n45214, 
        n38046, n4_adj_5247, n46836, n37857, n46835, n26286, n48177, 
        n38045, n45787, n45202, n38044, n48014, n28191, n41665, 
        n45198, n28190, n37856, n28189, n32652, n48162, n28188, 
        n37855, n38043, n45743, n38042, n45186, n45781, n45178, 
        n26432, n45172, n45162, n38041, n38040, n38039, n45156, 
        n37854, n38038, n37853, n38037, n38036, n37852, n37851, 
        n38035, n37850, n38034, n38033, n45150, n48147, n45148, 
        n28187, n45142, n37849, n45734, n26398, n45138, n45136, 
        n37848, n37467, n37847, n37846, n38032, n37466, n7_adj_5248, 
        n45124, n28185, n28184, n28183, n28182, n28181, n28180, 
        n45122, n28179, n43356, n42276, n45116, n48, n49, n50, 
        n51, n52, n53, n54, n55, n48130, n45110, n19799, n12_adj_5249, 
        n45106, n38031, n28178, n45773, n45100, n38456, n38455, 
        n45092, n38030, n48112, n38454, n45086, n28452, n28451, 
        n28450, n28449, n28448, n28447, n28446, n28445, n28444, 
        n28443, n28442, n28441, n28440, n28439, n28438, n28437, 
        n28433, n28432, n28431, n37845, n38453, n45082, n28428, 
        n28427, n28426, n28425, n28424, n28423, n28422, n28421, 
        n28420, n28419, n28177, n38452, n38029, n38028, n28176, 
        n28175, n28174, n28418, n28417, n28416, n28415, n28414, 
        n28413, n28412, n28411, n42166, n45076, n45074, n45062, 
        n47426, n7_adj_5250, n38451, n38450, n38449, n38448, n45056, 
        n28410, n28409, n28408, n28407, n28406, n28405, n28404, 
        n28403, n28402, n28401, n28400, n28399, n28398, n28397, 
        n28396, n28395, n28394, n28393, n28392, n28391, n28390, 
        n28389, n28387, n28384, n28383, n28382, n28381, n28380, 
        n28379, n45050, n45044, n45038, n45036, n10_adj_5251, n38447, 
        n38446, n45034, n28378, n28377, n28376, n28375, n28374, 
        n28373, n28372, n28371, n28370, n28369, n28368, n28367, 
        n28366, n28365, n47428, n38445, n42984, n28364, n28363, 
        n28362, n28361, n28360, n37844, n37843, n37432, n38444, 
        n37842, n38443, n38442, n38027, n38026, n28173, n28169, 
        n28168, n28167, n28166, n28359, n28358, n28357, n28356, 
        n28355, n28354, n28353, n28352, n38441, n38440, n37465, 
        n34048, n38025, n38439, n28165, n28164, n28163, n28162, 
        n28161, n28160, n28159, n28158, n28157, n28351, n28350, 
        n28349, n28348, n28347, n28346, n28345, n28344, n28343, 
        n38438, n26424, n34046, n38437, n45016, n37841, n38024, 
        n45010, n38436, n37431, n45008, n38435, n37464, n47434, 
        n37840, n38023, n28342, n28341, n28340, n41883, n28335, 
        n28331, n28330, n28329, n28328, n28327, n28326, n28325, 
        n28324, n28323, n28322, n28321, n28320, n28319, n28317, 
        n28316, n28315, n28314, n28313, n28312, n28311, n37463, 
        n37839, n38434, n28310, n28309, n28308, n28307, n28306, 
        n28305, n34042, n38433, n45002, n45000, n37462, n37461, 
        n37419, n38022, n20_adj_5252, n19_adj_5253, n38021, n17_adj_5254, 
        n38432, n38431, n38430, n38429, n38428, n38427, n38426, 
        n37838, n37837, n44990, n37430, n37836, n26482, n44984, 
        n42244, n37429, n34036, n44978, n38020, n37835, n37834, 
        n37833, n37832, n2_adj_5255, n3_adj_5256, n4_adj_5257, n5_adj_5258, 
        n6_adj_5259, n7_adj_5260, n8_adj_5261, n9_adj_5262, n10_adj_5263, 
        n11_adj_5264, n12_adj_5265, n13_adj_5266, n14_adj_5267, n15_adj_5268, 
        n16_adj_5269, n17_adj_5270, n18_adj_5271, n19_adj_5272, n20_adj_5273, 
        n21_adj_5274, n22_adj_5275, n23_adj_5276, n24_adj_5277, n25_adj_5278, 
        n26_adj_5279, n27_adj_5280, n28_adj_5281, n29_adj_5282, n30_adj_5283, 
        n31_adj_5284, n32_adj_5285, n33_adj_5286, n38019, n38018, 
        n44968, n38017, n44233, n38016, n37831, n44962, n37830, 
        n37829, n37460, n37828, n38015, n44956, n38014, n38013, 
        n37827, n38012, n38011, n44732, n37459, n38010, n44952, 
        n37458, n37826, n26285, n38009, n37457, n37825, n37824, 
        n44946, n37823, n37418, n44944, n38008, n37822, n44942, 
        n38007, n38006, n37821, n38005, n48229, n44926, n37456, 
        n37820, n37455, n38004, n44920, n38003, n38002, n47871, 
        n26296, n38001, n38000, n37999, n44914, n37998, n44908, 
        n47436, n44906, n37454, n37819, n37997, n37996, n37995, 
        n37818, n37994, n48088, n44896, n44894, n44892, n44890, 
        n44888, n37993, n37992, n37991, n37990, n37817, n37989, 
        n37988, n37987, n37986, n37816, n37428, n37815, n37985, 
        n44886, n44884, n37814, n37453, n37984, n37983, n37813, 
        n37812, n37982, n37811, n37452, n37451, n37810, n44882, 
        n37809, n37427, n44880, n44878, n37450, n37808, n44876, 
        n37807, n37981, n37449, n44874, n37980, n44872, n44870, 
        n37448, n37979, n44724, n44860, n37978, n38246, n38245, 
        n37806, n37417, n38244, n37805, n37447, n38243, n37977, 
        n38242, n37446, n38241, n38240, n38239, n38238, n38237, 
        n37426, n38236, n38235, n37425, n38234, n38233, n38232, 
        n44858, n37445, n37804, n38231, n38230, n37976, n38229, 
        n38228, n38227, n37803, n37416, n37444, n37443, n37802, 
        n38226, n44856, n37442, n38225, n38224, n44854, n37975, 
        n37441, n38223, n42251, n38222, n38221, n37440, n38220, 
        n38219, n38218, n38217, n38216, n38215, n38214, n37974, 
        n38213, n43270, n38212, n38211, n38210, n37415, n44852, 
        n38209, n37973, n44850, n38208, n38207, n7_adj_5287, n38206, 
        n37801, n37972, n38205, n13_adj_5288, n37424, n15_adj_5289, 
        n17_adj_5290, n38204, n21_adj_5291, n38203, n25_adj_5292, 
        n38202, n38201, n33292, n37, n39, n38200, n37800, n37439, 
        n37971, n38199, n38198, n37423, n7649, n38197, n43746, 
        n37799;
    
    VCC i2 (.Y(VCC_net));
    SB_LUT4 i14759_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n44019), 
            .I3(GND_net), .O(n28273));   // verilog/coms.v(127[12] 300[6])
    defparam i14759_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i14760_3_lut (.I0(\data_out_frame[22] [7]), .I1(current[7]), 
            .I2(n23622), .I3(GND_net), .O(n28274));   // verilog/coms.v(127[12] 300[6])
    defparam i14760_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5281), .I3(n38430), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_5148));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5172));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut (.I0(n2617), .I1(n45384), .I2(n2616), .I3(n45534), 
            .O(n45386));
    defparam i1_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n38430), 
            .I0(GND_net), .I1(n28_adj_5281), .CO(n38431));
    SB_DFFE dti_177 (.Q(dti), .C(CLK_c), .E(n27620), .D(dti_N_416));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i1_4_lut_adj_1571 (.I0(n2613), .I1(n2614), .I2(n45386), .I3(n2615), 
            .O(n45392));
    defparam i1_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5271));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33329_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n45392), 
            .O(n2643));
    defparam i33329_4_lut.LUT_INIT = 16'h0001;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_prev_i0 (.Q(commutation_state_prev[0]), .C(CLK_c), 
           .D(commutation_state[0]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_99[0]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4103[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5282), .I3(n38429), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n38440), 
            .I0(GND_net), .I1(n18_adj_5271), .CO(n38441));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n38429), 
            .I0(GND_net), .I1(n29_adj_5282), .CO(n38430));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5283), .I3(n38428), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5271), .I3(n38440), .O(n18)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .GND_net(GND_net), .CLK_c(CLK_c), .\state[1] (state[1]), .n41203(n41203), 
            .VCC_net(VCC_net), .timer({timer}), .neopxl_color({neopxl_color}), 
            .n43011(n43011), .\state_3__N_528[1] (state_3__N_528[1]), .n27791(n27791), 
            .n28195(n28195), .n28165(n28165), .LED_c(LED_c), .n28649(n28649), 
            .n28648(n28648), .n28647(n28647), .n28646(n28646), .n28645(n28645), 
            .n28644(n28644), .n28643(n28643), .n28642(n28642), .n28641(n28641), 
            .n28640(n28640), .n28639(n28639), .n28638(n28638), .n28637(n28637), 
            .n28636(n28636), .n28635(n28635), .n28634(n28634), .n28633(n28633), 
            .n28632(n28632), .n28631(n28631), .n28630(n28630), .n28629(n28629), 
            .n28628(n28628), .n28627(n28627), .n28626(n28626), .n28625(n28625), 
            .n28624(n28624), .n28623(n28623), .n28622(n28622), .n28621(n28621), 
            .n28620(n28620), .n28619(n28619), .NEOPXL_c(NEOPXL_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_CARRY add_224_8 (.CI(n37451), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n37452));
    SB_LUT4 unary_minus_10_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5147));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n7072), 
            .D(n1085), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2625_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n37526), 
            .O(n7647)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_5146));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2625_6 (.CI(n37526), .I0(n622), .I1(GND_net), .CO(n37527));
    SB_LUT4 unary_minus_10_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5145));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2625_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n37525), 
            .O(n7648)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n38428), 
            .I0(GND_net), .I1(n30_adj_5283), .CO(n38429));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5284), .I3(n38427), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32294_3_lut (.I0(n2445), .I1(n2346), .I2(n47428), .I3(GND_net), 
            .O(n47426));
    defparam i32294_3_lut.LUT_INIT = 16'h7f7f;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n38427), 
            .I0(GND_net), .I1(n31_adj_5284), .CO(n38428));
    SB_LUT4 i32302_3_lut (.I0(n2346), .I1(n2247), .I2(n2148), .I3(GND_net), 
            .O(n47434));
    defparam i32302_3_lut.LUT_INIT = 16'h7f7f;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n38441), 
            .I0(GND_net), .I1(n17_adj_5270), .CO(n38442));
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n37785), .O(n1094_adj_5230)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14761_3_lut (.I0(\data_out_frame[22] [6]), .I1(current[6]), 
            .I2(n23622), .I3(GND_net), .O(n28275));   // verilog/coms.v(127[12] 300[6])
    defparam i14761_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n37785), .I0(n1027), 
            .I1(VCC_net), .CO(n37786));
    SB_LUT4 mux_238_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[11]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5285), .I3(n38426), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32739_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n47871));
    defparam i32739_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14762_3_lut (.I0(\data_out_frame[22] [5]), .I1(current[5]), 
            .I2(n23622), .I3(GND_net), .O(n28276));   // verilog/coms.v(127[12] 300[6])
    defparam i14762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14644_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n27617), .I3(GND_net), .O(n28158));   // verilog/coms.v(127[12] 300[6])
    defparam i14644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1449_rep_33_3_lut (.I0(n2193), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n45746));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1449_rep_33_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1516_rep_31_3_lut (.I0(n45746), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n45743));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1516_rep_31_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32480_3_lut (.I0(n45743), .I1(n2126), .I2(n47434), .I3(GND_net), 
            .O(n47612));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32480_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32481_3_lut (.I0(n47612), .I1(n2490), .I2(n2445), .I3(GND_net), 
            .O(n2522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32481_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5141));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1649_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1649_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14763_3_lut (.I0(\data_out_frame[22] [4]), .I1(current[4]), 
            .I2(n23622), .I3(GND_net), .O(n28277));   // verilog/coms.v(127[12] 300[6])
    defparam i14763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32408_3_lut (.I0(n2028), .I1(n2392), .I2(n2346), .I3(GND_net), 
            .O(n47540));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32409_3_lut (.I0(n47540), .I1(n2491), .I2(n2445), .I3(GND_net), 
            .O(n47541));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14764_3_lut (.I0(\data_out_frame[22] [3]), .I1(current[3]), 
            .I2(n23622), .I3(GND_net), .O(n28278));   // verilog/coms.v(127[12] 300[6])
    defparam i14764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14645_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n27617), .I3(GND_net), .O(n28159));   // verilog/coms.v(127[12] 300[6])
    defparam i14645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14765_3_lut (.I0(\data_out_frame[22] [2]), .I1(current[2]), 
            .I2(n23622), .I3(GND_net), .O(n28279));   // verilog/coms.v(127[12] 300[6])
    defparam i14765_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14766_3_lut (.I0(\data_out_frame[22] [1]), .I1(current[1]), 
            .I2(n23622), .I3(GND_net), .O(n28280));   // verilog/coms.v(127[12] 300[6])
    defparam i14766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1651_3_lut (.I0(n47541), .I1(n45757), 
            .I2(n47426), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5173));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32370_3_lut (.I0(n2327), .I1(n2394), .I2(n2346), .I3(GND_net), 
            .O(n2426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32370_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14767_3_lut (.I0(\data_out_frame[22] [0]), .I1(current[0]), 
            .I2(n23622), .I3(GND_net), .O(n28281));   // verilog/coms.v(127[12] 300[6])
    defparam i14767_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14768_3_lut (.I0(\data_out_frame[21] [4]), .I1(current[12]), 
            .I2(n23622), .I3(GND_net), .O(n28282));   // verilog/coms.v(127[12] 300[6])
    defparam i14768_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32371_3_lut (.I0(n2426), .I1(n2493), .I2(n2445), .I3(GND_net), 
            .O(n2525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32371_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32372_3_lut (.I0(n2328), .I1(n2395), .I2(n2346), .I3(GND_net), 
            .O(n2427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14769_3_lut (.I0(\data_out_frame[21] [3]), .I1(current[11]), 
            .I2(n23622), .I3(GND_net), .O(n28283));   // verilog/coms.v(127[12] 300[6])
    defparam i14769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32373_3_lut (.I0(n2427), .I1(n2494), .I2(n2445), .I3(GND_net), 
            .O(n2526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14770_3_lut (.I0(\data_out_frame[21] [2]), .I1(current[10]), 
            .I2(n23622), .I3(GND_net), .O(n28284));   // verilog/coms.v(127[12] 300[6])
    defparam i14770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32139_3_lut (.I0(n2425), .I1(n2492), .I2(n2445), .I3(GND_net), 
            .O(n2524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32139_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[12]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33263_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48395));
    defparam i33263_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_5140));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[13]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_238_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[14]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n38426), 
            .I0(GND_net), .I1(n32_adj_5285), .CO(n38427));
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5286), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i33232_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48364));
    defparam i33232_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25), .I2(encoder0_position[31]), .I3(GND_net), .O(n950));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5286), .CO(n38426));
    SB_LUT4 i33354_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48486));
    defparam i33354_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_238_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[15]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_10_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_5139));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1572 (.I0(n2527), .I1(n2524), .I2(n2526), .I3(n2525), 
            .O(n44906));
    defparam i1_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1573 (.I0(n2523), .I1(n2521), .I2(n2528), .I3(n2522), 
            .O(n44908));
    defparam i1_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i14771_3_lut (.I0(\data_out_frame[21] [1]), .I1(current[9]), 
            .I2(n23622), .I3(GND_net), .O(n28285));   // verilog/coms.v(127[12] 300[6])
    defparam i14771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[16]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5174));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20526_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n34036));
    defparam i20526_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1574 (.I0(n2519), .I1(n2520), .I2(n44908), .I3(n44906), 
            .O(n44914));
    defparam i1_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1575 (.I0(n2529), .I1(n34036), .I2(n2530), .I3(n2531), 
            .O(n43352));
    defparam i1_4_lut_adj_1575.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1576 (.I0(n2517), .I1(n43352), .I2(n2518), .I3(n44914), 
            .O(n44920));
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1577 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n44920), 
            .O(n44926));
    defparam i1_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i33357_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n44926), 
            .O(n2544));
    defparam i33357_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_238_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[17]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i32758_2_lut (.I0(n23805), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(dti_N_416));
    defparam i32758_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_5217), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33416_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48548));
    defparam i33416_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5265));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5266));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14772_3_lut (.I0(\data_out_frame[21] [0]), .I1(current[8]), 
            .I2(n23622), .I3(GND_net), .O(n28286));   // verilog/coms.v(127[12] 300[6])
    defparam i14772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14773_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n23622), .I3(GND_net), .O(n28287));   // verilog/coms.v(127[12] 300[6])
    defparam i14773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14782_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n23622), .I3(GND_net), .O(n28296));   // verilog/coms.v(127[12] 300[6])
    defparam i14782_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1518_rep_22_3_lut (.I0(n2294), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n45734));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1518_rep_22_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14783_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n23622), .I3(GND_net), .O(n28297));   // verilog/coms.v(127[12] 300[6])
    defparam i14783_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5175));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5176));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32557_3_lut (.I0(n2224), .I1(n2291), .I2(n2247), .I3(GND_net), 
            .O(n2323));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32557_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32475_3_lut (.I0(n2323), .I1(n2390), .I2(n2346), .I3(GND_net), 
            .O(n2422));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32475_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5177));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1593_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1593_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5178));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24), .I2(encoder0_position[31]), .I3(GND_net), .O(n949));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5179));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5180));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32533_3_lut (.I0(n2225), .I1(n2292), .I2(n2247), .I3(GND_net), 
            .O(n2324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32533_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32477_3_lut (.I0(n2324), .I1(n2391), .I2(n2346), .I3(GND_net), 
            .O(n2423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32477_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32478_3_lut (.I0(n45757), .I1(n2028), .I2(n47428), .I3(GND_net), 
            .O(n2325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32478_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32479_3_lut (.I0(n2325), .I1(n2392), .I2(n2346), .I3(GND_net), 
            .O(n2424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32479_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n7072), 
            .D(n1084), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n7072), 
            .D(n1083), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n7072), 
            .D(n1082), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n7072), 
            .D(n1081), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n7072), 
            .D(n1080), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n7072), 
            .D(n1079), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n7072), 
            .D(n1078), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i33381_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48513));
    defparam i33381_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n7072), 
            .D(n1077), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i12_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n7270), .I2(n27874), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n41451));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i12_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_5204), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n935));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(n2426), .I1(n2428), .I2(n2424), .I3(n2423), 
            .O(n45342));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(n2427), .I1(n45342), .I2(n2422), .I3(n2425), 
            .O(n45344));
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(244[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5_adj_5224), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n405));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5267));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5270), .I3(n38441), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20589_4_lut (.I0(n949), .I1(n2431), .I2(n2432), .I3(n2433), 
            .O(n34100));
    defparam i20589_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1580 (.I0(n2419), .I1(n2420), .I2(n45344), .I3(n2421), 
            .O(n45350));
    defparam i1_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(n2429), .I1(n2430), .I2(GND_net), .I3(GND_net), 
            .O(n45538));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(n2418), .I1(n45538), .I2(n45350), .I3(n34100), 
            .O(n45354));
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'hfefa;
    SB_LUT4 i14774_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n23622), .I3(GND_net), .O(n28288));   // verilog/coms.v(127[12] 300[6])
    defparam i14774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[18]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_scaled_23__I_4_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_279));   // verilog/TinyFPGA_B.v(321[33:52])
    defparam encoder1_position_scaled_23__I_4_4_lut.LUT_INIT = 16'hccc8;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n38442), 
            .I0(GND_net), .I1(n16_adj_5269), .CO(n38443));
    SB_LUT4 unary_minus_10_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n37784), .O(n1095_adj_5231)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n37784), .I0(n1028), 
            .I1(VCC_net), .CO(n37785));
    SB_LUT4 i1_4_lut_adj_1582 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n45354), 
            .O(n45360));
    defparam i1_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5181));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33387_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n45360), 
            .O(n2445));
    defparam i33387_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n37783), .O(n1096_adj_5232)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4551_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(107[7:14])
    defparam i4551_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5268));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1520_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2625_5 (.CI(n37525), .I0(n623), .I1(VCC_net), .CO(n37526));
    SB_LUT4 encoder0_position_31__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23), .I2(encoder0_position[31]), .I3(GND_net), .O(n948));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5182));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32296_3_lut (.I0(n2247), .I1(n2148), .I2(n2049), .I3(GND_net), 
            .O(n47428));
    defparam i32296_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 encoder0_position_31__I_0_i1383_rep_46_3_lut (.I0(n2095), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n45760));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1383_rep_46_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1450_rep_45_3_lut (.I0(n45760), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n45757));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1450_rep_45_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1518_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33168_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48300));
    defparam i33168_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1519_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14646_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n27617), .I3(GND_net), .O(n28160));   // verilog/coms.v(127[12] 300[6])
    defparam i14646_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1583 (.I0(n2323), .I1(n2327), .I2(n2326), .I3(n2325), 
            .O(n45074));
    defparam i1_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(n2322), .I1(n2328), .I2(n2324), .I3(GND_net), 
            .O(n45076));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i20591_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n34102));
    defparam i20591_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1584 (.I0(n2320), .I1(n2321), .I2(n45076), .I3(n45074), 
            .O(n45082));
    defparam i1_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1585 (.I0(n2329), .I1(n2330), .I2(GND_net), .I3(GND_net), 
            .O(n45330));
    defparam i1_2_lut_adj_1585.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1586 (.I0(n45330), .I1(n2319), .I2(n45082), .I3(n34102), 
            .O(n45086));
    defparam i1_4_lut_adj_1586.LUT_INIT = 16'hfefc;
    SB_LUT4 i19677_2_lut (.I0(pwm_out), .I1(GHC), .I2(GND_net), .I3(GND_net), 
            .O(INHC_c_0));   // verilog/TinyFPGA_B.v(84[16:31])
    defparam i19677_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1587 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n45086), 
            .O(n45092));
    defparam i1_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i33421_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n45092), 
            .O(n2346));
    defparam i33421_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19676_2_lut (.I0(pwm_out), .I1(GHB), .I2(GND_net), .I3(GND_net), 
            .O(INHB_c_0));   // verilog/TinyFPGA_B.v(82[16:31])
    defparam i19676_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19974_2_lut (.I0(pwm_out), .I1(GHA), .I2(GND_net), .I3(GND_net), 
            .O(INHA_c_0));   // verilog/TinyFPGA_B.v(80[16:31])
    defparam i19974_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22), .I2(encoder0_position[31]), .I3(GND_net), .O(n947));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33097_1_lut (.I0(n34196), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48229));
    defparam i33097_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32470_3_lut (.I0(n45773), .I1(n1827), .I2(n47436), .I3(GND_net), 
            .O(n2124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32470_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32471_3_lut (.I0(n2124), .I1(n2191), .I2(n2148), .I3(GND_net), 
            .O(n2223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32471_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2188_3_lut (.I0(n3217), .I1(n3284), 
            .I2(n3237), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2194_3_lut (.I0(n3223), .I1(n3290), 
            .I2(n3237), .I3(GND_net), .O(n25_adj_5292));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2200_3_lut (.I0(n3229), .I1(n3296), 
            .I2(n3237), .I3(GND_net), .O(n13_adj_5288));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32472_3_lut (.I0(n2028), .I1(n2095), .I2(n2049), .I3(GND_net), 
            .O(n2127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32472_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5290));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2196_3_lut (.I0(n3225), .I1(n3292), 
            .I2(n3237), .I3(GND_net), .O(n21_adj_5291));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1588 (.I0(n3220), .I1(n21_adj_5291), .I2(n3287), 
            .I3(n3237), .O(n44848));
    defparam i1_4_lut_adj_1588.LUT_INIT = 16'heefc;
    SB_LUT4 i32473_3_lut (.I0(n2127), .I1(n2194), .I2(n2148), .I3(GND_net), 
            .O(n2226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32473_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1589 (.I0(n2226), .I1(n2224), .I2(n2225), .I3(n2227), 
            .O(n45308));
    defparam i1_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5289));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20532_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n34042));
    defparam i20532_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1590 (.I0(n3219), .I1(n37), .I2(n3286), .I3(n3237), 
            .O(n44852));
    defparam i1_4_lut_adj_1590.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1591 (.I0(n2222), .I1(n45308), .I2(n2223), .I3(n2228), 
            .O(n45312));
    defparam i1_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1592 (.I0(n2229), .I1(n34042), .I2(n2230), .I3(n2231), 
            .O(n43363));
    defparam i1_4_lut_adj_1592.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1593 (.I0(n3222), .I1(n25_adj_5292), .I2(n3289), 
            .I3(n3237), .O(n44850));
    defparam i1_4_lut_adj_1593.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1594 (.I0(n2220), .I1(n43363), .I2(n2221), .I3(n45312), 
            .O(n45318));
    defparam i1_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1595 (.I0(n2217), .I1(n2218), .I2(n2219), .I3(n45318), 
            .O(n45324));
    defparam i1_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i32745_4_lut (.I0(n2215), .I1(n2214), .I2(n2216), .I3(n45324), 
            .O(n2247));
    defparam i32745_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14647_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n27617), .I3(GND_net), .O(n28161));   // verilog/coms.v(127[12] 300[6])
    defparam i14647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14648_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n27617), .I3(GND_net), .O(n28162));   // verilog/coms.v(127[12] 300[6])
    defparam i14648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14649_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n27617), .I3(GND_net), .O(n28163));   // verilog/coms.v(127[12] 300[6])
    defparam i14649_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2187_3_lut (.I0(n3216), .I1(n3283), 
            .I2(n3237), .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2187_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1596 (.I0(n44848), .I1(n3221), .I2(n3288), .I3(n3237), 
            .O(n44860));
    defparam i1_4_lut_adj_1596.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_31__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1597 (.I0(n3218), .I1(n13_adj_5288), .I2(n3285), 
            .I3(n3237), .O(n44854));
    defparam i1_4_lut_adj_1597.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1598 (.I0(n3224), .I1(n17_adj_5290), .I2(n3291), 
            .I3(n3237), .O(n44858));
    defparam i1_4_lut_adj_1598.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1389_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1599 (.I0(n3226), .I1(n15_adj_5289), .I2(n3293), 
            .I3(n3237), .O(n44856));
    defparam i1_4_lut_adj_1599.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1600 (.I0(n44860), .I1(n39), .I2(n44850), .I3(n44852), 
            .O(n44870));
    defparam i1_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21), .I2(encoder0_position[31]), .I3(GND_net), .O(n946));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32304_3_lut (.I0(n2049), .I1(n1950), .I2(n1851), .I3(GND_net), 
            .O(n47436));
    defparam i32304_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 i1_4_lut_adj_1601 (.I0(n44870), .I1(n44856), .I2(n44858), 
            .I3(n44854), .O(n44872));
    defparam i1_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1246_rep_69_3_lut (.I0(n1894), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n45781));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1246_rep_69_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1313_rep_61_3_lut (.I0(n45781), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n45773));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1313_rep_61_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1602 (.I0(n3215), .I1(n44872), .I2(n3282), .I3(n3237), 
            .O(n44874));
    defparam i1_4_lut_adj_1602.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20396_4_lut (.I0(n652), .I1(n957), .I2(n3301), .I3(n3237), 
            .O(n33903));
    defparam i20396_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_31__I_0_i2203_3_lut (.I0(n3232), .I1(n3299), 
            .I2(n3237), .I3(GND_net), .O(n7_adj_5287));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2203_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n46883), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5240));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1603 (.I0(n3214), .I1(n44874), .I2(n3281), .I3(n3237), 
            .O(n44876));
    defparam i1_4_lut_adj_1603.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20508_4_lut (.I0(n33903), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n34018));
    defparam i20508_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 encoder0_position_31__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32785_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n47917));
    defparam i32785_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1604 (.I0(n34018), .I1(n44876), .I2(n5_adj_5240), 
            .I3(n7_adj_5287), .O(n44878));
    defparam i1_4_lut_adj_1604.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1605 (.I0(n2126), .I1(n2128), .I2(n2127), .I3(GND_net), 
            .O(n45000));
    defparam i1_3_lut_adj_1605.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_adj_1606 (.I0(n2123), .I1(n2125), .I2(n2124), .I3(GND_net), 
            .O(n45002));
    defparam i1_3_lut_adj_1606.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1607 (.I0(n3213), .I1(n44878), .I2(n3280), .I3(n3237), 
            .O(n44880));
    defparam i1_4_lut_adj_1607.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1608 (.I0(n3212), .I1(n44880), .I2(n3279), .I3(n3237), 
            .O(n44882));
    defparam i1_4_lut_adj_1608.LUT_INIT = 16'heefc;
    SB_LUT4 i20595_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n34106));
    defparam i20595_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1609 (.I0(n2121), .I1(n2122), .I2(n45002), .I3(n45000), 
            .O(n45008));
    defparam i1_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1610 (.I0(n3211), .I1(n44882), .I2(n3278), .I3(n3237), 
            .O(n44884));
    defparam i1_4_lut_adj_1610.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1611 (.I0(n3210), .I1(n44884), .I2(n3277), .I3(n3237), 
            .O(n44886));
    defparam i1_4_lut_adj_1611.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1612 (.I0(n2129), .I1(n45008), .I2(n34106), .I3(n2130), 
            .O(n45010));
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1613 (.I0(n3209), .I1(n44886), .I2(n3276), .I3(n3237), 
            .O(n44888));
    defparam i1_4_lut_adj_1613.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1614 (.I0(n2118), .I1(n2119), .I2(n45010), .I3(n2120), 
            .O(n45016));
    defparam i1_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i32789_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n45016), 
            .O(n2148));
    defparam i32789_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1615 (.I0(n3208), .I1(n44888), .I2(n3275), .I3(n3237), 
            .O(n44890));
    defparam i1_4_lut_adj_1615.LUT_INIT = 16'heefc;
    SB_LUT4 i14784_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n23622), .I3(GND_net), .O(n28298));   // verilog/coms.v(127[12] 300[6])
    defparam i14784_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14785_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n23622), .I3(GND_net), .O(n28299));   // verilog/coms.v(127[12] 300[6])
    defparam i14785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1616 (.I0(n3207), .I1(n44890), .I2(n3274), .I3(n3237), 
            .O(n44892));
    defparam i1_4_lut_adj_1616.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1617 (.I0(n3206), .I1(n44892), .I2(n3273), .I3(n3237), 
            .O(n44894));
    defparam i1_4_lut_adj_1617.LUT_INIT = 16'heefc;
    SB_LUT4 i14786_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n23622), .I3(GND_net), .O(n28300));   // verilog/coms.v(127[12] 300[6])
    defparam i14786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1618 (.I0(n3205), .I1(n44894), .I2(n3272), .I3(n3237), 
            .O(n44896));
    defparam i1_4_lut_adj_1618.LUT_INIT = 16'heefc;
    SB_LUT4 i33100_4_lut (.I0(n44896), .I1(n3204), .I2(n3271), .I3(n3237), 
            .O(n34196));
    defparam i33100_4_lut.LUT_INIT = 16'h1105;
    SB_LUT4 encoder0_position_31__I_0_i1316_rep_67_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1316_rep_67_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1111_rep_84_3_lut (.I0(n1695), .I1(n1794), 
            .I2(n1752), .I3(GND_net), .O(n45796));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1111_rep_84_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14650_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n27617), .I3(GND_net), .O(n28164));   // verilog/coms.v(127[12] 300[6])
    defparam i14650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31769_2_lut (.I0(n1752), .I1(n1653), .I2(GND_net), .I3(GND_net), 
            .O(n46900));
    defparam i31769_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_31__I_0_i1178_rep_75_3_lut (.I0(n45796), .I1(n1893), 
            .I2(n1851), .I3(GND_net), .O(n45787));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1178_rep_75_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14651_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n41203), .I3(GND_net), .O(n28165));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32468_4_lut (.I0(n45787), .I1(n1628), .I2(n1851), .I3(n46900), 
            .O(n47600));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32468_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i32469_3_lut (.I0(n47600), .I1(n1992), .I2(n1950), .I3(GND_net), 
            .O(n2024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32469_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32360_3_lut (.I0(n1827), .I1(n1894), .I2(n1851), .I3(GND_net), 
            .O(n1926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32360_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32361_3_lut (.I0(n1926), .I1(n1993), .I2(n1950), .I3(GND_net), 
            .O(n2025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32361_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32362_3_lut (.I0(n1828), .I1(n1895), .I2(n1851), .I3(GND_net), 
            .O(n1927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32362_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32363_3_lut (.I0(n1927), .I1(n1994), .I2(n1950), .I3(GND_net), 
            .O(n2026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14787_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n23622), .I3(GND_net), .O(n28301));   // verilog/coms.v(127[12] 300[6])
    defparam i14787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20), .I2(encoder0_position[31]), .I3(GND_net), .O(n945));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32882_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48014));
    defparam i32882_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20536_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n34046));
    defparam i20536_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1619 (.I0(n2026), .I1(n2027), .I2(GND_net), .I3(GND_net), 
            .O(n45278));
    defparam i1_2_lut_adj_1619.LUT_INIT = 16'heeee;
    SB_LUT4 i14653_3_lut (.I0(h3), .I1(reg_B[0]), .I2(n44732), .I3(GND_net), 
            .O(n28167));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14653_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14654_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n44019), .I3(GND_net), .O(n28168));   // verilog/coms.v(127[12] 300[6])
    defparam i14654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1620 (.I0(n2025), .I1(n45278), .I2(n2024), .I3(n2028), 
            .O(n45282));
    defparam i1_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1621 (.I0(n2029), .I1(n34046), .I2(n2030), .I3(n2031), 
            .O(n43356));
    defparam i1_4_lut_adj_1621.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1622 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n45282), 
            .O(n45288));
    defparam i1_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1623 (.I0(n2019), .I1(n2020), .I2(n45288), .I3(n43356), 
            .O(n45294));
    defparam i1_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32885_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n45294), 
            .O(n2049));
    defparam i32885_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14655_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28169));   // verilog/coms.v(127[12] 300[6])
    defparam i14655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14659_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[1]), .I2(n5_adj_5186), 
            .I3(n26445), .O(n28173));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14659_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14660_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[2]), .I2(n5_adj_5196), 
            .I3(n26445), .O(n28174));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14660_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19), .I2(encoder0_position[31]), .I3(GND_net), .O(n944));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5269), .I3(n38442), .O(n16_adj_5151)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14661_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[3]), .I2(n33328), 
            .I3(n26445), .O(n28175));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14661_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14662_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[4]), .I2(n9_adj_5198), 
            .I3(n26440), .O(n28176));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14662_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14663_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[5]), .I2(n5_adj_5186), 
            .I3(n26440), .O(n28177));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14663_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32379_3_lut (.I0(n1727), .I1(n1794), .I2(n1752), .I3(GND_net), 
            .O(n1826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14664_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[6]), .I2(n5_adj_5196), 
            .I3(n26440), .O(n28178));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14664_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32357_3_lut (.I0(n1826), .I1(n1893), .I2(n1851), .I3(GND_net), 
            .O(n1925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32357_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14665_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[7]), .I2(n33328), 
            .I3(n26440), .O(n28179));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14665_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n37783), .I0(n1029), 
            .I1(GND_net), .CO(n37784));
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n37782), .O(n1097_adj_5233)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14666_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[8]), .I2(n9_adj_5198), 
            .I3(n26435), .O(n28180));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14666_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n37782), .I0(n1030), 
            .I1(GND_net), .CO(n37783));
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n37781), .O(n1098_adj_5234)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14667_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[9]), .I2(n5_adj_5186), 
            .I3(n26435), .O(n28181));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14667_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14668_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[10]), .I2(n5_adj_5196), 
            .I3(n26435), .O(n28182));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14668_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14669_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[11]), .I2(n33328), 
            .I3(n26435), .O(n28183));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14669_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14670_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[12]), .I2(n9_adj_5198), 
            .I3(n26432), .O(n28184));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14670_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32381_3_lut (.I0(n1726), .I1(n1793), .I2(n1752), .I3(GND_net), 
            .O(n1825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32355_3_lut (.I0(n1825), .I1(n1892), .I2(n1851), .I3(GND_net), 
            .O(n1924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32355_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32906_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48038));
    defparam i32906_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1624 (.I0(n1927), .I1(n1926), .I2(n1925), .I3(n1928), 
            .O(n44978));
    defparam i1_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20538_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n34048));
    defparam i20538_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1625 (.I0(n1922), .I1(n1923), .I2(n44978), .I3(n1924), 
            .O(n44984));
    defparam i1_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14671_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[15]), .I2(n33328), 
            .I3(n26432), .O(n28185));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14671_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_4_lut_adj_1626 (.I0(n1929), .I1(n34048), .I2(n1930), .I3(n1931), 
            .O(n43320));
    defparam i1_4_lut_adj_1626.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n37781), .I0(n1031), 
            .I1(VCC_net), .CO(n37782));
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n37780), .O(n1099_adj_5235)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n38443), 
            .I0(GND_net), .I1(n15_adj_5268), .CO(n38444));
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n37780), .I0(n1032), 
            .I1(GND_net), .CO(n37781));
    SB_DFFSR pwm_setpoint__i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_23__N_191[0]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5268), .I3(n38443), .O(n15_adj_5187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n37779), .O(n1100_adj_5236)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14673_4_lut (.I0(state_7__N_4103[3]), .I1(data[1]), .I2(n10_adj_5251), 
            .I3(n26424), .O(n28187));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14673_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14674_4_lut (.I0(state_7__N_4103[3]), .I1(data[2]), .I2(n4_adj_5218), 
            .I3(n26409), .O(n28188));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14674_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i33130_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48262));
    defparam i33130_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1627 (.I0(n1920), .I1(n43320), .I2(n1921), .I3(n44984), 
            .O(n44990));
    defparam i1_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i32909_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n44990), 
            .O(n1950));
    defparam i32909_4_lut.LUT_INIT = 16'h0001;
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n7072), 
            .D(n1088), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14675_4_lut (.I0(state_7__N_4103[3]), .I1(data[3]), .I2(n4_adj_5218), 
            .I3(n26424), .O(n28189));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14675_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1628 (.I0(n3220), .I1(n3225), .I2(n3221), .I3(n3219), 
            .O(n45490));
    defparam i1_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i14676_4_lut (.I0(state_7__N_4103[3]), .I1(data[4]), .I2(n4_adj_5192), 
            .I3(n26409), .O(n28190));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14676_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n38444), 
            .I0(GND_net), .I1(n14_adj_5267), .CO(n38445));
    SB_LUT4 i14677_4_lut (.I0(state_7__N_4103[3]), .I1(data[5]), .I2(n4_adj_5192), 
            .I3(n26424), .O(n28191));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14677_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2625_4_lut (.I0(GND_net), .I1(n405), .I2(GND_net), .I3(n37524), 
            .O(n7649)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n7072), 
            .D(n1096), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n37779), .I0(n1033), 
            .I1(VCC_net), .CO(n37780));
    SB_LUT4 i14678_4_lut (.I0(state_7__N_4103[3]), .I1(data[6]), .I2(n33292), 
            .I3(n26409), .O(n28192));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14678_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101_adj_5237)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n7072), 
            .D(n1095), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i20573_4_lut (.I0(n957), .I1(n3231), .I2(n3232), .I3(n3233), 
            .O(n34084));
    defparam i20573_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14679_4_lut (.I0(state_7__N_4103[3]), .I1(data[7]), .I2(n33292), 
            .I3(n26424), .O(n28193));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14679_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i1_3_lut_adj_1629 (.I0(n3216), .I1(n3218), .I2(n45490), .I3(GND_net), 
            .O(n45494));
    defparam i1_3_lut_adj_1629.LUT_INIT = 16'hfefe;
    SB_LUT4 i14681_4_lut (.I0(n43011), .I1(state[1]), .I2(state_3__N_528[1]), 
            .I3(n27791), .O(n28195));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14681_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2625_4 (.CI(n37524), .I0(n405), .I1(GND_net), .CO(n37525));
    SB_LUT4 i14682_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_5200), 
            .I3(n26390), .O(n28196));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14682_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14683_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_5184), 
            .I3(n26398), .O(n28197));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14683_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5267), .I3(n38444), .O(n14_adj_5188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14684_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_5184), 
            .I3(n26390), .O(n28198));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14684_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n38445), 
            .I0(GND_net), .I1(n13_adj_5266), .CO(n38446));
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n37779));
    SB_LUT4 i1_2_lut_adj_1630 (.I0(n3229), .I1(n3230), .I2(GND_net), .I3(GND_net), 
            .O(n45546));
    defparam i1_2_lut_adj_1630.LUT_INIT = 16'h8888;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n38446), 
            .I0(GND_net), .I1(n12_adj_5265), .CO(n38447));
    SB_LUT4 add_2625_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n37523), 
            .O(n7650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5266), .I3(n38445), .O(n13_adj_5189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1631 (.I0(n3228), .I1(n3226), .I2(n3223), .I3(n3222), 
            .O(n45510));
    defparam i1_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1180_rep_77_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1180_rep_77_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1632 (.I0(n3217), .I1(n45510), .I2(n3227), .I3(n3224), 
            .O(n45514));
    defparam i1_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1633 (.I0(n3213), .I1(n3214), .I2(n3215), .I3(n45514), 
            .O(n45520));
    defparam i1_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 add_224_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n37450), .O(encoder1_position_scaled_23__N_75[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n37778), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n37777), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14685_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_5199), 
            .I3(n26398), .O(n28199));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14685_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n37777), .I0(n928), 
            .I1(VCC_net), .CO(n37778));
    SB_CARRY add_224_7 (.CI(n37450), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n37451));
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n37776), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n7072), 
            .D(n1087), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY add_2625_3 (.CI(n37523), .I0(n625), .I1(VCC_net), .CO(n37524));
    SB_LUT4 add_2625_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n7651)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1634 (.I0(n3209), .I1(n3210), .I2(n3211), .I3(n45520), 
            .O(n45526));
    defparam i1_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n37776), .I0(n929), 
            .I1(GND_net), .CO(n37777));
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1635 (.I0(n3212), .I1(n45546), .I2(n45494), .I3(n34084), 
            .O(n45498));
    defparam i1_4_lut_adj_1635.LUT_INIT = 16'hfefa;
    SB_LUT4 add_224_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n37468), .O(encoder1_position_scaled_23__N_75[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2625_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n37523));
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n37775), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n7072), 
            .D(n1108), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 unary_minus_10_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_setpoint_23__N_215), 
            .I3(n37522), .O(pwm_setpoint_23__N_191[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n37467), .O(encoder1_position_scaled_23__N_75[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n37775), .I0(n930), 
            .I1(GND_net), .CO(n37776));
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n37774), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n37774), .I0(n931), 
            .I1(VCC_net), .CO(n37775));
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n37773), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1636 (.I0(n3207), .I1(n3206), .I2(n3208), .I3(n45526), 
            .O(n44592));
    defparam i1_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18), .I2(encoder0_position[31]), .I3(GND_net), .O(n943));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32932_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48064));
    defparam i32932_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33134_4_lut (.I0(n3205), .I1(n44592), .I2(n3204), .I3(n45498), 
            .O(n3237));
    defparam i33134_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1637 (.I0(n1825), .I1(n1828), .I2(n1826), .I3(n1827), 
            .O(n45252));
    defparam i1_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i20544_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n34054));
    defparam i20544_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1638 (.I0(n1823), .I1(n1824), .I2(n45252), .I3(GND_net), 
            .O(n45256));
    defparam i1_3_lut_adj_1638.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1639 (.I0(n1829), .I1(n34054), .I2(n1830), .I3(n1831), 
            .O(n43335));
    defparam i1_4_lut_adj_1639.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i2041_3_lut (.I0(n3006), .I1(n3073), 
            .I2(n3039), .I3(GND_net), .O(n3105));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2041_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n7072), 
            .D(n1086), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1640 (.I0(n1821), .I1(n1822), .I2(n43335), .I3(n45256), 
            .O(n45262));
    defparam i1_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i32935_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n45262), 
            .O(n1851));
    defparam i32935_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n37773), .I0(n932), 
            .I1(GND_net), .CO(n37774));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5279), .I3(n38432), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n37772), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5280), .I3(n38431), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15167_3_lut (.I0(current[12]), .I1(data_adj_5353[12]), .I2(n43722), 
            .I3(GND_net), .O(n28681));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15168_3_lut (.I0(current[11]), .I1(data_adj_5353[11]), .I2(n43722), 
            .I3(GND_net), .O(n28682));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5272));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14790_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n23622), .I3(GND_net), .O(n28304));   // verilog/coms.v(127[12] 300[6])
    defparam i14790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14791_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n23622), .I3(GND_net), .O(n28305));   // verilog/coms.v(127[12] 300[6])
    defparam i14791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14686_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_5199), 
            .I3(n26390), .O(n28200));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14686_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14792_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n23622), .I3(GND_net), .O(n28306));   // verilog/coms.v(127[12] 300[6])
    defparam i14792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14793_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n44019), 
            .I3(GND_net), .O(n28307));   // verilog/coms.v(127[12] 300[6])
    defparam i14793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15169_3_lut (.I0(current[10]), .I1(data_adj_5353[10]), .I2(n43722), 
            .I3(GND_net), .O(n28683));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14642_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n27617), .I3(GND_net), .O(n28156));   // verilog/coms.v(127[12] 300[6])
    defparam i14642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[20]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14794_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n23622), .I3(GND_net), .O(n28308));   // verilog/coms.v(127[12] 300[6])
    defparam i14794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14687_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n33332), 
            .I3(n26398), .O(n28201));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14687_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i14795_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n44019), 
            .I3(GND_net), .O(n28309));   // verilog/coms.v(127[12] 300[6])
    defparam i14795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n37772), .I0(n933), 
            .I1(VCC_net), .CO(n37773));
    SB_LUT4 i15170_3_lut (.I0(current[9]), .I1(data_adj_5353[9]), .I2(n43722), 
            .I3(GND_net), .O(n28684));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15171_3_lut (.I0(current[8]), .I1(data_adj_5353[8]), .I2(n43722), 
            .I3(GND_net), .O(n28685));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15171_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n38432), 
            .I0(GND_net), .I1(n26_adj_5279), .CO(n38433));
    SB_LUT4 i4798_2_lut (.I0(n2_adj_5227), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4798_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15172_3_lut (.I0(current[7]), .I1(data_adj_5353[7]), .I2(n43722), 
            .I3(GND_net), .O(n28686));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14796_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n44019), 
            .I3(GND_net), .O(n28310));   // verilog/coms.v(127[12] 300[6])
    defparam i14796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n38433), 
            .I0(GND_net), .I1(n25_adj_5278), .CO(n38434));
    SB_LUT4 i14797_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n44019), 
            .I3(GND_net), .O(n28311));   // verilog/coms.v(127[12] 300[6])
    defparam i14797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15173_3_lut (.I0(current[6]), .I1(data_adj_5353[6]), .I2(n43722), 
            .I3(GND_net), .O(n28687));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14798_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n23622), .I3(GND_net), .O(n28312));   // verilog/coms.v(127[12] 300[6])
    defparam i14798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14799_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n23622), .I3(GND_net), .O(n28313));   // verilog/coms.v(127[12] 300[6])
    defparam i14799_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[21]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15174_3_lut (.I0(current[5]), .I1(data_adj_5353[5]), .I2(n43722), 
            .I3(GND_net), .O(n28688));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5278), .I3(n38433), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n37772));
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n37771), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n37770), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n37770), .I0(n829), 
            .I1(GND_net), .CO(n37771));
    SB_LUT4 i14800_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n44019), 
            .I3(GND_net), .O(n28314));   // verilog/coms.v(127[12] 300[6])
    defparam i14800_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14801_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_4087[0]), 
            .I3(enable_slow_N_4190), .O(n28315));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14801_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i15175_3_lut (.I0(current[4]), .I1(data_adj_5353[4]), .I2(n43722), 
            .I3(GND_net), .O(n28689));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n37769), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n37769), .I0(n830), 
            .I1(GND_net), .CO(n37770));
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n37768), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_238_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[22]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14802_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28316));   // verilog/coms.v(127[12] 300[6])
    defparam i14802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14803_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n23622), .I3(GND_net), .O(n28317));   // verilog/coms.v(127[12] 300[6])
    defparam i14803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[23]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15176_3_lut (.I0(current[3]), .I1(data_adj_5353[3]), .I2(n43722), 
            .I3(GND_net), .O(n28690));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n3), 
            .I3(n37521), .O(pwm_setpoint_23__N_191[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n37768), .I0(n831), 
            .I1(VCC_net), .CO(n37769));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n38434), 
            .I0(GND_net), .I1(n24_adj_5277), .CO(n38435));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5277), .I3(n38434), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n38435), 
            .I0(GND_net), .I1(n23_adj_5276), .CO(n38436));
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5276), .I3(n38435), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_24 (.CI(n37521), .I0(GND_net), .I1(n3), 
            .CO(n37522));
    SB_LUT4 unary_minus_10_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n4), 
            .I3(n37520), .O(pwm_setpoint_23__N_191[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15177_3_lut (.I0(current[2]), .I1(data_adj_5353[2]), .I2(n43722), 
            .I3(GND_net), .O(n28691));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15177_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_24 (.CI(n37467), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n37468));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n38436), 
            .I0(GND_net), .I1(n22_adj_5275), .CO(n38437));
    SB_LUT4 add_224_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n37466), .O(encoder1_position_scaled_23__N_75[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5275), .I3(n38436), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n38437), 
            .I0(GND_net), .I1(n21_adj_5274), .CO(n38438));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5265), .I3(n38446), .O(n12_adj_5202)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n37449), .O(encoder1_position_scaled_23__N_75[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632_adj_5239), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_23 (.CI(n37466), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n37467));
    SB_LUT4 add_224_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n37465), .O(encoder1_position_scaled_23__N_75[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n37767), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n37767), .I0(n832), 
            .I1(GND_net), .CO(n37768));
    SB_LUT4 i15178_3_lut (.I0(current[1]), .I1(data_adj_5353[1]), .I2(n43722), 
            .I3(GND_net), .O(n28692));   // verilog/tli4970.v(33[10] 66[6])
    defparam i15178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n37766), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_22 (.CI(n37465), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n37466));
    SB_LUT4 add_224_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n37464), .O(encoder1_position_scaled_23__N_75[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n37766), .I0(n833), 
            .I1(VCC_net), .CO(n37767));
    SB_CARRY add_224_21 (.CI(n37464), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n37465));
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n37463), .O(encoder1_position_scaled_23__N_75[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_23 (.CI(n37520), .I0(GND_net), .I1(n4), 
            .CO(n37521));
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14805_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n44019), 
            .I3(GND_net), .O(n28319));   // verilog/coms.v(127[12] 300[6])
    defparam i14805_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17), .I2(encoder0_position[31]), .I3(GND_net), .O(n942));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_20 (.CI(n37463), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n37464));
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n5), 
            .I3(n37519), .O(pwm_setpoint_23__N_191[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n37462), .O(encoder1_position_scaled_23__N_75[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_19 (.CI(n37462), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n37463));
    SB_LUT4 add_224_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n37461), .O(encoder1_position_scaled_23__N_75[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14806_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n23622), 
            .I3(GND_net), .O(n28320));   // verilog/coms.v(127[12] 300[6])
    defparam i14806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32956_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48088));
    defparam i32956_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14807_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n23622), 
            .I3(GND_net), .O(n28321));   // verilog/coms.v(127[12] 300[6])
    defparam i14807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33059_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48191));
    defparam i33059_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14808_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n23622), 
            .I3(GND_net), .O(n28322));   // verilog/coms.v(127[12] 300[6])
    defparam i14808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14809_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n23622), 
            .I3(GND_net), .O(n28323));   // verilog/coms.v(127[12] 300[6])
    defparam i14809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14810_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28324));   // verilog/coms.v(127[12] 300[6])
    defparam i14810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14811_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n23622), 
            .I3(GND_net), .O(n28325));   // verilog/coms.v(127[12] 300[6])
    defparam i14811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14812_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n23622), 
            .I3(GND_net), .O(n28326));   // verilog/coms.v(127[12] 300[6])
    defparam i14812_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_18 (.CI(n37461), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n37462));
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n37766));
    SB_LUT4 i14813_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n23622), 
            .I3(GND_net), .O(n28327));   // verilog/coms.v(127[12] 300[6])
    defparam i14813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14814_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28328));   // verilog/coms.v(127[12] 300[6])
    defparam i14814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_224_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n37460), .O(encoder1_position_scaled_23__N_75[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14815_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n23622), 
            .I3(GND_net), .O(n28329));   // verilog/coms.v(127[12] 300[6])
    defparam i14815_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_22 (.CI(n37519), .I0(GND_net), .I1(n5), 
            .CO(n37520));
    SB_LUT4 i1_3_lut_adj_1641 (.I0(n1727), .I1(n1728), .I2(n1726), .I3(GND_net), 
            .O(n45100));
    defparam i1_3_lut_adj_1641.LUT_INIT = 16'hfefe;
    SB_LUT4 i20607_4_lut (.I0(n942), .I1(n1731), .I2(n1732), .I3(n1733), 
            .O(n34118));
    defparam i20607_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 unary_minus_10_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n6_adj_5138), 
            .I3(n37518), .O(pwm_setpoint_23__N_191[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1642 (.I0(n1723), .I1(n1724), .I2(n45100), .I3(n1725), 
            .O(n45106));
    defparam i1_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1643 (.I0(n1729), .I1(n1730), .I2(GND_net), .I3(GND_net), 
            .O(n45242));
    defparam i1_2_lut_adj_1643.LUT_INIT = 16'h8888;
    SB_LUT4 i14816_4_lut (.I0(state_7__N_4103[3]), .I1(data[0]), .I2(n10_adj_5251), 
            .I3(n26409), .O(n28330));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14816_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14817_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n23622), 
            .I3(GND_net), .O(n28331));   // verilog/coms.v(127[12] 300[6])
    defparam i14817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14821_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n23622), 
            .I3(GND_net), .O(n28335));   // verilog/coms.v(127[12] 300[6])
    defparam i14821_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut_adj_1644 (.I0(state_adj_5377[0]), .I1(n46890), .I2(n6692), 
            .I3(n33185), .O(n8_adj_5241));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_adj_1644.LUT_INIT = 16'h3afa;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62_adj_5244), 
            .I2(delay_counter[31]), .I3(\ID_READOUT_FSM.state [0]), .O(n44724));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i14826_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28340));   // verilog/coms.v(127[12] 300[6])
    defparam i14826_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_10_add_3_21 (.CI(n37518), .I0(GND_net), .I1(n6_adj_5138), 
            .CO(n37519));
    SB_LUT4 i14827_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28341));   // verilog/coms.v(127[12] 300[6])
    defparam i14827_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1645 (.I0(n45242), .I1(n1722), .I2(n45106), .I3(n34118), 
            .O(n45110));
    defparam i1_4_lut_adj_1645.LUT_INIT = 16'hfefc;
    SB_LUT4 i32959_4_lut (.I0(n1720), .I1(n1719), .I2(n1721), .I3(n45110), 
            .O(n1752));
    defparam i32959_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_10_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n7), 
            .I3(n37517), .O(pwm_setpoint_23__N_191[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14828_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28342));   // verilog/coms.v(127[12] 300[6])
    defparam i14828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_145_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n37425), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_6 (.CI(n37449), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n37450));
    SB_LUT4 i14829_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n23622), 
            .I3(GND_net), .O(n28343));   // verilog/coms.v(127[12] 300[6])
    defparam i14829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14830_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n23622), 
            .I3(GND_net), .O(n28344));   // verilog/coms.v(127[12] 300[6])
    defparam i14830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14831_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n23622), 
            .I3(GND_net), .O(n28345));   // verilog/coms.v(127[12] 300[6])
    defparam i14831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14832_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n23622), 
            .I3(GND_net), .O(n28346));   // verilog/coms.v(127[12] 300[6])
    defparam i14832_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14833_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n23622), 
            .I3(GND_net), .O(n28347));   // verilog/coms.v(127[12] 300[6])
    defparam i14833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15193_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n42288), 
            .I3(GND_net), .O(n28707));   // verilog/coms.v(127[12] 300[6])
    defparam i15193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15194_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n42288), 
            .I3(GND_net), .O(n28708));   // verilog/coms.v(127[12] 300[6])
    defparam i15194_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14834_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n23622), 
            .I3(GND_net), .O(n28348));   // verilog/coms.v(127[12] 300[6])
    defparam i14834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15195_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n42288), 
            .I3(GND_net), .O(n28709));   // verilog/coms.v(127[12] 300[6])
    defparam i15195_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14835_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n23622), 
            .I3(GND_net), .O(n28349));   // verilog/coms.v(127[12] 300[6])
    defparam i14835_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14836_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n23622), 
            .I3(GND_net), .O(n28350));   // verilog/coms.v(127[12] 300[6])
    defparam i14836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15196_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n42288), 
            .I3(GND_net), .O(n28710));   // verilog/coms.v(127[12] 300[6])
    defparam i15196_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15197_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n42288), 
            .I3(GND_net), .O(n28711));   // verilog/coms.v(127[12] 300[6])
    defparam i15197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14837_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n23622), 
            .I3(GND_net), .O(n28351));   // verilog/coms.v(127[12] 300[6])
    defparam i14837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14838_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n23622), 
            .I3(GND_net), .O(n28352));   // verilog/coms.v(127[12] 300[6])
    defparam i14838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15198_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n42288), 
            .I3(GND_net), .O(n28712));   // verilog/coms.v(127[12] 300[6])
    defparam i15198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14839_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n23622), 
            .I3(GND_net), .O(n28353));   // verilog/coms.v(127[12] 300[6])
    defparam i14839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15199_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n42288), 
            .I3(GND_net), .O(n28713));   // verilog/coms.v(127[12] 300[6])
    defparam i15199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14840_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n23622), 
            .I3(GND_net), .O(n28354));   // verilog/coms.v(127[12] 300[6])
    defparam i14840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_IO CS_MISO_pad (.PACKAGE_PIN(CS_MISO), .OUTPUT_ENABLE(VCC_net), .D_IN_0(CS_MISO_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_MISO_pad.PIN_TYPE = 6'b000001;
    defparam CS_MISO_pad.PULLUP = 1'b0;
    defparam CS_MISO_pad.NEG_TRIGGER = 1'b0;
    defparam CS_MISO_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i14841_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n23622), 
            .I3(GND_net), .O(n28355));   // verilog/coms.v(127[12] 300[6])
    defparam i14841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14842_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n23622), 
            .I3(GND_net), .O(n28356));   // verilog/coms.v(127[12] 300[6])
    defparam i14842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5365_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GHC_N_403));   // verilog/TinyFPGA_B.v(185[7] 204[14])
    defparam i5365_3_lut_4_lut.LUT_INIT = 16'h21cc;
    SB_LUT4 i14843_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n23622), .I3(GND_net), .O(n28357));   // verilog/coms.v(127[12] 300[6])
    defparam i14843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14844_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n23622), .I3(GND_net), .O(n28358));   // verilog/coms.v(127[12] 300[6])
    defparam i14844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14845_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n23622), .I3(GND_net), .O(n28359));   // verilog/coms.v(127[12] 300[6])
    defparam i14845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14846_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n23622), .I3(GND_net), .O(n28360));   // verilog/coms.v(127[12] 300[6])
    defparam i14846_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15200_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n42288), 
            .I3(GND_net), .O(n28714));   // verilog/coms.v(127[12] 300[6])
    defparam i15200_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14847_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n23622), .I3(GND_net), .O(n28361));   // verilog/coms.v(127[12] 300[6])
    defparam i14847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14848_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n23622), .I3(GND_net), .O(n28362));   // verilog/coms.v(127[12] 300[6])
    defparam i14848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632_adj_5239));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14849_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n23622), .I3(GND_net), .O(n28363));   // verilog/coms.v(127[12] 300[6])
    defparam i14849_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14850_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n23622), .I3(GND_net), .O(n28364));   // verilog/coms.v(127[12] 300[6])
    defparam i14850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14851_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n23622), .I3(GND_net), .O(n28365));   // verilog/coms.v(127[12] 300[6])
    defparam i14851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14852_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n23622), .I3(GND_net), .O(n28366));   // verilog/coms.v(127[12] 300[6])
    defparam i14852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14853_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n23622), .I3(GND_net), .O(n28367));   // verilog/coms.v(127[12] 300[6])
    defparam i14853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14854_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n23622), .I3(GND_net), .O(n28368));   // verilog/coms.v(127[12] 300[6])
    defparam i14854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14855_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n23622), .I3(GND_net), .O(n28369));   // verilog/coms.v(127[12] 300[6])
    defparam i14855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16_adj_5151), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n941));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32980_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48112));
    defparam i32980_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20548_3_lut (.I0(n941), .I1(n1632_adj_5239), .I2(n1633), 
            .I3(GND_net), .O(n34058));
    defparam i20548_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i14856_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n23622), .I3(GND_net), .O(n28370));   // verilog/coms.v(127[12] 300[6])
    defparam i14856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14857_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n23622), .I3(GND_net), .O(n28371));   // verilog/coms.v(127[12] 300[6])
    defparam i14857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1646 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n45230));
    defparam i1_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i14858_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n23622), .I3(GND_net), .O(n28372));   // verilog/coms.v(127[12] 300[6])
    defparam i14858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14859_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n23622), .I3(GND_net), .O(n28373));   // verilog/coms.v(127[12] 300[6])
    defparam i14859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14860_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n23622), .I3(GND_net), .O(n28374));   // verilog/coms.v(127[12] 300[6])
    defparam i14860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1647 (.I0(n1629), .I1(n34058), .I2(n1630), .I3(n1631), 
            .O(n43298));
    defparam i1_4_lut_adj_1647.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1648 (.I0(n1623), .I1(n43298), .I2(n1624), .I3(n45230), 
            .O(n45236));
    defparam i1_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i14861_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n23622), .I3(GND_net), .O(n28375));   // verilog/coms.v(127[12] 300[6])
    defparam i14861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32983_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n45236), 
            .O(n1653));
    defparam i32983_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14862_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n23622), .I3(GND_net), .O(n28376));   // verilog/coms.v(127[12] 300[6])
    defparam i14862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_10_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14863_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n23622), .I3(GND_net), .O(n28377));   // verilog/coms.v(127[12] 300[6])
    defparam i14863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14864_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n23622), .I3(GND_net), .O(n28378));   // verilog/coms.v(127[12] 300[6])
    defparam i14864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14865_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n44019), 
            .I3(GND_net), .O(n28379));   // verilog/coms.v(127[12] 300[6])
    defparam i14865_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_224_17 (.CI(n37460), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n37461));
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_145_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n37417), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14866_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n23622), .I3(GND_net), .O(n28380));   // verilog/coms.v(127[12] 300[6])
    defparam i14866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14867_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28381));   // verilog/coms.v(127[12] 300[6])
    defparam i14867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14868_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n44019), 
            .I3(GND_net), .O(n28382));   // verilog/coms.v(127[12] 300[6])
    defparam i14868_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14453_2_lut (.I0(n27644), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n27973));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i14453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32674_4_lut (.I0(commutation_state[1]), .I1(n23805), .I2(dti), 
            .I3(commutation_state[2]), .O(n27644));
    defparam i32674_4_lut.LUT_INIT = 16'hc5cf;
    SB_LUT4 add_224_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n37459), .O(encoder1_position_scaled_23__N_75[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14869_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n44019), 
            .I3(GND_net), .O(n28383));   // verilog/coms.v(127[12] 300[6])
    defparam i14869_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_20 (.CI(n37517), .I0(GND_net), .I1(n7), 
            .CO(n37518));
    SB_LUT4 i1_4_lut_adj_1649 (.I0(n3124), .I1(n3121), .I2(n3125), .I3(n3118), 
            .O(n45034));
    defparam i1_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33045_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48177));
    defparam i33045_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14870_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n23622), .I3(GND_net), .O(n28384));   // verilog/coms.v(127[12] 300[6])
    defparam i14870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1650 (.I0(n3119), .I1(n3117), .I2(n3128), .I3(n3127), 
            .O(n45038));
    defparam i1_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i14875_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n23622), .I3(GND_net), .O(n28389));   // verilog/coms.v(127[12] 300[6])
    defparam i14875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14876_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n23622), .I3(GND_net), .O(n28390));   // verilog/coms.v(127[12] 300[6])
    defparam i14876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14877_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n23622), .I3(GND_net), .O(n28391));   // verilog/coms.v(127[12] 300[6])
    defparam i14877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14878_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n23622), .I3(GND_net), .O(n28392));   // verilog/coms.v(127[12] 300[6])
    defparam i14878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14879_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n23622), .I3(GND_net), .O(n28393));   // verilog/coms.v(127[12] 300[6])
    defparam i14879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1651 (.I0(n3126), .I1(n3122), .I2(n3123), .I3(n3120), 
            .O(n45036));
    defparam i1_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14880_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n23622), .I3(GND_net), .O(n28394));   // verilog/coms.v(127[12] 300[6])
    defparam i14880_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_5187), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n940));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15209_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n42287), 
            .I3(GND_net), .O(n28723));   // verilog/coms.v(127[12] 300[6])
    defparam i15209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20512_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n34022));
    defparam i20512_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY add_224_16 (.CI(n37459), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n37460));
    SB_LUT4 dti_counter_2188_add_4_9_lut (.I0(n46835), .I1(n33280), .I2(dti_counter[7]), 
            .I3(n38246), .O(n48)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_9_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 add_224_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n37458), .O(encoder1_position_scaled_23__N_75[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14881_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n23622), .I3(GND_net), .O(n28395));   // verilog/coms.v(127[12] 300[6])
    defparam i14881_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_15 (.CI(n37458), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n37459));
    SB_LUT4 dti_counter_2188_add_4_8_lut (.I0(n46836), .I1(n33280), .I2(dti_counter[6]), 
            .I3(n38245), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_8_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i14882_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n23622), .I3(GND_net), .O(n28396));   // verilog/coms.v(127[12] 300[6])
    defparam i14882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14883_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n23622), .I3(GND_net), .O(n28397));   // verilog/coms.v(127[12] 300[6])
    defparam i14883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15210_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n42287), 
            .I3(GND_net), .O(n28724));   // verilog/coms.v(127[12] 300[6])
    defparam i15210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15211_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n42287), 
            .I3(GND_net), .O(n28725));   // verilog/coms.v(127[12] 300[6])
    defparam i15211_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_2188_add_4_8 (.CI(n38245), .I0(n33280), .I1(dti_counter[6]), 
            .CO(n38246));
    SB_LUT4 dti_counter_2188_add_4_7_lut (.I0(n46837), .I1(n33280), .I2(dti_counter[5]), 
            .I3(n38244), .O(n50)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_7_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 encoder0_position_31__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1652 (.I0(n3116), .I1(n45036), .I2(n45038), .I3(n45034), 
            .O(n45044));
    defparam i1_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i14884_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n23622), .I3(GND_net), .O(n28398));   // verilog/coms.v(127[12] 300[6])
    defparam i14884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14885_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n23622), .I3(GND_net), .O(n28399));   // verilog/coms.v(127[12] 300[6])
    defparam i14885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15212_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n42287), 
            .I3(GND_net), .O(n28726));   // verilog/coms.v(127[12] 300[6])
    defparam i15212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14886_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n23622), .I3(GND_net), .O(n28400));   // verilog/coms.v(127[12] 300[6])
    defparam i14886_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1653 (.I0(n3129), .I1(n34022), .I2(n3130), .I3(n3131), 
            .O(n43381));
    defparam i1_4_lut_adj_1653.LUT_INIT = 16'ha080;
    SB_LUT4 i15213_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n42287), 
            .I3(GND_net), .O(n28727));   // verilog/coms.v(127[12] 300[6])
    defparam i15213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14887_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n23622), .I3(GND_net), .O(n28401));   // verilog/coms.v(127[12] 300[6])
    defparam i14887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14888_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n23622), .I3(GND_net), .O(n28402));   // verilog/coms.v(127[12] 300[6])
    defparam i14888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32998_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48130));
    defparam i32998_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15214_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n42287), 
            .I3(GND_net), .O(n28728));   // verilog/coms.v(127[12] 300[6])
    defparam i15214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14889_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n23622), .I3(GND_net), .O(n28403));   // verilog/coms.v(127[12] 300[6])
    defparam i14889_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2188_add_4_7 (.CI(n38244), .I0(n33280), .I1(dti_counter[5]), 
            .CO(n38245));
    SB_LUT4 i1_4_lut_adj_1654 (.I0(n43381), .I1(n3114), .I2(n3115), .I3(n45044), 
            .O(n45050));
    defparam i1_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 dti_counter_2188_add_4_6_lut (.I0(n46838), .I1(n33280), .I2(dti_counter[4]), 
            .I3(n38243), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_6_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i14890_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n23622), .I3(GND_net), .O(n28404));   // verilog/coms.v(127[12] 300[6])
    defparam i14890_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15215_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n42287), 
            .I3(GND_net), .O(n28729));   // verilog/coms.v(127[12] 300[6])
    defparam i15215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14891_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n23622), .I3(GND_net), .O(n28405));   // verilog/coms.v(127[12] 300[6])
    defparam i14891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14892_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n23622), .I3(GND_net), .O(n28406));   // verilog/coms.v(127[12] 300[6])
    defparam i14892_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2188_add_4_6 (.CI(n38243), .I0(n33280), .I1(dti_counter[4]), 
            .CO(n38244));
    SB_LUT4 i14893_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n23622), .I3(GND_net), .O(n28407));   // verilog/coms.v(127[12] 300[6])
    defparam i14893_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14894_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n23622), .I3(GND_net), .O(n28408));   // verilog/coms.v(127[12] 300[6])
    defparam i14894_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15216_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n42287), 
            .I3(GND_net), .O(n28730));   // verilog/coms.v(127[12] 300[6])
    defparam i15216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1655 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n45050), 
            .O(n45056));
    defparam i1_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1656 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n45116));
    defparam i1_2_lut_adj_1656.LUT_INIT = 16'heeee;
    SB_LUT4 i14895_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n23622), .I3(GND_net), .O(n28409));   // verilog/coms.v(127[12] 300[6])
    defparam i14895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20611_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n34122));
    defparam i20611_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 dti_counter_2188_add_4_5_lut (.I0(n46839), .I1(n33280), .I2(dti_counter[3]), 
            .I3(n38242), .O(n52)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_5_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i14896_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n23622), .I3(GND_net), .O(n28410));   // verilog/coms.v(127[12] 300[6])
    defparam i14896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14897_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n23622), .I3(GND_net), .O(n28411));   // verilog/coms.v(127[12] 300[6])
    defparam i14897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14898_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n23622), .I3(GND_net), .O(n28412));   // verilog/coms.v(127[12] 300[6])
    defparam i14898_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2188_add_4_5 (.CI(n38242), .I0(n33280), .I1(dti_counter[3]), 
            .CO(n38243));
    SB_LUT4 i14899_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n23622), .I3(GND_net), .O(n28413));   // verilog/coms.v(127[12] 300[6])
    defparam i14899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14900_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n23622), .I3(GND_net), .O(n28414));   // verilog/coms.v(127[12] 300[6])
    defparam i14900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14901_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n23622), .I3(GND_net), .O(n28415));   // verilog/coms.v(127[12] 300[6])
    defparam i14901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1657 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n45116), 
            .O(n45122));
    defparam i1_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 dti_counter_2188_add_4_4_lut (.I0(n46840), .I1(n33280), .I2(dti_counter[2]), 
            .I3(n38241), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_4_lut.LUT_INIT = 16'hE22E;
    SB_LUT4 i1_4_lut_adj_1658 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n45056), 
            .O(n45062));
    defparam i1_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 i33171_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n45062), 
            .O(n3138));
    defparam i33171_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(n1529), .I1(n45122), .I2(n34122), .I3(n1530), 
            .O(n45124));
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'heccc;
    SB_LUT4 i33001_4_lut (.I0(n1522), .I1(n1521), .I2(n45124), .I3(n1523), 
            .O(n1554));
    defparam i33001_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14902_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n23622), .I3(GND_net), .O(n28416));   // verilog/coms.v(127[12] 300[6])
    defparam i14902_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY dti_counter_2188_add_4_4 (.CI(n38241), .I0(n33280), .I1(dti_counter[2]), 
            .CO(n38242));
    SB_LUT4 i14903_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n23622), .I3(GND_net), .O(n28417));   // verilog/coms.v(127[12] 300[6])
    defparam i14903_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14904_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n23622), .I3(GND_net), .O(n28418));   // verilog/coms.v(127[12] 300[6])
    defparam i14904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14905_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n23622), .I3(GND_net), .O(n28419));   // verilog/coms.v(127[12] 300[6])
    defparam i14905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 dti_counter_2188_add_4_3_lut (.I0(n46841), .I1(n33280), .I2(dti_counter[1]), 
            .I3(n38240), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_3_lut.LUT_INIT = 16'hE22E;
    SB_DFF dti_counter_2188__i7 (.Q(dti_counter[7]), .C(CLK_c), .D(n48));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i6 (.Q(dti_counter[6]), .C(CLK_c), .D(n49));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i5 (.Q(dti_counter[5]), .C(CLK_c), .D(n50));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i4 (.Q(dti_counter[4]), .C(CLK_c), .D(n51));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i3 (.Q(dti_counter[3]), .C(CLK_c), .D(n52));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i2 (.Q(dti_counter[2]), .C(CLK_c), .D(n53));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFF dti_counter_2188__i1 (.Q(dti_counter[1]), .C(CLK_c), .D(n54));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n7072), 
            .D(n1107), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i14906_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n23622), .I3(GND_net), .O(n28420));   // verilog/coms.v(127[12] 300[6])
    defparam i14906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY dti_counter_2188_add_4_3 (.CI(n38240), .I0(n33280), .I1(dti_counter[1]), 
            .CO(n38241));
    SB_LUT4 dti_counter_2188_add_4_2_lut (.I0(n46878), .I1(n1964), .I2(dti_counter[0]), 
            .I3(VCC_net), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam dti_counter_2188_add_4_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY dti_counter_2188_add_4_2 (.CI(VCC_net), .I0(n1964), .I1(dti_counter[0]), 
            .CO(n38240));
    SB_LUT4 encoder0_position_31__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n7072), 
            .D(n1094), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 add_2693_25_lut (.I0(n48205), .I1(n2_adj_5255), .I2(n1059), 
            .I3(n38239), .O(encoder0_position_scaled_23__N_51[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_2693_24_lut (.I0(n48191), .I1(n2_adj_5255), .I2(n1158), 
            .I3(n38238), .O(encoder0_position_scaled_23__N_51[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_24 (.CI(n38238), .I0(n2_adj_5255), .I1(n1158), .CO(n38239));
    SB_LUT4 i14907_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n23622), .I3(GND_net), .O(n28421));   // verilog/coms.v(127[12] 300[6])
    defparam i14907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14908_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n23622), .I3(GND_net), .O(n28422));   // verilog/coms.v(127[12] 300[6])
    defparam i14908_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n7072), 
            .D(n1106), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 add_2693_23_lut (.I0(n48177), .I1(n2_adj_5255), .I2(n1257), 
            .I3(n38237), .O(encoder0_position_scaled_23__N_51[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14909_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n23622), .I3(GND_net), .O(n28423));   // verilog/coms.v(127[12] 300[6])
    defparam i14909_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2693_23 (.CI(n38237), .I0(n2_adj_5255), .I1(n1257), .CO(n38238));
    SB_LUT4 i14910_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n44019), 
            .I3(GND_net), .O(n28424));   // verilog/coms.v(127[12] 300[6])
    defparam i14910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_22_lut (.I0(n48162), .I1(n2_adj_5255), .I2(n1356), 
            .I3(n38236), .O(encoder0_position_scaled_23__N_51[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i5367_3_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state[0]), .I3(dir), .O(GLC_N_412));   // verilog/TinyFPGA_B.v(185[7] 204[14])
    defparam i5367_3_lut_4_lut.LUT_INIT = 16'hcc21;
    SB_CARRY add_2693_22 (.CI(n38236), .I0(n2_adj_5255), .I1(n1356), .CO(n38237));
    SB_LUT4 i14911_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n23622), .I3(GND_net), .O(n28425));   // verilog/coms.v(127[12] 300[6])
    defparam i14911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_21_lut (.I0(n48147), .I1(n2_adj_5255), .I2(n1455), 
            .I3(n38235), .O(encoder0_position_scaled_23__N_51[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14912_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n44019), 
            .I3(GND_net), .O(n28426));   // verilog/coms.v(127[12] 300[6])
    defparam i14912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2693_21 (.CI(n38235), .I0(n2_adj_5255), .I1(n1455), .CO(n38236));
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_20_lut (.I0(n48130), .I1(n2_adj_5255), .I2(n1554), 
            .I3(n38234), .O(encoder0_position_scaled_23__N_51[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14913_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n44824), .I3(GND_net), 
            .O(n28427));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i14913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15225_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n42285), 
            .I3(GND_net), .O(n28739));   // verilog/coms.v(127[12] 300[6])
    defparam i15225_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15226_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n42285), 
            .I3(GND_net), .O(n28740));   // verilog/coms.v(127[12] 300[6])
    defparam i15226_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14914_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28428));   // verilog/coms.v(127[12] 300[6])
    defparam i14914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33030_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48162));
    defparam i33030_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14918_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28432));   // verilog/coms.v(127[12] 300[6])
    defparam i14918_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_145_13 (.CI(n37425), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n37426));
    SB_LUT4 encoder0_position_31__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2693_20 (.CI(n38234), .I0(n2_adj_5255), .I1(n1554), .CO(n38235));
    SB_LUT4 unary_minus_10_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n8), 
            .I3(n37516), .O(pwm_setpoint_23__N_191[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14919_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n23622), .I3(GND_net), .O(n28433));   // verilog/coms.v(127[12] 300[6])
    defparam i14919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14923_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_5200), 
            .I3(n26398), .O(n28437));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14923_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2693_19_lut (.I0(n48112), .I1(n2_adj_5255), .I2(n1653), 
            .I3(n38233), .O(encoder0_position_scaled_23__N_51[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14924_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n23622), .I3(GND_net), .O(n28438));   // verilog/coms.v(127[12] 300[6])
    defparam i14924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15227_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n42285), 
            .I3(GND_net), .O(n28741));   // verilog/coms.v(127[12] 300[6])
    defparam i15227_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14925_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n23622), .I3(GND_net), .O(n28439));   // verilog/coms.v(127[12] 300[6])
    defparam i14925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15228_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n42285), 
            .I3(GND_net), .O(n28742));   // verilog/coms.v(127[12] 300[6])
    defparam i15228_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14926_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n23622), .I3(GND_net), .O(n28440));   // verilog/coms.v(127[12] 300[6])
    defparam i14926_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2693_19 (.CI(n38233), .I0(n2_adj_5255), .I1(n1653), .CO(n38234));
    SB_LUT4 add_2693_18_lut (.I0(n48088), .I1(n2_adj_5255), .I2(n1752), 
            .I3(n38232), .O(encoder0_position_scaled_23__N_51[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_18 (.CI(n38232), .I0(n2_adj_5255), .I1(n1752), .CO(n38233));
    SB_LUT4 add_2693_17_lut (.I0(n48064), .I1(n2_adj_5255), .I2(n1851), 
            .I3(n38231), .O(encoder0_position_scaled_23__N_51[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2693_17 (.CI(n38231), .I0(n2_adj_5255), .I1(n1851), .CO(n38232));
    SB_LUT4 add_2693_16_lut (.I0(n48038), .I1(n2_adj_5255), .I2(n1950), 
            .I3(n38230), .O(encoder0_position_scaled_23__N_51[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_16 (.CI(n38230), .I0(n2_adj_5255), .I1(n1950), .CO(n38231));
    SB_LUT4 add_2693_15_lut (.I0(n48014), .I1(n2_adj_5255), .I2(n2049), 
            .I3(n38229), .O(encoder0_position_scaled_23__N_51[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_15 (.CI(n38229), .I0(n2_adj_5255), .I1(n2049), .CO(n38230));
    SB_LUT4 add_2693_14_lut (.I0(n47917), .I1(n2_adj_5255), .I2(n2148), 
            .I3(n38228), .O(encoder0_position_scaled_23__N_51[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_14 (.CI(n38228), .I0(n2_adj_5255), .I1(n2148), .CO(n38229));
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_19 (.CI(n37516), .I0(GND_net), .I1(n8), 
            .CO(n37517));
    SB_LUT4 add_2693_13_lut (.I0(n47871), .I1(n2_adj_5255), .I2(n2247), 
            .I3(n38227), .O(encoder0_position_scaled_23__N_51[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_13 (.CI(n38227), .I0(n2_adj_5255), .I1(n2247), .CO(n38228));
    SB_LUT4 add_2693_12_lut (.I0(n48548), .I1(n2_adj_5255), .I2(n2346), 
            .I3(n38226), .O(encoder0_position_scaled_23__N_51[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_5188), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n939));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2693_12 (.CI(n38226), .I0(n2_adj_5255), .I1(n2346), .CO(n38227));
    SB_LUT4 add_2693_11_lut (.I0(n48513), .I1(n2_adj_5255), .I2(n2445), 
            .I3(n38225), .O(encoder0_position_scaled_23__N_51[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_11 (.CI(n38225), .I0(n2_adj_5255), .I1(n2445), .CO(n38226));
    SB_LUT4 add_2693_10_lut (.I0(n48486), .I1(n2_adj_5255), .I2(n2544), 
            .I3(n38224), .O(encoder0_position_scaled_23__N_51[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_10 (.CI(n38224), .I0(n2_adj_5255), .I1(n2544), .CO(n38225));
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_9_lut (.I0(n48457), .I1(n2_adj_5255), .I2(n2643), 
            .I3(n38223), .O(encoder0_position_scaled_23__N_51[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_9 (.CI(n38223), .I0(n2_adj_5255), .I1(n2643), .CO(n38224));
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_8_lut (.I0(n48428), .I1(n2_adj_5255), .I2(n2742), 
            .I3(n38222), .O(encoder0_position_scaled_23__N_51[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_8 (.CI(n38222), .I0(n2_adj_5255), .I1(n2742), .CO(n38223));
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2693_7_lut (.I0(n48395), .I1(n2_adj_5255), .I2(n2841), 
            .I3(n38221), .O(encoder0_position_scaled_23__N_51[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_7 (.CI(n38221), .I0(n2_adj_5255), .I1(n2841), .CO(n38222));
    SB_LUT4 add_2693_6_lut (.I0(n48364), .I1(n2_adj_5255), .I2(n2940), 
            .I3(n38220), .O(encoder0_position_scaled_23__N_51[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_6 (.CI(n38220), .I0(n2_adj_5255), .I1(n2940), .CO(n38221));
    SB_LUT4 add_2693_5_lut (.I0(n48333), .I1(n2_adj_5255), .I2(n3039), 
            .I3(n38219), .O(encoder0_position_scaled_23__N_51[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_5 (.CI(n38219), .I0(n2_adj_5255), .I1(n3039), .CO(n38220));
    SB_LUT4 add_2693_4_lut (.I0(n48300), .I1(n2_adj_5255), .I2(n3138), 
            .I3(n38218), .O(encoder0_position_scaled_23__N_51[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_4 (.CI(n38218), .I0(n2_adj_5255), .I1(n3138), .CO(n38219));
    SB_LUT4 add_2693_3_lut (.I0(n48262), .I1(n2_adj_5255), .I2(n3237), 
            .I3(n38217), .O(encoder0_position_scaled_23__N_51[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15229_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n42285), 
            .I3(GND_net), .O(n28743));   // verilog/coms.v(127[12] 300[6])
    defparam i15229_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2693_3 (.CI(n38217), .I0(n2_adj_5255), .I1(n3237), .CO(n38218));
    SB_LUT4 add_2693_2_lut (.I0(n48229), .I1(n2_adj_5255), .I2(n34196), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_51[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2693_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2693_2 (.CI(VCC_net), .I0(n2_adj_5255), .I1(n34196), 
            .CO(n38217));
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(GND_net), .I1(n3204), 
            .I2(VCC_net), .I3(n38216), .O(n3271)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n38215), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n38215), .I0(n3205), 
            .I1(VCC_net), .CO(n38216));
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n38214), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n38214), .I0(n3206), 
            .I1(VCC_net), .CO(n38215));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n38213), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n38213), .I0(n3207), 
            .I1(VCC_net), .CO(n38214));
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n38212), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n38212), .I0(n3208), 
            .I1(VCC_net), .CO(n38213));
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n38211), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n38211), .I0(n3209), 
            .I1(VCC_net), .CO(n38212));
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n38210), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n38210), .I0(n3210), 
            .I1(VCC_net), .CO(n38211));
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n38209), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n38209), .I0(n3211), 
            .I1(VCC_net), .CO(n38210));
    SB_LUT4 i15230_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n42285), 
            .I3(GND_net), .O(n28744));   // verilog/coms.v(127[12] 300[6])
    defparam i15230_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n38208), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n38208), .I0(n3212), 
            .I1(VCC_net), .CO(n38209));
    SB_LUT4 i14788_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n23622), .I3(GND_net), .O(n28302));   // verilog/coms.v(127[12] 300[6])
    defparam i14788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n38207), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n38207), .I0(n3213), 
            .I1(VCC_net), .CO(n38208));
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n38206), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n38206), .I0(n3214), 
            .I1(VCC_net), .CO(n38207));
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n38205), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n38205), .I0(n3215), 
            .I1(VCC_net), .CO(n38206));
    SB_LUT4 i15231_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n42285), 
            .I3(GND_net), .O(n28745));   // verilog/coms.v(127[12] 300[6])
    defparam i15231_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n38204), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n38204), .I0(n3216), 
            .I1(VCC_net), .CO(n38205));
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n38203), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n38203), .I0(n3217), 
            .I1(VCC_net), .CO(n38204));
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n38202), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n38202), .I0(n3218), 
            .I1(VCC_net), .CO(n38203));
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n38201), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n38201), .I0(n3219), 
            .I1(VCC_net), .CO(n38202));
    SB_LUT4 i14927_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n23622), .I3(GND_net), .O(n28441));   // verilog/coms.v(127[12] 300[6])
    defparam i14927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n38200), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n38200), .I0(n3220), 
            .I1(VCC_net), .CO(n38201));
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n38199), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n38199), .I0(n3221), 
            .I1(VCC_net), .CO(n38200));
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n38198), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n38198), .I0(n3222), 
            .I1(VCC_net), .CO(n38199));
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n38197), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n38197), .I0(n3223), 
            .I1(VCC_net), .CO(n38198));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n38196), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n38196), .I0(n3224), 
            .I1(VCC_net), .CO(n38197));
    SB_LUT4 i14928_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n23622), .I3(GND_net), .O(n28442));   // verilog/coms.v(127[12] 300[6])
    defparam i14928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14929_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n23622), .I3(GND_net), .O(n28443));   // verilog/coms.v(127[12] 300[6])
    defparam i14929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n38195), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n38195), .I0(n3225), 
            .I1(VCC_net), .CO(n38196));
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n38194), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n9), 
            .I3(n37515), .O(pwm_setpoint_23__N_191[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n38194), .I0(n3226), 
            .I1(VCC_net), .CO(n38195));
    SB_CARRY unary_minus_10_add_3_18 (.CI(n37515), .I0(GND_net), .I1(n9), 
            .CO(n37516));
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n38193), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c_0));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(CS_CLK_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 add_224_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n37457), .O(encoder1_position_scaled_23__N_75[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n38193), .I0(n3227), 
            .I1(VCC_net), .CO(n38194));
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n38192), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n38192), .I0(n3228), 
            .I1(VCC_net), .CO(n38193));
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n38191), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n38191), .I0(n3229), 
            .I1(GND_net), .CO(n38192));
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n38190), .O(n46883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n38190), .I0(n3230), 
            .I1(GND_net), .CO(n38191));
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n38189), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n38189), .I0(n3231), 
            .I1(VCC_net), .CO(n38190));
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n38188), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n38188), .I0(n3232), 
            .I1(GND_net), .CO(n38189));
    SB_LUT4 i33015_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48147));
    defparam i33015_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14930_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n23622), .I3(GND_net), .O(n28444));   // verilog/coms.v(127[12] 300[6])
    defparam i14930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14931_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n23622), .I3(GND_net), .O(n28445));   // verilog/coms.v(127[12] 300[6])
    defparam i14931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14932_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n23622), .I3(GND_net), .O(n28446));   // verilog/coms.v(127[12] 300[6])
    defparam i14932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14933_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n23622), .I3(GND_net), .O(n28447));   // verilog/coms.v(127[12] 300[6])
    defparam i14933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15232_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n42285), 
            .I3(GND_net), .O(n28746));   // verilog/coms.v(127[12] 300[6])
    defparam i15232_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20552_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n34062));
    defparam i20552_3_lut.LUT_INIT = 16'hc8c8;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n38187), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14688_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28202));   // verilog/coms.v(127[12] 300[6])
    defparam i14688_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n38187), .I0(n3233), 
            .I1(VCC_net), .CO(n38188));
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n38186), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n38186), .I0(n957), 
            .I1(GND_net), .CO(n38187));
    SB_LUT4 i14934_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n23622), .I3(GND_net), .O(n28448));   // verilog/coms.v(127[12] 300[6])
    defparam i14934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14935_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n23622), .I3(GND_net), .O(n28449));   // verilog/coms.v(127[12] 300[6])
    defparam i14935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_224_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n37448), .O(encoder1_position_scaled_23__N_75[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1660 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n45214));
    defparam i1_2_lut_adj_1660.LUT_INIT = 16'heeee;
    SB_LUT4 i14936_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n23622), .I3(GND_net), .O(n28450));   // verilog/coms.v(127[12] 300[6])
    defparam i14936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1661 (.I0(n1429), .I1(n34062), .I2(n1430), .I3(n1431), 
            .O(n43289));
    defparam i1_4_lut_adj_1661.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14689_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n33332), 
            .I3(n26390), .O(n28203));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14689_4_lut.LUT_INIT = 16'hccac;
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n652), 
            .I1(VCC_net), .CO(n38186));
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n48300), .I1(n3105), 
            .I2(VCC_net), .I3(n38185), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14937_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n23622), .I3(GND_net), .O(n28451));   // verilog/coms.v(127[12] 300[6])
    defparam i14937_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_14 (.CI(n37457), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n37458));
    SB_LUT4 i1_4_lut_adj_1662 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n45214), 
            .O(n45220));
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n38184), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n38184), .I0(n3106), 
            .I1(VCC_net), .CO(n38185));
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n38183), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n38183), .I0(n3107), 
            .I1(VCC_net), .CO(n38184));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2), .I3(n37749), .O(displacement_23__N_99[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_5182), .I3(n37748), .O(displacement_23__N_99[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_5 (.CI(n37417), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n37418));
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n38182), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n37748), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_5182), .CO(n37749));
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n38182), .I0(n3108), 
            .I1(VCC_net), .CO(n38183));
    SB_LUT4 i33018_4_lut (.I0(n1423), .I1(n1422), .I2(n45220), .I3(n43289), 
            .O(n1455));
    defparam i33018_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_10_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n10), 
            .I3(n37514), .O(pwm_setpoint_23__N_191[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n38181), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_17 (.CI(n37514), .I0(GND_net), .I1(n10), 
            .CO(n37515));
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n38181), .I0(n3109), 
            .I1(VCC_net), .CO(n38182));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_5181), .I3(n37747), .O(displacement_23__N_99[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n11), 
            .I3(n37513), .O(pwm_setpoint_23__N_191[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n38180), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n38180), .I0(n3110), 
            .I1(VCC_net), .CO(n38181));
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n38179), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n38179), .I0(n3111), 
            .I1(VCC_net), .CO(n38180));
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n38178), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n38178), .I0(n3112), 
            .I1(VCC_net), .CO(n38179));
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n38177), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n38177), .I0(n3113), 
            .I1(VCC_net), .CO(n38178));
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n38176), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n38176), .I0(n3114), 
            .I1(VCC_net), .CO(n38177));
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n38175), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n38175), .I0(n3115), 
            .I1(VCC_net), .CO(n38176));
    SB_LUT4 i14938_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n23622), .I3(GND_net), .O(n28452));   // verilog/coms.v(127[12] 300[6])
    defparam i14938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14939_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n23622), .I3(GND_net), .O(n28453));   // verilog/coms.v(127[12] 300[6])
    defparam i14939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n38174), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14940_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n23622), .I3(GND_net), .O(n28454));   // verilog/coms.v(127[12] 300[6])
    defparam i14940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14941_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n23622), .I3(GND_net), .O(n28455));   // verilog/coms.v(127[12] 300[6])
    defparam i14941_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n37747), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_5181), .CO(n37748));
    SB_LUT4 add_224_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n37456), .O(encoder1_position_scaled_23__N_75[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14690_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28204));   // verilog/coms.v(127[12] 300[6])
    defparam i14690_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n38174), .I0(n3116), 
            .I1(VCC_net), .CO(n38175));
    SB_LUT4 i14691_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28205));   // verilog/coms.v(127[12] 300[6])
    defparam i14691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n38173), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14942_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n23622), .I3(GND_net), .O(n28456));   // verilog/coms.v(127[12] 300[6])
    defparam i14942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_16 (.CI(n37513), .I0(GND_net), .I1(n11), 
            .CO(n37514));
    SB_LUT4 i14943_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n44019), .I3(GND_net), .O(n28457));   // verilog/coms.v(127[12] 300[6])
    defparam i14943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14692_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28206));   // verilog/coms.v(127[12] 300[6])
    defparam i14692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14944_4_lut (.I0(CS_MISO_c), .I1(data_adj_5353[0]), .I2(n11_adj_5197), 
            .I3(state_7__N_4293), .O(n28458));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14944_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n38173), .I0(n3117), 
            .I1(VCC_net), .CO(n38174));
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n38172), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n38172), .I0(n3118), 
            .I1(VCC_net), .CO(n38173));
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n38171), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n38171), .I0(n3119), 
            .I1(VCC_net), .CO(n38172));
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n38170), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n38170), .I0(n3120), 
            .I1(VCC_net), .CO(n38171));
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14693_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28207));   // verilog/coms.v(127[12] 300[6])
    defparam i14693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n38169), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n38169), .I0(n3121), 
            .I1(VCC_net), .CO(n38170));
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n38168), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14694_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28208));   // verilog/coms.v(127[12] 300[6])
    defparam i14694_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n38168), .I0(n3122), 
            .I1(VCC_net), .CO(n38169));
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n38167), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n38167), .I0(n3123), 
            .I1(VCC_net), .CO(n38168));
    SB_CARRY add_224_13 (.CI(n37456), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n37457));
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14695_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n44019), 
            .I3(GND_net), .O(n28209));   // verilog/coms.v(127[12] 300[6])
    defparam i14695_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n38166), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n38166), .I0(n3124), 
            .I1(VCC_net), .CO(n38167));
    SB_LUT4 unary_minus_10_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n12), 
            .I3(n37512), .O(pwm_setpoint_23__N_191[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14696_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n44019), 
            .I3(GND_net), .O(n28210));   // verilog/coms.v(127[12] 300[6])
    defparam i14696_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n38165), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_15 (.CI(n37512), .I0(GND_net), .I1(n12), 
            .CO(n37513));
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n38165), .I0(n3125), 
            .I1(VCC_net), .CO(n38166));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_5180), .I3(n37746), .O(displacement_23__N_99[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n37746), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_5180), .CO(n37747));
    SB_LUT4 i14948_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n23622), 
            .I3(GND_net), .O(n28462));   // verilog/coms.v(127[12] 300[6])
    defparam i14948_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_5 (.CI(n37448), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n37449));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_5179), .I3(n37745), .O(displacement_23__N_99[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n38164), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n38164), .I0(n3126), 
            .I1(VCC_net), .CO(n38165));
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n38163), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n38163), .I0(n3127), 
            .I1(VCC_net), .CO(n38164));
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n38162), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n37745), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_5179), .CO(n37746));
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n38162), .I0(n3128), 
            .I1(VCC_net), .CO(n38163));
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n38161), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_5178), .I3(n37744), .O(displacement_23__N_99[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n38161), .I0(n3129), 
            .I1(GND_net), .CO(n38162));
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n38160), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n38160), .I0(n3130), 
            .I1(GND_net), .CO(n38161));
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14697_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28211));   // verilog/coms.v(127[12] 300[6])
    defparam i14697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n38159), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14949_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n23622), 
            .I3(GND_net), .O(n28463));   // verilog/coms.v(127[12] 300[6])
    defparam i14949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14950_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n23622), 
            .I3(GND_net), .O(n28464));   // verilog/coms.v(127[12] 300[6])
    defparam i14950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13_adj_5189), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n938));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n38159), .I0(n3131), 
            .I1(VCC_net), .CO(n38160));
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n38158), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n37744), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_5178), .CO(n37745));
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n38158), .I0(n3132), 
            .I1(GND_net), .CO(n38159));
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n38157), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_5177), .I3(n37743), .O(displacement_23__N_99[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n38157), .I0(n3133), 
            .I1(VCC_net), .CO(n38158));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n37743), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_5177), .CO(n37744));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_5176), .I3(n37742), .O(displacement_23__N_99[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n37742), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_5176), .CO(n37743));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_5175), .I3(n37741), .O(displacement_23__N_99[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n13), 
            .I3(n37511), .O(pwm_setpoint_23__N_191[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n38157));
    SB_LUT4 i14698_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n44019), 
            .I3(GND_net), .O(n28212));   // verilog/coms.v(127[12] 300[6])
    defparam i14698_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(GND_net), .I1(n3006), 
            .I2(VCC_net), .I3(n38156), .O(n3073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n38155), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n38155), .I0(n3007), 
            .I1(VCC_net), .CO(n38156));
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n38154), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14699_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n44019), 
            .I3(GND_net), .O(n28213));   // verilog/coms.v(127[12] 300[6])
    defparam i14699_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n38154), .I0(n3008), 
            .I1(VCC_net), .CO(n38155));
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n38153), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n38153), .I0(n3009), 
            .I1(VCC_net), .CO(n38154));
    SB_LUT4 i14951_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n23622), 
            .I3(GND_net), .O(n28465));   // verilog/coms.v(127[12] 300[6])
    defparam i14951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n38152), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n38152), .I0(n3010), 
            .I1(VCC_net), .CO(n38153));
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n38151), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n38151), .I0(n3011), 
            .I1(VCC_net), .CO(n38152));
    SB_LUT4 encoder0_position_31__I_0_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n37741), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_5175), .CO(n37742));
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n38150), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n38150), .I0(n3012), 
            .I1(VCC_net), .CO(n38151));
    SB_LUT4 add_224_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n37455), .O(encoder1_position_scaled_23__N_75[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n38149), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n38149), .I0(n3013), 
            .I1(VCC_net), .CO(n38150));
    SB_CARRY add_224_12 (.CI(n37455), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n37456));
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n38148), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_14 (.CI(n37511), .I0(GND_net), .I1(n13), 
            .CO(n37512));
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n38148), .I0(n3014), 
            .I1(VCC_net), .CO(n38149));
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n38147), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n38147), .I0(n3015), 
            .I1(VCC_net), .CO(n38148));
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n38146), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n38146), .I0(n3016), 
            .I1(VCC_net), .CO(n38147));
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n38145), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n38145), .I0(n3017), 
            .I1(VCC_net), .CO(n38146));
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n38144), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n38144), .I0(n3018), 
            .I1(VCC_net), .CO(n38145));
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n38143), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n38143), .I0(n3019), 
            .I1(VCC_net), .CO(n38144));
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n38142), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n38142), .I0(n3020), 
            .I1(VCC_net), .CO(n38143));
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n38141), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n38141), .I0(n3021), 
            .I1(VCC_net), .CO(n38142));
    SB_LUT4 i14700_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n44019), 
            .I3(GND_net), .O(n28214));   // verilog/coms.v(127[12] 300[6])
    defparam i14700_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n38140), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n38140), .I0(n3022), 
            .I1(VCC_net), .CO(n38141));
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n38139), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n38139), .I0(n3023), 
            .I1(VCC_net), .CO(n38140));
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n38138), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14701_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n27617), .I3(GND_net), .O(n28215));   // verilog/coms.v(127[12] 300[6])
    defparam i14701_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_5174), .I3(n37740), .O(displacement_23__N_99[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n38138), .I0(n3024), 
            .I1(VCC_net), .CO(n38139));
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n38137), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n38137), .I0(n3025), 
            .I1(VCC_net), .CO(n38138));
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n38136), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20554_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n34064));
    defparam i20554_3_lut.LUT_INIT = 16'hc8c8;
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n38136), .I0(n3026), 
            .I1(VCC_net), .CO(n38137));
    SB_LUT4 unary_minus_10_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n14_adj_5139), 
            .I3(n37510), .O(pwm_setpoint_23__N_191[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1663 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n45186));
    defparam i1_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i14952_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n23622), 
            .I3(GND_net), .O(n28466));   // verilog/coms.v(127[12] 300[6])
    defparam i14952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n38135), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n38135), .I0(n3027), 
            .I1(VCC_net), .CO(n38136));
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n38134), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n38134), .I0(n3028), 
            .I1(VCC_net), .CO(n38135));
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n38133), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n38133), .I0(n3029), 
            .I1(GND_net), .CO(n38134));
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n38132), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n38132), .I0(n3030), 
            .I1(GND_net), .CO(n38133));
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n38131), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n38131), .I0(n3031), 
            .I1(VCC_net), .CO(n38132));
    SB_LUT4 i14953_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n23622), 
            .I3(GND_net), .O(n28467));   // verilog/coms.v(127[12] 300[6])
    defparam i14953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14954_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n23622), 
            .I3(GND_net), .O(n28468));   // verilog/coms.v(127[12] 300[6])
    defparam i14954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n38130), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n38130), .I0(n3032), 
            .I1(GND_net), .CO(n38131));
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n38129), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n38129), .I0(n3033), 
            .I1(VCC_net), .CO(n38130));
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n38129));
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n7072), 
            .D(n1105), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n48364), .I1(n2907), 
            .I2(VCC_net), .I3(n38128), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14955_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n23622), 
            .I3(GND_net), .O(n28469));   // verilog/coms.v(127[12] 300[6])
    defparam i14955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n38127), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n38127), .I0(n2908), 
            .I1(VCC_net), .CO(n38128));
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n38126), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n38126), .I0(n2909), 
            .I1(VCC_net), .CO(n38127));
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n38125), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n38125), .I0(n2910), 
            .I1(VCC_net), .CO(n38126));
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n38124), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n38124), .I0(n2911), 
            .I1(VCC_net), .CO(n38125));
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n38123), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n38123), .I0(n2912), 
            .I1(VCC_net), .CO(n38124));
    GND i1 (.Y(GND_net));
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n38122), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n38122), .I0(n2913), 
            .I1(VCC_net), .CO(n38123));
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n38121), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n38121), .I0(n2914), 
            .I1(VCC_net), .CO(n38122));
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n38120), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n38120), .I0(n2915), 
            .I1(VCC_net), .CO(n38121));
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n38119), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n38119), .I0(n2916), 
            .I1(VCC_net), .CO(n38120));
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n38118), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n38118), .I0(n2917), 
            .I1(VCC_net), .CO(n38119));
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n38117), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n38117), .I0(n2918), 
            .I1(VCC_net), .CO(n38118));
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n38116), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n38116), .I0(n2919), 
            .I1(VCC_net), .CO(n38117));
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n38115), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n38115), .I0(n2920), 
            .I1(VCC_net), .CO(n38116));
    SB_CARRY unary_minus_10_add_3_13 (.CI(n37510), .I0(GND_net), .I1(n14_adj_5139), 
            .CO(n37511));
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n38114), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n38114), .I0(n2921), 
            .I1(VCC_net), .CO(n38115));
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n38113), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n38113), .I0(n2922), 
            .I1(VCC_net), .CO(n38114));
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n38112), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n38112), .I0(n2923), 
            .I1(VCC_net), .CO(n38113));
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n38111), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n38111), .I0(n2924), 
            .I1(VCC_net), .CO(n38112));
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n38110), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n38110), .I0(n2925), 
            .I1(VCC_net), .CO(n38111));
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n38109), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n38109), .I0(n2926), 
            .I1(VCC_net), .CO(n38110));
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n38108), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n38108), .I0(n2927), 
            .I1(VCC_net), .CO(n38109));
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n7072), 
            .D(n1104), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n38107), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n38107), .I0(n2928), 
            .I1(VCC_net), .CO(n38108));
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n38106), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n38106), .I0(n2929), 
            .I1(GND_net), .CO(n38107));
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n38105), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1664 (.I0(n1329), .I1(n34064), .I2(n1330), .I3(n1331), 
            .O(n43270));
    defparam i1_4_lut_adj_1664.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n38105), .I0(n2930), 
            .I1(GND_net), .CO(n38106));
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n38104), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n38104), .I0(n2931), 
            .I1(VCC_net), .CO(n38105));
    SB_LUT4 unary_minus_10_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_5144));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n37740), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_5174), .CO(n37741));
    SB_LUT4 unary_minus_10_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n15_adj_5140), 
            .I3(n37509), .O(pwm_setpoint_23__N_191[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n38103), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut (.I0(n32652), .I1(n20_adj_5252), .I2(n42251), .I3(n122), 
            .O(n43746));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n38103), .I0(n2932), 
            .I1(GND_net), .CO(n38104));
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33034_4_lut (.I0(n43270), .I1(n1323), .I2(n1324), .I3(n45186), 
            .O(n1356));
    defparam i33034_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n38102), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n38102), .I0(n2933), 
            .I1(VCC_net), .CO(n38103));
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n38102));
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n48395), .I1(n2808), 
            .I2(VCC_net), .I3(n38101), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n38100), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n38100), .I0(n2809), 
            .I1(VCC_net), .CO(n38101));
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n38099), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n38099), .I0(n2810), 
            .I1(VCC_net), .CO(n38100));
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n38098), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i769_3_lut (.I0(n1126), .I1(n1193), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n38098), .I0(n2811), 
            .I1(VCC_net), .CO(n38099));
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n38097), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n38097), .I0(n2812), 
            .I1(VCC_net), .CO(n38098));
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n38096), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n38096), .I0(n2813), 
            .I1(VCC_net), .CO(n38097));
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n38095), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n38095), .I0(n2814), 
            .I1(VCC_net), .CO(n38096));
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n38094), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n38094), .I0(n2815), 
            .I1(VCC_net), .CO(n38095));
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n38093), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut_adj_1665 (.I0(n43746), .I1(\FRAME_MATCHER.state_31__N_2788 [2]), 
            .I2(n7_adj_5248), .I3(n26482), .O(n8_adj_5183));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1665.LUT_INIT = 16'hfafe;
    SB_LUT4 i4_4_lut (.I0(\FRAME_MATCHER.state_31__N_2660 [2]), .I1(n8_adj_5183), 
            .I2(n62), .I3(n42244), .O(n48873));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut.LUT_INIT = 16'hefcf;
    SB_LUT4 i14957_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n44019), .I3(GND_net), .O(n28471));   // verilog/coms.v(127[12] 300[6])
    defparam i14957_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14958_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n44019), .I3(GND_net), .O(n28472));   // verilog/coms.v(127[12] 300[6])
    defparam i14958_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY unary_minus_10_add_3_12 (.CI(n37509), .I0(GND_net), .I1(n15_adj_5140), 
            .CO(n37510));
    SB_LUT4 unary_minus_10_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n16), 
            .I3(n37508), .O(pwm_setpoint_23__N_191[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_11 (.CI(n37508), .I0(GND_net), .I1(n16), 
            .CO(n37509));
    SB_LUT4 add_224_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n37454), .O(encoder1_position_scaled_23__N_75[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n38093), .I0(n2816), 
            .I1(VCC_net), .CO(n38094));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_5173), .I3(n37739), .O(displacement_23__N_99[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n38092), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_11 (.CI(n37454), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n37455));
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n38092), .I0(n2817), 
            .I1(VCC_net), .CO(n38093));
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n38091), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n38091), .I0(n2818), 
            .I1(VCC_net), .CO(n38092));
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14959_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n44019), .I3(GND_net), .O(n28473));   // verilog/coms.v(127[12] 300[6])
    defparam i14959_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n37453), .O(encoder1_position_scaled_23__N_75[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_10 (.CI(n37453), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n37454));
    SB_LUT4 unary_minus_10_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n17_adj_5141), 
            .I3(n37507), .O(pwm_setpoint_23__N_191[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_10 (.CI(n37507), .I0(GND_net), .I1(n17_adj_5141), 
            .CO(n37508));
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n38090), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14960_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n44019), .I3(GND_net), .O(n28474));   // verilog/coms.v(127[12] 300[6])
    defparam i14960_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n38090), .I0(n2819), 
            .I1(VCC_net), .CO(n38091));
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n38089), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14961_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n44019), .I3(GND_net), .O(n28475));   // verilog/coms.v(127[12] 300[6])
    defparam i14961_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14962_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n44019), .I3(GND_net), .O(n28476));   // verilog/coms.v(127[12] 300[6])
    defparam i14962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33325_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48457));
    defparam i33325_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14963_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n44019), .I3(GND_net), .O(n28477));   // verilog/coms.v(127[12] 300[6])
    defparam i14963_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n38089), .I0(n2820), 
            .I1(VCC_net), .CO(n38090));
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195_adj_5238), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n37739), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_5173), .CO(n37740));
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n37452), .O(encoder1_position_scaled_23__N_75[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n38088), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n38088), .I0(n2821), 
            .I1(VCC_net), .CO(n38089));
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n38087), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n38087), .I0(n2822), 
            .I1(VCC_net), .CO(n38088));
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n38086), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n38086), .I0(n2823), 
            .I1(VCC_net), .CO(n38087));
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n38085), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n38085), .I0(n2824), 
            .I1(VCC_net), .CO(n38086));
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n38084), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n38084), .I0(n2825), 
            .I1(VCC_net), .CO(n38085));
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n38083), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n38083), .I0(n2826), 
            .I1(VCC_net), .CO(n38084));
    SB_LUT4 i14964_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n44019), .I3(GND_net), .O(n28478));   // verilog/coms.v(127[12] 300[6])
    defparam i14964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14965_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n44019), .I3(GND_net), .O(n28479));   // verilog/coms.v(127[12] 300[6])
    defparam i14965_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_5202), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n937));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20556_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n34066));
    defparam i20556_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n38082), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1666 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n45202));
    defparam i1_3_lut_adj_1666.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n38082), .I0(n2827), 
            .I1(VCC_net), .CO(n38083));
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n38081), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n38081), .I0(n2828), 
            .I1(VCC_net), .CO(n38082));
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n38080), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n38080), .I0(n2829), 
            .I1(GND_net), .CO(n38081));
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n38079), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n38079), .I0(n2830), 
            .I1(GND_net), .CO(n38080));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_224_9 (.CI(n37452), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n37453));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_5172), .I3(n37738), .O(displacement_23__N_99[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n38078), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n38078), .I0(n2831), 
            .I1(VCC_net), .CO(n38079));
    SB_LUT4 i33201_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48333));
    defparam i33201_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(n1229), .I1(n34066), .I2(n1230), .I3(n1231), 
            .O(n43273));
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'ha080;
    SB_LUT4 i33049_4_lut (.I0(n1225), .I1(n1224), .I2(n43273), .I3(n45202), 
            .O(n1257));
    defparam i33049_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i20514_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n34024));
    defparam i20514_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1668 (.I0(n3021), .I1(n3027), .I2(n3028), .I3(n3023), 
            .O(n45452));
    defparam i1_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093_adj_5229), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098_adj_5234), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14968_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n44019), .I3(GND_net), .O(n28482));   // verilog/coms.v(127[12] 300[6])
    defparam i14968_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097_adj_5233), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096_adj_5232), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14703_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n44019), .I3(GND_net), .O(n28217));   // verilog/coms.v(127[12] 300[6])
    defparam i14703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14969_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n44019), .I3(GND_net), .O(n28483));   // verilog/coms.v(127[12] 300[6])
    defparam i14969_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14973_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n44019), .I3(GND_net), .O(n28487));   // verilog/coms.v(127[12] 300[6])
    defparam i14973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1669 (.I0(n3025), .I1(n3019), .I2(n3024), .I3(GND_net), 
            .O(n45450));
    defparam i1_3_lut_adj_1669.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(n45450), .I1(n45452), .I2(n3020), .I3(n3022), 
            .O(n45456));
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1671 (.I0(n3029), .I1(n34024), .I2(n3030), .I3(n3031), 
            .O(n43421));
    defparam i1_4_lut_adj_1671.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095_adj_5231), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i702_3_lut (.I0(n1027), .I1(n1094_adj_5230), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n38077), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n38077), .I0(n2832), 
            .I1(GND_net), .CO(n38078));
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n38076), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_99[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n38076), .I0(n2833), 
            .I1(VCC_net), .CO(n38077));
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_99[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_i709_3_lut (.I0(n935), .I1(n1101_adj_5237), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100_adj_5236), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14974_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n44019), .I3(GND_net), .O(n28488));   // verilog/coms.v(127[12] 300[6])
    defparam i14974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14975_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n44019), .I3(GND_net), .O(n28489));   // verilog/coms.v(127[12] 300[6])
    defparam i14975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5160));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_99[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_99[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_99[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_99[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_99[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_99[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i1_4_lut_adj_1672 (.I0(n3013), .I1(n3015), .I2(n43421), .I3(n45456), 
            .O(n45462));
    defparam i1_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099_adj_5235), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_5203), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n936));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_99[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_99[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i14976_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n44019), .I3(GND_net), .O(n28490));   // verilog/coms.v(127[12] 300[6])
    defparam i14976_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_99[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_99[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_99[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_99[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_99[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_99[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_99[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_99[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_99[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_99[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_99[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_99[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_99[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i14704_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28218));   // verilog/coms.v(127[12] 300[6])
    defparam i14704_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14977_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n44019), .I3(GND_net), .O(n28491));   // verilog/coms.v(127[12] 300[6])
    defparam i14977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1673 (.I0(n3016), .I1(n3017), .I2(n3018), .I3(n3026), 
            .O(n45476));
    defparam i1_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5161));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14705_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n44019), .I3(GND_net), .O(n28219));   // verilog/coms.v(127[12] 300[6])
    defparam i14705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14978_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n44019), .I3(GND_net), .O(n28492));   // verilog/coms.v(127[12] 300[6])
    defparam i14978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(n3009), .I1(n3011), .I2(n3012), .I3(n45462), 
            .O(n45468));
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i14979_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n44019), .I3(GND_net), .O(n28493));   // verilog/coms.v(127[12] 300[6])
    defparam i14979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1675 (.I0(n3008), .I1(n3010), .I2(n3014), .I3(n45476), 
            .O(n45482));
    defparam i1_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1676 (.I0(n20_adj_5252), .I1(n43068), .I2(n42244), 
            .I3(n43094), .O(n44847));
    defparam i3_4_lut_adj_1676.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_3_lut_adj_1677 (.I0(\FRAME_MATCHER.state [0]), .I1(n44847), 
            .I2(n23516), .I3(GND_net), .O(n17_adj_5254));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_adj_1677.LUT_INIT = 16'h8c8c;
    SB_LUT4 i1_4_lut_adj_1678 (.I0(n6_adj_5159), .I1(n17_adj_5254), .I2(n60), 
            .I3(\FRAME_MATCHER.state [3]), .O(n41665));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1678.LUT_INIT = 16'hcdcc;
    SB_LUT4 i14980_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n44019), .I3(GND_net), .O(n28494));   // verilog/coms.v(127[12] 300[6])
    defparam i14980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33204_4_lut (.I0(n3007), .I1(n45482), .I2(n45468), .I3(n3006), 
            .O(n3039));
    defparam i33204_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i20619_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n34130));
    defparam i20619_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i14707_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28221));   // verilog/coms.v(127[12] 300[6])
    defparam i14707_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i14981_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n44019), .I3(GND_net), .O(n28495));   // verilog/coms.v(127[12] 300[6])
    defparam i14981_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_75[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_75[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_LUT4 i1_3_lut_adj_1679 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n45178));
    defparam i1_3_lut_adj_1679.LUT_INIT = 16'hfefe;
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n38076));
    SB_LUT4 i14708_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n44019), 
            .I3(GND_net), .O(n28222));   // verilog/coms.v(127[12] 300[6])
    defparam i14708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14709_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n44019), 
            .I3(GND_net), .O(n28223));   // verilog/coms.v(127[12] 300[6])
    defparam i14709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14982_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n44019), .I3(GND_net), .O(n28496));   // verilog/coms.v(127[12] 300[6])
    defparam i14982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14710_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n44019), 
            .I3(GND_net), .O(n28224));   // verilog/coms.v(127[12] 300[6])
    defparam i14710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(n48428), .I1(n2709), 
            .I2(VCC_net), .I3(n38075), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n38074), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n37738), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_5172), .CO(n37739));
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n38074), .I0(n2710), 
            .I1(VCC_net), .CO(n38075));
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n38073), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n38073), .I0(n2711), 
            .I1(VCC_net), .CO(n38074));
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n38072), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n38072), .I0(n2712), 
            .I1(VCC_net), .CO(n38073));
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n38071), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n38071), .I0(n2713), 
            .I1(VCC_net), .CO(n38072));
    SB_LUT4 add_145_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n37424), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n38070), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n38070), .I0(n2714), 
            .I1(VCC_net), .CO(n38071));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_5171), .I3(n37737), .O(displacement_23__N_99[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n38069), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n38069), .I0(n2715), 
            .I1(VCC_net), .CO(n38070));
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n38068), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n38068), .I0(n2716), 
            .I1(VCC_net), .CO(n38069));
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n38067), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n37737), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_5171), .CO(n37738));
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n38067), .I0(n2717), 
            .I1(VCC_net), .CO(n38068));
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n38066), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n38066), .I0(n2718), 
            .I1(VCC_net), .CO(n38067));
    SB_LUT4 i14983_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n44019), .I3(GND_net), .O(n28497));   // verilog/coms.v(127[12] 300[6])
    defparam i14983_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n38065), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_5170), .I3(n37736), .O(displacement_23__N_99[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n38065), .I0(n2719), 
            .I1(VCC_net), .CO(n38066));
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n38064), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n38064), .I0(n2720), 
            .I1(VCC_net), .CO(n38065));
    SB_LUT4 unary_minus_10_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n18_adj_5142), 
            .I3(n37506), .O(pwm_setpoint_23__N_191[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n38063), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n38063), .I0(n2721), 
            .I1(VCC_net), .CO(n38064));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n37736), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_5170), .CO(n37737));
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n38062), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_5169), .I3(n37735), .O(displacement_23__N_99[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n37735), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_5169), .CO(n37736));
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n38062), .I0(n2722), 
            .I1(VCC_net), .CO(n38063));
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n38061), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n38061), .I0(n2723), 
            .I1(VCC_net), .CO(n38062));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_5168), .I3(n37734), .O(displacement_23__N_99[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n37734), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_5168), .CO(n37735));
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n38060), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n38060), .I0(n2724), 
            .I1(VCC_net), .CO(n38061));
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n38059), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n38059), .I0(n2725), 
            .I1(VCC_net), .CO(n38060));
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n38058), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n38058), .I0(n2726), 
            .I1(VCC_net), .CO(n38059));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_5167), .I3(n37733), .O(displacement_23__N_99[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n38057), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n38057), .I0(n2727), 
            .I1(VCC_net), .CO(n38058));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n38056), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n37447), .O(encoder1_position_scaled_23__N_75[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n38056), .I0(n2728), 
            .I1(VCC_net), .CO(n38057));
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n38055), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n38055), .I0(n2729), 
            .I1(GND_net), .CO(n38056));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n37733), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_5167), .CO(n37734));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_5166), .I3(n37732), .O(displacement_23__N_99[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n37732), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_5166), .CO(n37733));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_5165), .I3(n37731), .O(displacement_23__N_99[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n37731), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_5165), .CO(n37732));
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n28486));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY unary_minus_10_add_3_9 (.CI(n37506), .I0(GND_net), .I1(n18_adj_5142), 
            .CO(n37507));
    SB_DFF commutation_state_i1 (.Q(commutation_state[1]), .C(CLK_c), .D(n42087));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i14711_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n44019), 
            .I3(GND_net), .O(n28225));   // verilog/coms.v(127[12] 300[6])
    defparam i14711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_5164), .I3(n37730), .O(displacement_23__N_99[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n37730), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_5164), .CO(n37731));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_5163), .I3(n37729), .O(displacement_23__N_99[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14984_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n44019), .I3(GND_net), .O(n28498));   // verilog/coms.v(127[12] 300[6])
    defparam i14984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n19_adj_5143), 
            .I3(n37505), .O(pwm_setpoint_23__N_191[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n37729), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_5163), .CO(n37730));
    SB_LUT4 i14712_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n44019), 
            .I3(GND_net), .O(n28226));   // verilog/coms.v(127[12] 300[6])
    defparam i14712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_5162), .I3(n37728), .O(displacement_23__N_99[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n37728), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_5162), .CO(n37729));
    SB_LUT4 add_145_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n37416), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n38054), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14985_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n44019), .I3(GND_net), .O(n28499));   // verilog/coms.v(127[12] 300[6])
    defparam i14985_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n38054), .I0(n2730), 
            .I1(GND_net), .CO(n38055));
    SB_CARRY add_145_12 (.CI(n37424), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n37425));
    SB_LUT4 i14986_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n44019), .I3(GND_net), .O(n28500));   // verilog/coms.v(127[12] 300[6])
    defparam i14986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n38053), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14713_3_lut (.I0(current[0]), .I1(data_adj_5353[0]), .I2(n43722), 
            .I3(GND_net), .O(n28227));   // verilog/tli4970.v(33[10] 66[6])
    defparam i14713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(enable_slow_N_4190), .I1(data_ready), 
            .I2(state_adj_5349[1]), .I3(state_adj_5349[0]), .O(n41973));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'hccd0;
    SB_LUT4 i1_2_lut_adj_1681 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n45198));
    defparam i1_2_lut_adj_1681.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14987_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n44019), .I3(GND_net), .O(n28501));   // verilog/coms.v(127[12] 300[6])
    defparam i14987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33063_4_lut (.I0(n45198), .I1(n1125), .I2(n45178), .I3(n34130), 
            .O(n1158));
    defparam i33063_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 i14715_4_lut (.I0(rw), .I1(state_adj_5349[0]), .I2(state_adj_5349[1]), 
            .I3(n5615), .O(n28229));   // verilog/eeprom.v(26[8] 58[4])
    defparam i14715_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i14991_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n44019), .I3(GND_net), .O(n28505));   // verilog/coms.v(127[12] 300[6])
    defparam i14991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_5161), .I3(n37727), .O(displacement_23__N_99[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14718_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28232));   // verilog/coms.v(127[12] 300[6])
    defparam i14718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14719_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n44019), 
            .I3(GND_net), .O(n28233));   // verilog/coms.v(127[12] 300[6])
    defparam i14719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14992_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n44019), .I3(GND_net), .O(n28506));   // verilog/coms.v(127[12] 300[6])
    defparam i14992_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n38053), .I0(n2731), 
            .I1(VCC_net), .CO(n38054));
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n38052), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n38052), .I0(n2732), 
            .I1(GND_net), .CO(n38053));
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n38051), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n38051), .I0(n2733), 
            .I1(VCC_net), .CO(n38052));
    SB_LUT4 i14993_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n44019), .I3(GND_net), .O(n28507));   // verilog/coms.v(127[12] 300[6])
    defparam i14993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n38051));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n37727), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_5161), .CO(n37728));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_5160), .I3(VCC_net), .O(displacement_23__N_99[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_5160), .CO(n37727));
    SB_LUT4 i14720_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n44019), 
            .I3(GND_net), .O(n28234));   // verilog/coms.v(127[12] 300[6])
    defparam i14720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14994_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n44019), .I3(GND_net), .O(n28508));   // verilog/coms.v(127[12] 300[6])
    defparam i14994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(n48457), .I1(n2610), 
            .I2(VCC_net), .I3(n38050), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n38049), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n38049), .I0(n2611), 
            .I1(VCC_net), .CO(n38050));
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n38048), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_DFF dti_counter_2188__i0 (.Q(dti_counter[0]), .C(CLK_c), .D(n55));   // verilog/TinyFPGA_B.v(159[23:37])
    SB_CARRY add_224_4 (.CI(n37447), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n37448));
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n38048), .I0(n2612), 
            .I1(VCC_net), .CO(n38049));
    SB_LUT4 i14995_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n44019), .I3(GND_net), .O(n28509));   // verilog/coms.v(127[12] 300[6])
    defparam i14995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n37446), .O(encoder1_position_scaled_23__N_75[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_8 (.CI(n37505), .I0(GND_net), .I1(n19_adj_5143), 
            .CO(n37506));
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n38047), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n20_adj_5144), 
            .I3(n37504), .O(pwm_setpoint_23__N_191[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_7 (.CI(n37504), .I0(GND_net), .I1(n20_adj_5144), 
            .CO(n37505));
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n38047), .I0(n2613), 
            .I1(VCC_net), .CO(n38048));
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n38046), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14996_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n44019), .I3(GND_net), .O(n28510));   // verilog/coms.v(127[12] 300[6])
    defparam i14996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15000_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n44019), .I3(GND_net), .O(n28514));   // verilog/coms.v(127[12] 300[6])
    defparam i15000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14721_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5364[1]), .I2(n18934), 
            .I3(n4_adj_5153), .O(n28235));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14721_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i15001_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n44019), .I3(GND_net), .O(n28515));   // verilog/coms.v(127[12] 300[6])
    defparam i15001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14722_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28236));   // verilog/coms.v(127[12] 300[6])
    defparam i14722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14723_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28237));   // verilog/coms.v(127[12] 300[6])
    defparam i14723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33073_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48205));
    defparam i33073_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20560_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n34070));
    defparam i20560_3_lut.LUT_INIT = 16'hc8c8;
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[23]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[22]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[21]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[20]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[19]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[18]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[17]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[16]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[15]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[14]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[13]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[12]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[11]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_51[10]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[9]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[8]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[7]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[6]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[5]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[4]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[3]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[2]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_51[1]));   // verilog/TinyFPGA_B.v(319[10] 323[6])
    SB_DFF commutation_state_prev_i2 (.Q(commutation_state_prev[2]), .C(CLK_c), 
           .D(commutation_state[2]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i15002_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n44019), .I3(GND_net), .O(n28516));   // verilog/coms.v(127[12] 300[6])
    defparam i15002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14724_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28238));   // verilog/coms.v(127[12] 300[6])
    defparam i14724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14725_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28239));   // verilog/coms.v(127[12] 300[6])
    defparam i14725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15003_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n44019), .I3(GND_net), .O(n28517));   // verilog/coms.v(127[12] 300[6])
    defparam i15003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14726_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n23622), .I3(GND_net), .O(n28240));   // verilog/coms.v(127[12] 300[6])
    defparam i14726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14727_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28241));   // verilog/coms.v(127[12] 300[6])
    defparam i14727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14728_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n23622), .I3(GND_net), .O(n28242));   // verilog/coms.v(127[12] 300[6])
    defparam i14728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14729_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n44019), 
            .I3(GND_net), .O(n28243));   // verilog/coms.v(127[12] 300[6])
    defparam i14729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15004_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n44019), .I3(GND_net), .O(n28518));   // verilog/coms.v(127[12] 300[6])
    defparam i15004_3_lut.LUT_INIT = 16'hacac;
    SB_DFF commutation_state_prev_i1 (.Q(commutation_state_prev[1]), .C(CLK_c), 
           .D(commutation_state[1]));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n38046), .I0(n2614), 
            .I1(VCC_net), .CO(n38047));
    SB_LUT4 i1_4_lut_adj_1682 (.I0(n1029), .I1(n34070), .I2(n1030), .I3(n1031), 
            .O(n43278));
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'ha080;
    SB_LUT4 i33076_4_lut (.I0(n1026), .I1(n43278), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i33076_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n38045), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15005_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n44019), .I3(GND_net), .O(n28519));   // verilog/coms.v(127[12] 300[6])
    defparam i15005_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHC_184 (.Q(GHC), .C(CLK_c), .E(n27644), .D(GHC_N_403), 
            .R(n27973));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i15006_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n44019), .I3(GND_net), .O(n28520));   // verilog/coms.v(127[12] 300[6])
    defparam i15006_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15007_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n44019), .I3(GND_net), .O(n28521));   // verilog/coms.v(127[12] 300[6])
    defparam i15007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15008_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n44019), .I3(GND_net), .O(n28522));   // verilog/coms.v(127[12] 300[6])
    defparam i15008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15009_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n42276), .I3(GND_net), .O(n28523));   // verilog/coms.v(127[12] 300[6])
    defparam i15009_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15010_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n42276), .I3(GND_net), .O(n28524));   // verilog/coms.v(127[12] 300[6])
    defparam i15010_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15011_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n42276), .I3(GND_net), .O(n28525));   // verilog/coms.v(127[12] 300[6])
    defparam i15011_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15012_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n42276), .I3(GND_net), .O(n28526));   // verilog/coms.v(127[12] 300[6])
    defparam i15012_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15013_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n42276), .I3(GND_net), .O(n28527));   // verilog/coms.v(127[12] 300[6])
    defparam i15013_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n38045), .I0(n2615), 
            .I1(VCC_net), .CO(n38046));
    SB_LUT4 i15014_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n42276), .I3(GND_net), .O(n28528));   // verilog/coms.v(127[12] 300[6])
    defparam i15014_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15015_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n42276), .I3(GND_net), .O(n28529));   // verilog/coms.v(127[12] 300[6])
    defparam i15015_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n7072), 
            .D(n1103), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n7072), 
            .D(n1093), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n7072), 
            .D(n1102), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n7072), 
            .D(n1101), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i14730_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n23622), .I3(GND_net), .O(n28244));   // verilog/coms.v(127[12] 300[6])
    defparam i14730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14731_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n23622), .I3(GND_net), .O(n28245));   // verilog/coms.v(127[12] 300[6])
    defparam i14731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14732_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n23622), .I3(GND_net), .O(n28246));   // verilog/coms.v(127[12] 300[6])
    defparam i14732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15016_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n42276), .I3(GND_net), .O(n28530));   // verilog/coms.v(127[12] 300[6])
    defparam i15016_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14733_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n23622), .I3(GND_net), .O(n28247));   // verilog/coms.v(127[12] 300[6])
    defparam i14733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14734_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n23622), .I3(GND_net), .O(n28248));   // verilog/coms.v(127[12] 300[6])
    defparam i14734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5255));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14738_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n23622), .I3(GND_net), .O(n28252));   // verilog/coms.v(127[12] 300[6])
    defparam i14738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14735_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n23622), .I3(GND_net), .O(n28249));   // verilog/coms.v(127[12] 300[6])
    defparam i14735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14736_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n23622), .I3(GND_net), .O(n28250));   // verilog/coms.v(127[12] 300[6])
    defparam i14736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15025_3_lut (.I0(\data_in_frame[19] [7]), .I1(rx_data[7]), 
            .I2(n42277), .I3(GND_net), .O(n28539));   // verilog/coms.v(127[12] 300[6])
    defparam i15025_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15026_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n42277), .I3(GND_net), .O(n28540));   // verilog/coms.v(127[12] 300[6])
    defparam i15026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15027_3_lut (.I0(\data_in_frame[19] [5]), .I1(rx_data[5]), 
            .I2(n42277), .I3(GND_net), .O(n28541));   // verilog/coms.v(127[12] 300[6])
    defparam i15027_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15028_3_lut (.I0(\data_in_frame[19] [4]), .I1(rx_data[4]), 
            .I2(n42277), .I3(GND_net), .O(n28542));   // verilog/coms.v(127[12] 300[6])
    defparam i15028_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15029_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n42277), .I3(GND_net), .O(n28543));   // verilog/coms.v(127[12] 300[6])
    defparam i15029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15030_3_lut (.I0(\data_in_frame[19] [2]), .I1(rx_data[2]), 
            .I2(n42277), .I3(GND_net), .O(n28544));   // verilog/coms.v(127[12] 300[6])
    defparam i15030_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15031_3_lut (.I0(\data_in_frame[19] [1]), .I1(rx_data[1]), 
            .I2(n42277), .I3(GND_net), .O(n28545));   // verilog/coms.v(127[12] 300[6])
    defparam i15031_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5162));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15032_3_lut (.I0(\data_in_frame[19] [0]), .I1(rx_data[0]), 
            .I2(n42277), .I3(GND_net), .O(n28546));   // verilog/coms.v(127[12] 300[6])
    defparam i15032_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n38044), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n38044), .I0(n2616), 
            .I1(VCC_net), .CO(n38045));
    SB_CARRY add_224_3 (.CI(n37446), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n37447));
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n38043), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n38043), .I0(n2617), 
            .I1(VCC_net), .CO(n38044));
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n7072), 
            .D(n1100), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n7072), 
            .D(n1092), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n7072), 
            .D(n1091), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n38042), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n38042), .I0(n2618), 
            .I1(VCC_net), .CO(n38043));
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n38041), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n38041), .I0(n2619), 
            .I1(VCC_net), .CO(n38042));
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n38040), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n38040), .I0(n2620), 
            .I1(VCC_net), .CO(n38041));
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n38039), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n38039), .I0(n2621), 
            .I1(VCC_net), .CO(n38040));
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n38038), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n38038), .I0(n2622), 
            .I1(VCC_net), .CO(n38039));
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n38037), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n38037), .I0(n2623), 
            .I1(VCC_net), .CO(n38038));
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n7072), 
            .D(n1099), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n38036), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n38036), .I0(n2624), 
            .I1(VCC_net), .CO(n38037));
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n38035), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n38035), .I0(n2625), 
            .I1(VCC_net), .CO(n38036));
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n7072), 
            .D(n1090), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n38034), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n7072), 
            .D(n1089), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n38034), .I0(n2626), 
            .I1(VCC_net), .CO(n38035));
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n38033), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n38033), .I0(n2627), 
            .I1(VCC_net), .CO(n38034));
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n38032), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n38032), .I0(n2628), 
            .I1(VCC_net), .CO(n38033));
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n38031), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n38031), .I0(n2629), 
            .I1(GND_net), .CO(n38032));
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n38030), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n38030), .I0(n2630), 
            .I1(GND_net), .CO(n38031));
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n38029), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n38029), .I0(n2631), 
            .I1(VCC_net), .CO(n38030));
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n38028), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n38028), .I0(n2632), 
            .I1(GND_net), .CO(n38029));
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n38027), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n38027), .I0(n2633), 
            .I1(VCC_net), .CO(n38028));
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR pwm_setpoint__i23 (.Q(pwm_setpoint[23]), .C(CLK_c), .D(pwm_setpoint_23__N_191[23]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_23__N_191[22]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_23__N_191[21]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_23__N_191[20]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_23__N_191[19]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_23__N_191[18]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_23__N_191[17]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_23__N_191[16]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_23__N_191[15]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_23__N_191[14]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_23__N_191[13]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFFSR pwm_setpoint__i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_23__N_191[12]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n38027));
    SB_DFFSR pwm_setpoint__i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_23__N_191[11]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_23__N_191[10]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_23__N_191[9]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_23__N_191[8]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_23__N_191[7]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_23__N_191[6]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_23__N_191[5]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_23__N_191[4]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_23__N_191[3]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_23__N_191[2]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_DFFSR pwm_setpoint__i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_23__N_191[1]), 
            .R(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n48486), .I1(n2511), 
            .I2(VCC_net), .I3(n38026), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n38025), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n38025), .I0(n2512), 
            .I1(VCC_net), .CO(n38026));
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n38024), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n38024), .I0(n2513), 
            .I1(VCC_net), .CO(n38025));
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n38023), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n38023), .I0(n2514), 
            .I1(VCC_net), .CO(n38024));
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n38022), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n38022), .I0(n2515), 
            .I1(VCC_net), .CO(n38023));
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n38021), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GHB_182 (.Q(GHB), .C(CLK_c), .E(n27644), .D(GHB_N_389), 
            .R(n27973));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n38021), .I0(n2516), 
            .I1(VCC_net), .CO(n38022));
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n38020), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n38020), .I0(n2517), 
            .I1(VCC_net), .CO(n38021));
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n38019), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n38019), .I0(n2518), 
            .I1(VCC_net), .CO(n38020));
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n38018), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n38018), .I0(n2519), 
            .I1(VCC_net), .CO(n38019));
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n38017), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n38017), .I0(n2520), 
            .I1(VCC_net), .CO(n38018));
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n38016), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n38016), .I0(n2521), 
            .I1(VCC_net), .CO(n38017));
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n38015), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_3_lut (.I0(h1), .I1(h3), .I2(h2), .I3(GND_net), 
            .O(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n38015), .I0(n2522), 
            .I1(VCC_net), .CO(n38016));
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n38014), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n38014), .I0(n2523), 
            .I1(VCC_net), .CO(n38015));
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n38013), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n38013), .I0(n2524), 
            .I1(VCC_net), .CO(n38014));
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15256_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n27617), .I3(GND_net), .O(n28770));   // verilog/coms.v(127[12] 300[6])
    defparam i15256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n38012), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n38012), .I0(n2525), 
            .I1(VCC_net), .CO(n38013));
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n38011), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n38011), .I0(n2526), 
            .I1(VCC_net), .CO(n38012));
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n38010), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n38010), .I0(n2527), 
            .I1(VCC_net), .CO(n38011));
    SB_LUT4 i15257_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n27617), .I3(GND_net), .O(n28771));   // verilog/coms.v(127[12] 300[6])
    defparam i15257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15057_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n42267), .I3(GND_net), .O(n28571));   // verilog/coms.v(127[12] 300[6])
    defparam i15057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15058_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n42267), .I3(GND_net), .O(n28572));   // verilog/coms.v(127[12] 300[6])
    defparam i15058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15258_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n27617), .I3(GND_net), .O(n28772));   // verilog/coms.v(127[12] 300[6])
    defparam i15258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15059_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n42267), .I3(GND_net), .O(n28573));   // verilog/coms.v(127[12] 300[6])
    defparam i15059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15060_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n42267), .I3(GND_net), .O(n28574));   // verilog/coms.v(127[12] 300[6])
    defparam i15060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15061_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n42267), .I3(GND_net), .O(n28575));   // verilog/coms.v(127[12] 300[6])
    defparam i15061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15062_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n42267), .I3(GND_net), .O(n28576));   // verilog/coms.v(127[12] 300[6])
    defparam i15062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5143));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15063_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n42267), .I3(GND_net), .O(n28577));   // verilog/coms.v(127[12] 300[6])
    defparam i15063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15259_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n27617), .I3(GND_net), .O(n28773));   // verilog/coms.v(127[12] 300[6])
    defparam i15259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15260_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n27617), .I3(GND_net), .O(n28774));   // verilog/coms.v(127[12] 300[6])
    defparam i15260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n38009), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n38009), .I0(n2528), 
            .I1(VCC_net), .CO(n38010));
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n38008), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n38008), .I0(n2529), 
            .I1(GND_net), .CO(n38009));
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15064_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n42267), .I3(GND_net), .O(n28578));   // verilog/coms.v(127[12] 300[6])
    defparam i15064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n38007), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_224_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_279), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_75[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14739_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n23622), .I3(GND_net), .O(n28253));   // verilog/coms.v(127[12] 300[6])
    defparam i14739_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n38007), .I0(n2530), 
            .I1(GND_net), .CO(n38008));
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n38006), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_224_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_279), 
            .CO(n37446));
    SB_LUT4 i15065_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28579));   // verilog/coms.v(127[12] 300[6])
    defparam i15065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14740_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n23622), .I3(GND_net), .O(n28254));   // verilog/coms.v(127[12] 300[6])
    defparam i14740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n38006), .I0(n2531), 
            .I1(VCC_net), .CO(n38007));
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n38005), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n38005), .I0(n2532), 
            .I1(GND_net), .CO(n38006));
    SB_LUT4 i15261_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n27617), .I3(GND_net), .O(n28775));   // verilog/coms.v(127[12] 300[6])
    defparam i15261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15066_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28580));   // verilog/coms.v(127[12] 300[6])
    defparam i15066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1922_3_lut (.I0(n2823), .I1(n2890), 
            .I2(n2841), .I3(GND_net), .O(n2922));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n38004), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n38004), .I0(n2533), 
            .I1(VCC_net), .CO(n38005));
    SB_LUT4 i14741_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n23622), .I3(GND_net), .O(n28255));   // verilog/coms.v(127[12] 300[6])
    defparam i14741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15262_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n27617), .I3(GND_net), .O(n28776));   // verilog/coms.v(127[12] 300[6])
    defparam i15262_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n41451));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15067_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28581));   // verilog/coms.v(127[12] 300[6])
    defparam i15067_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n38004));
    SB_LUT4 i15263_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n27617), .I3(GND_net), .O(n28777));   // verilog/coms.v(127[12] 300[6])
    defparam i15263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n48513), .I1(n2412), 
            .I2(VCC_net), .I3(n38003), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n38002), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n38002), .I0(n2413), 
            .I1(VCC_net), .CO(n38003));
    SB_LUT4 i15264_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n27617), .I3(GND_net), .O(n28778));   // verilog/coms.v(127[12] 300[6])
    defparam i15264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5163));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15265_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n27617), .I3(GND_net), .O(n28779));   // verilog/coms.v(127[12] 300[6])
    defparam i15265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5164));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15068_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28582));   // verilog/coms.v(127[12] 300[6])
    defparam i15068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n38001), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15266_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n27617), .I3(GND_net), .O(n28780));   // verilog/coms.v(127[12] 300[6])
    defparam i15266_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n38001), .I0(n2414), 
            .I1(VCC_net), .CO(n38002));
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n38000), .O(n2482)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n38000), .I0(n2415), 
            .I1(VCC_net), .CO(n38001));
    SB_LUT4 encoder0_position_31__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n37999), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15267_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n27617), .I3(GND_net), .O(n28781));   // verilog/coms.v(127[12] 300[6])
    defparam i15267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_145_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n37445), .O(n1077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15069_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28583));   // verilog/coms.v(127[12] 300[6])
    defparam i15069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15268_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n27617), .I3(GND_net), .O(n28782));   // verilog/coms.v(127[12] 300[6])
    defparam i15268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15070_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28584));   // verilog/coms.v(127[12] 300[6])
    defparam i15070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15071_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n42255), .I3(GND_net), .O(n28585));   // verilog/coms.v(127[12] 300[6])
    defparam i15071_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n37999), .I0(n2416), 
            .I1(VCC_net), .CO(n38000));
    SB_LUT4 i15072_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28586));   // verilog/coms.v(127[12] 300[6])
    defparam i15072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n37998), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n37998), .I0(n2417), 
            .I1(VCC_net), .CO(n37999));
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n37997), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n37997), .I0(n2418), 
            .I1(VCC_net), .CO(n37998));
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15269_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n27617), .I3(GND_net), .O(n28783));   // verilog/coms.v(127[12] 300[6])
    defparam i15269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(h3), .I1(commutation_state[1]), .I2(h2), 
            .I3(h1), .O(n42087));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'hd054;
    SB_LUT4 i15073_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n42255), .I3(GND_net), .O(n28587));   // verilog/coms.v(127[12] 300[6])
    defparam i15073_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15074_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n42255), .I3(GND_net), .O(n28588));   // verilog/coms.v(127[12] 300[6])
    defparam i15074_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n37996), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15075_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n44019), .I3(GND_net), .O(n28589));   // verilog/coms.v(127[12] 300[6])
    defparam i15075_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n37996), .I0(n2419), 
            .I1(VCC_net), .CO(n37997));
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n37995), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n37995), .I0(n2420), 
            .I1(VCC_net), .CO(n37996));
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15076_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n44019), .I3(GND_net), .O(n28590));   // verilog/coms.v(127[12] 300[6])
    defparam i15076_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1684 (.I0(state_adj_5349[1]), .I1(read), .I2(n42289), 
            .I3(GND_net), .O(n12_adj_5242));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut_adj_1684.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n33881), .I1(n12_adj_5242), .I2(state_adj_5349[0]), 
            .I3(n42289), .O(n41869));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'h88a8;
    SB_LUT4 i15077_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n44019), .I3(GND_net), .O(n28591));   // verilog/coms.v(127[12] 300[6])
    defparam i15077_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n37994), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n37994), .I0(n2421), 
            .I1(VCC_net), .CO(n37995));
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n37993), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n37993), .I0(n2422), 
            .I1(VCC_net), .CO(n37994));
    SB_LUT4 i15078_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n44019), .I3(GND_net), .O(n28592));   // verilog/coms.v(127[12] 300[6])
    defparam i15078_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15079_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n44019), .I3(GND_net), .O(n28593));   // verilog/coms.v(127[12] 300[6])
    defparam i15079_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR GHA_180 (.Q(GHA), .C(CLK_c), .E(n27644), .D(GHA_N_367), 
            .R(n27973));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 i14742_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n23622), .I3(GND_net), .O(n28256));   // verilog/coms.v(127[12] 300[6])
    defparam i14742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14743_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n23622), .I3(GND_net), .O(n28257));   // verilog/coms.v(127[12] 300[6])
    defparam i14743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n7270), .I1(n4_adj_5216), .I2(data_ready), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n42984));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'heaee;
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n37992), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n37992), .I0(n2423), 
            .I1(VCC_net), .CO(n37993));
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n37991), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n37991), .I0(n2424), 
            .I1(VCC_net), .CO(n37992));
    SB_LUT4 i15080_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n44019), .I3(GND_net), .O(n28594));   // verilog/coms.v(127[12] 300[6])
    defparam i15080_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1687 (.I0(\ID_READOUT_FSM.state [0]), .I1(n33250), 
            .I2(\ID_READOUT_FSM.state [1]), .I3(n42984), .O(n27874));
    defparam i2_4_lut_adj_1687.LUT_INIT = 16'h4c00;
    SB_LUT4 i14972_3_lut (.I0(n27874), .I1(\ID_READOUT_FSM.state [0]), .I2(n7270), 
            .I3(GND_net), .O(n28486));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i14972_3_lut.LUT_INIT = 16'h4646;
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n37990), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n37990), .I0(n2425), 
            .I1(VCC_net), .CO(n37991));
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n37989), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n37989), .I0(n2426), 
            .I1(VCC_net), .CO(n37990));
    SB_LUT4 i15081_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n44019), .I3(GND_net), .O(n28595));   // verilog/coms.v(127[12] 300[6])
    defparam i15081_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14744_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n23622), .I3(GND_net), .O(n28258));   // verilog/coms.v(127[12] 300[6])
    defparam i14744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15082_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n44019), .I3(GND_net), .O(n28596));   // verilog/coms.v(127[12] 300[6])
    defparam i15082_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n37988), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n37988), .I0(n2427), 
            .I1(VCC_net), .CO(n37989));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n37987), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n37987), .I0(n2428), 
            .I1(VCC_net), .CO(n37988));
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14917_3_lut (.I0(n28125), .I1(r_Bit_Index[0]), .I2(n27844), 
            .I3(GND_net), .O(n28431));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14917_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i14873_3_lut (.I0(n28123), .I1(r_Bit_Index_adj_5366[0]), .I2(n27840), 
            .I3(GND_net), .O(n28387));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14873_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i15083_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n44019), .I3(GND_net), .O(n28597));   // verilog/coms.v(127[12] 300[6])
    defparam i15083_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14745_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n23622), .I3(GND_net), .O(n28259));   // verilog/coms.v(127[12] 300[6])
    defparam i14745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5165));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15084_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n44019), .I3(GND_net), .O(n28598));   // verilog/coms.v(127[12] 300[6])
    defparam i15084_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14746_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n23622), .I3(GND_net), .O(n28260));   // verilog/coms.v(127[12] 300[6])
    defparam i14746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5166));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15085_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n44019), .I3(GND_net), .O(n28599));   // verilog/coms.v(127[12] 300[6])
    defparam i15085_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n37986), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n37986), .I0(n2429), 
            .I1(GND_net), .CO(n37987));
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n37985), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n37985), .I0(n2430), 
            .I1(GND_net), .CO(n37986));
    SB_LUT4 i14747_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n23622), .I3(GND_net), .O(n28261));   // verilog/coms.v(127[12] 300[6])
    defparam i14747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15086_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n42255), .I3(GND_net), .O(n28600));   // verilog/coms.v(127[12] 300[6])
    defparam i15086_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14748_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n23622), .I3(GND_net), .O(n28262));   // verilog/coms.v(127[12] 300[6])
    defparam i14748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5273));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(n2924), .I1(n2922), .I2(n2920), .I3(n2928), 
            .O(n44942));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'hfffe;
    SB_LUT4 i14749_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n23622), .I3(GND_net), .O(n28263));   // verilog/coms.v(127[12] 300[6])
    defparam i14749_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n37984), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n37984), .I0(n2431), 
            .I1(VCC_net), .CO(n37985));
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n37983), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n7072), 
            .D(n1098), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 i14750_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n44019), 
            .I3(GND_net), .O(n28264));   // verilog/coms.v(127[12] 300[6])
    defparam i14750_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5167));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15087_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n42255), .I3(GND_net), .O(n28601));   // verilog/coms.v(127[12] 300[6])
    defparam i15087_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1689 (.I0(n2919), .I1(n2921), .I2(n2926), .I3(GND_net), 
            .O(n44944));
    defparam i1_3_lut_adj_1689.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5168));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n44942), .I1(n2927), .I2(n2925), .I3(n2923), 
            .O(n44946));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n37983), .I0(n2432), 
            .I1(GND_net), .CO(n37984));
    SB_LUT4 i15088_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n42255), .I3(GND_net), .O(n28602));   // verilog/coms.v(127[12] 300[6])
    defparam i15088_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20579_4_lut (.I0(n954), .I1(n2931), .I2(n2932), .I3(n2933), 
            .O(n34090));
    defparam i20579_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i15089_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n42255), .I3(GND_net), .O(n28603));   // verilog/coms.v(127[12] 300[6])
    defparam i15089_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n37982), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n37982), .I0(n2433), 
            .I1(VCC_net), .CO(n37983));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5169));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n37982));
    SB_LUT4 i14751_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n44019), 
            .I3(GND_net), .O(n28265));   // verilog/coms.v(127[12] 300[6])
    defparam i14751_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n48548), .I1(n2313), 
            .I2(VCC_net), .I3(n37981), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n37980), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n37980), .I0(n2314), 
            .I1(VCC_net), .CO(n37981));
    SB_LUT4 i4_4_lut_adj_1691 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5150));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i4_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 i15090_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n42255), .I3(GND_net), .O(n28604));   // verilog/coms.v(127[12] 300[6])
    defparam i15090_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_5150), .I2(control_mode[2]), 
            .I3(GND_net), .O(n26429));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15091_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n44824), .I3(GND_net), 
            .O(n28605));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15091_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28091_4_lut (.I0(n7_adj_5250), .I1(state_adj_5349[0]), .I2(n6), 
            .I3(state_adj_5377[0]), .O(n43114));
    defparam i28091_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i15092_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n44824), .I3(GND_net), 
            .O(n28606));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15092_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n37979), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n37979), .I0(n2315), 
            .I1(VCC_net), .CO(n37980));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5274), .I3(n38437), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n37978), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15093_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n44824), .I3(GND_net), 
            .O(n28607));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15093_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n37978), .I0(n2316), 
            .I1(VCC_net), .CO(n37979));
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n37977), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15094_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n44824), .I3(GND_net), 
            .O(n28608));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15094_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n33881), .I1(n42289), .I2(state_adj_5349[0]), 
            .I3(read), .O(n41883));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'h8280;
    SB_LUT4 i15095_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n44824), .I3(GND_net), 
            .O(n28609));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15095_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n37977), .I0(n2317), 
            .I1(VCC_net), .CO(n37978));
    SB_LUT4 unary_minus_10_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_5142));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n37976), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15096_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n44824), .I3(GND_net), 
            .O(n28610));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15096_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14752_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n23622), .I3(GND_net), .O(n28266));   // verilog/coms.v(127[12] 300[6])
    defparam i14752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n44824));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i14753_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n44019), 
            .I3(GND_net), .O(n28267));   // verilog/coms.v(127[12] 300[6])
    defparam i14753_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15097_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n44824), .I3(GND_net), 
            .O(n28611));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i15097_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5170));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n37976), .I0(n2318), 
            .I1(VCC_net), .CO(n37977));
    SB_LUT4 i15098_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n42266), .I3(GND_net), .O(n28612));   // verilog/coms.v(127[12] 300[6])
    defparam i15098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n37975), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15099_3_lut (.I0(h1), .I1(reg_B[2]), .I2(n44732), .I3(GND_net), 
            .O(n28613));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i15099_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n37975), .I0(n2319), 
            .I1(VCC_net), .CO(n37976));
    SB_LUT4 i15100_3_lut (.I0(h2), .I1(reg_B[1]), .I2(n44732), .I3(GND_net), 
            .O(n28614));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i15100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n37974), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1693 (.I0(n26277), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5158));   // verilog/TinyFPGA_B.v(268[5:22])
    defparam i1_2_lut_adj_1693.LUT_INIT = 16'hbbbb;
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n37974), .I0(n2320), 
            .I1(VCC_net), .CO(n37975));
    SB_LUT4 i15101_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n42266), .I3(GND_net), .O(n28615));   // verilog/coms.v(127[12] 300[6])
    defparam i15101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15102_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n42266), .I3(GND_net), .O(n28616));   // verilog/coms.v(127[12] 300[6])
    defparam i15102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15103_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n42266), .I3(GND_net), .O(n28617));   // verilog/coms.v(127[12] 300[6])
    defparam i15103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1694 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n26429), .I3(GND_net), .O(n15_adj_5191));   // verilog/TinyFPGA_B.v(267[5:22])
    defparam i2_3_lut_adj_1694.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n2917), .I1(n2918), .I2(n44946), .I3(n44944), 
            .O(n44952));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 i15104_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n42266), .I3(GND_net), .O(n28618));   // verilog/coms.v(127[12] 300[6])
    defparam i15104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[19]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15105_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n41203), .I3(GND_net), .O(n28619));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15106_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n41203), .I3(GND_net), .O(n28620));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31923_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[0]), .O(n46878));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31923_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i15107_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n41203), .I3(GND_net), .O(n28621));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31931_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[1]), .O(n46841));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31931_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n37973), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n37973), .I0(n2321), 
            .I1(VCC_net), .CO(n37974));
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n37972), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n37972), .I0(n2322), 
            .I1(VCC_net), .CO(n37973));
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n37971), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n37971), .I0(n2323), 
            .I1(VCC_net), .CO(n37972));
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n37970), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15108_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n41203), .I3(GND_net), .O(n28622));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5171));   // verilog/TinyFPGA_B.v(322[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15109_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n41203), .I3(GND_net), .O(n28623));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14754_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n44019), 
            .I3(GND_net), .O(n28268));   // verilog/coms.v(127[12] 300[6])
    defparam i14754_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31930_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[2]), .O(n46840));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31930_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 i31929_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[3]), .O(n46839));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31929_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n37970), .I0(n2324), 
            .I1(VCC_net), .CO(n37971));
    SB_LUT4 i15110_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n41203), .I3(GND_net), .O(n28624));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1696 (.I0(n2929), .I1(n2930), .I2(GND_net), .I3(GND_net), 
            .O(n45484));
    defparam i1_2_lut_adj_1696.LUT_INIT = 16'h8888;
    SB_LUT4 i31928_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[4]), .O(n46838));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31928_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n37969), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14755_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n44019), 
            .I3(GND_net), .O(n28269));   // verilog/coms.v(127[12] 300[6])
    defparam i14755_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n37969), .I0(n2325), 
            .I1(VCC_net), .CO(n37970));
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n37968), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(n45484), .I1(n2916), .I2(n44952), .I3(n34090), 
            .O(n44956));
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'hfefc;
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n37968), .I0(n2326), 
            .I1(VCC_net), .CO(n37969));
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n37967), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n37967), .I0(n2327), 
            .I1(VCC_net), .CO(n37968));
    SB_LUT4 i33296_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n48428));
    defparam i33296_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n37966), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15111_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n41203), .I3(GND_net), .O(n28625));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15111_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n37966), .I0(n2328), 
            .I1(VCC_net), .CO(n37967));
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n37965), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n37965), .I0(n2329), 
            .I1(GND_net), .CO(n37966));
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n2913), .I1(n2914), .I2(n2915), .I3(n44956), 
            .O(n44962));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 i15112_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n41203), .I3(GND_net), .O(n28626));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n37964), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15113_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n41203), .I3(GND_net), .O(n28627));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31927_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[5]), .O(n46837));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31927_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n37964), .I0(n2330), 
            .I1(GND_net), .CO(n37965));
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n37963), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31893_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[6]), .O(n46836));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31893_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n37963), .I0(n2331), 
            .I1(VCC_net), .CO(n37964));
    SB_LUT4 mux_238_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[0]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14737_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n23622), .I3(GND_net), .O(n28251));   // verilog/coms.v(127[12] 300[6])
    defparam i14737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n37962), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15114_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n41203), .I3(GND_net), .O(n28628));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31868_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_counter[7]), .O(n46835));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i31868_2_lut_4_lut.LUT_INIT = 16'h2100;
    SB_LUT4 add_145_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n37444), .O(n1078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut (.I0(commutation_state[0]), .I1(n4_adj_5247), 
            .I2(commutation_state_prev[0]), .I3(dti_N_416), .O(n27620));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 i15115_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n41203), .I3(GND_net), .O(n28629));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15116_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n41203), .I3(GND_net), .O(n28630));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15116_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n37962), .I0(n2332), 
            .I1(GND_net), .CO(n37963));
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n2910), .I1(n2911), .I2(n2912), .I3(n44962), 
            .O(n44968));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 i14756_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n44019), 
            .I3(GND_net), .O(n28270));   // verilog/coms.v(127[12] 300[6])
    defparam i14756_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n37961), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15117_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n41203), .I3(GND_net), .O(n28631));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14775_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n23622), .I3(GND_net), .O(n28289));   // verilog/coms.v(127[12] 300[6])
    defparam i14775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15118_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n41203), .I3(GND_net), .O(n28632));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15119_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n41203), .I3(GND_net), .O(n28633));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15120_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n41203), .I3(GND_net), .O(n28634));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15121_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n41203), .I3(GND_net), .O(n28635));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15121_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n37961), .I0(n2333), 
            .I1(VCC_net), .CO(n37962));
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n37961));
    SB_LUT4 i1_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26285), .I3(GND_net), .O(n7072));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i19753_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26285), .I3(n1195), .O(n33250));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i19753_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfbb;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26285), .I3(n1195), .O(n7270));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i15122_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n41203), .I3(GND_net), .O(n28636));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33236_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n44968), 
            .O(n2940));
    defparam i33236_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i15123_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n41203), .I3(GND_net), .O(n28637));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5269));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14776_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n23622), .I3(GND_net), .O(n28290));   // verilog/coms.v(127[12] 300[6])
    defparam i14776_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15124_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n41203), .I3(GND_net), .O(n28638));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19783_2_lut (.I0(n23805), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n33280));
    defparam i19783_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15125_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n41203), .I3(GND_net), .O(n28639));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[1]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26285), .I3(GND_net), .O(n26286));   // verilog/TinyFPGA_B.v(375[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i15126_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n41203), .I3(GND_net), .O(n28640));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15127_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n41203), .I3(GND_net), .O(n28641));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15128_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n41203), .I3(GND_net), .O(n28642));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15129_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n41203), .I3(GND_net), .O(n28643));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15130_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n41203), .I3(GND_net), .O(n28644));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15131_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n41203), .I3(GND_net), .O(n28645));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15132_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n41203), .I3(GND_net), .O(n28646));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[2]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15133_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n41203), .I3(GND_net), .O(n28647));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15134_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n41203), .I3(GND_net), .O(n28648));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1855_3_lut (.I0(n2724), .I1(n2791), 
            .I2(n2742), .I3(GND_net), .O(n2823));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1855_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15135_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n41203), .I3(GND_net), .O(n28649));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15136_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n42266), .I3(GND_net), .O(n28650));   // verilog/coms.v(127[12] 300[6])
    defparam i15136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(n47871), .I1(n2214), 
            .I2(VCC_net), .I3(n37960), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n37959), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n37423), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n21_adj_5145), 
            .I3(n37503), .O(pwm_setpoint_23__N_191[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_6 (.CI(n37503), .I0(GND_net), .I1(n21_adj_5145), 
            .CO(n37504));
    SB_LUT4 unary_minus_10_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n22_adj_5146), 
            .I3(n37502), .O(pwm_setpoint_23__N_191[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n37959), .I0(n2215), 
            .I1(VCC_net), .CO(n37960));
    SB_LUT4 mux_238_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[3]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n37958), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n37958), .I0(n2216), 
            .I1(VCC_net), .CO(n37959));
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n37957), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n37957), .I0(n2217), 
            .I1(VCC_net), .CO(n37958));
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n37956), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n37956), .I0(n2218), 
            .I1(VCC_net), .CO(n37957));
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n37955), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n37955), .I0(n2219), 
            .I1(VCC_net), .CO(n37956));
    SB_CARRY unary_minus_10_add_3_5 (.CI(n37502), .I0(GND_net), .I1(n22_adj_5146), 
            .CO(n37503));
    SB_LUT4 unary_minus_10_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n23_adj_5147), 
            .I3(n37501), .O(pwm_setpoint_23__N_191[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_32 (.CI(n37444), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n37445));
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n37954), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_4 (.CI(n37501), .I0(GND_net), .I1(n23_adj_5147), 
            .CO(n37502));
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n37954), .I0(n2220), 
            .I1(VCC_net), .CO(n37955));
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n37953), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n37953), .I0(n2221), 
            .I1(VCC_net), .CO(n37954));
    SB_LUT4 add_145_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n37443), .O(n1079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n37952), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n37952), .I0(n2222), 
            .I1(VCC_net), .CO(n37953));
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n37951), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_31 (.CI(n37443), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n37444));
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n37951), .I0(n2223), 
            .I1(VCC_net), .CO(n37952));
    SB_LUT4 unary_minus_10_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n24_adj_5148), 
            .I3(n37500), .O(pwm_setpoint_23__N_191[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n37950), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n37950), .I0(n2224), 
            .I1(VCC_net), .CO(n37951));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n37949), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n37949), .I0(n2225), 
            .I1(VCC_net), .CO(n37950));
    SB_CARRY add_145_4 (.CI(n37416), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n37417));
    SB_CARRY add_145_11 (.CI(n37423), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n37424));
    SB_CARRY unary_minus_10_add_3_3 (.CI(n37500), .I0(GND_net), .I1(n24_adj_5148), 
            .CO(n37501));
    SB_LUT4 unary_minus_10_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n25_adj_5149), 
            .I3(VCC_net), .O(pwm_setpoint_23__N_191[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_10_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_10_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_5149), 
            .CO(n37500));
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n37948), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n37948), .I0(n2226), 
            .I1(VCC_net), .CO(n37949));
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n37947), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n37947), .I0(n2227), 
            .I1(VCC_net), .CO(n37948));
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n37946), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n37946), .I0(n2228), 
            .I1(VCC_net), .CO(n37947));
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n37945), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n37945), .I0(n2229), 
            .I1(GND_net), .CO(n37946));
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n37944), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n37944), .I0(n2230), 
            .I1(GND_net), .CO(n37945));
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n37943), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n37943), .I0(n2231), 
            .I1(VCC_net), .CO(n37944));
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15137_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n42266), .I3(GND_net), .O(n28651));   // verilog/coms.v(127[12] 300[6])
    defparam i15137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15138_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n42266), .I3(GND_net), .O(n28652));   // verilog/coms.v(127[12] 300[6])
    defparam i15138_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n37942), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n37942), .I0(n2232), 
            .I1(GND_net), .CO(n37943));
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n37941), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS commutation_state_i0 (.Q(commutation_state[0]), .C(CLK_c), 
            .E(n6_adj_5228), .D(commutation_state_7__N_216[0]), .S(commutation_state_7__N_224));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n37941), .I0(n2233), 
            .I1(VCC_net), .CO(n37942));
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n7072), 
            .D(n1097), .R(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n37941));
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n47917), .I1(n2115), 
            .I2(VCC_net), .I3(n37940), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n37939), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n37939), .I0(n2116), 
            .I1(VCC_net), .CO(n37940));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n37938), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n37938), .I0(n2117), 
            .I1(VCC_net), .CO(n37939));
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n37937), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLA_181 (.Q(INLA_c_0), .C(CLK_c), .E(n27644), .D(GLA_N_384), 
            .R(n27973));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n37937), .I0(n2118), 
            .I1(VCC_net), .CO(n37938));
    SB_LUT4 mux_238_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[4]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n37936), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n37936), .I0(n2119), 
            .I1(VCC_net), .CO(n37937));
    SB_LUT4 encoder0_position_31__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[5]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n37935), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_10_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n37935), .I0(n2120), 
            .I1(VCC_net), .CO(n37936));
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n37934), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n37934), .I0(n2121), 
            .I1(VCC_net), .CO(n37935));
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n37933), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n37933), .I0(n2122), 
            .I1(VCC_net), .CO(n37934));
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n37932), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n37932), .I0(n2123), 
            .I1(VCC_net), .CO(n37933));
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n37931), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n37931), .I0(n2124), 
            .I1(VCC_net), .CO(n37932));
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n37930), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n37930), .I0(n2125), 
            .I1(VCC_net), .CO(n37931));
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n37929), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n37929), .I0(n2126), 
            .I1(VCC_net), .CO(n37930));
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n37928), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n37928), .I0(n2127), 
            .I1(VCC_net), .CO(n37929));
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n37927), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n37927), .I0(n2128), 
            .I1(VCC_net), .CO(n37928));
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n37926), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n37926), .I0(n2129), 
            .I1(GND_net), .CO(n37927));
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n37925), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n37925), .I0(n2130), 
            .I1(GND_net), .CO(n37926));
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n37924), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n37924), .I0(n2131), 
            .I1(VCC_net), .CO(n37925));
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n37923), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n37923), .I0(n2132), 
            .I1(GND_net), .CO(n37924));
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n37922), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n37922), .I0(n2133), 
            .I1(VCC_net), .CO(n37923));
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n37922));
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n48014), .I1(n2016), 
            .I2(VCC_net), .I3(n37921), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i28072_2_lut (.I0(n26494), .I1(n4452), .I2(GND_net), .I3(GND_net), 
            .O(n43094));
    defparam i28072_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n37920), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n37920), .I0(n2017), 
            .I1(VCC_net), .CO(n37921));
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n37919), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n37919), .I0(n2018), 
            .I1(VCC_net), .CO(n37920));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n37918), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n37422), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n37918), .I0(n2019), 
            .I1(VCC_net), .CO(n37919));
    SB_LUT4 add_145_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n37442), .O(n1080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_30 (.CI(n37442), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n37443));
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n37917), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n37917), .I0(n2020), 
            .I1(VCC_net), .CO(n37918));
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n37916), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n37916), .I0(n2021), 
            .I1(VCC_net), .CO(n37917));
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n37915), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n37915), .I0(n2022), 
            .I1(VCC_net), .CO(n37916));
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n37914), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_10 (.CI(n37422), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n37423));
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n37914), .I0(n2023), 
            .I1(VCC_net), .CO(n37915));
    SB_LUT4 add_145_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n37441), .O(n1081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n37913), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n37913), .I0(n2024), 
            .I1(VCC_net), .CO(n37914));
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n37912), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_29 (.CI(n37441), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n37442));
    SB_LUT4 add_145_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n37415), .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n37912), .I0(n2025), 
            .I1(VCC_net), .CO(n37913));
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n37911), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n37911), .I0(n2026), 
            .I1(VCC_net), .CO(n37912));
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n37910), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n37910), .I0(n2027), 
            .I1(VCC_net), .CO(n37911));
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n37909), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n37909), .I0(n2028), 
            .I1(VCC_net), .CO(n37910));
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n37908), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_3 (.CI(n37415), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n37416));
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n37908), .I0(n2029), 
            .I1(GND_net), .CO(n37909));
    SB_LUT4 add_145_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n37440), .O(n1082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_28 (.CI(n37440), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n37441));
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n37907), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n37421), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n37907), .I0(n2030), 
            .I1(GND_net), .CO(n37908));
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n37906), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_9 (.CI(n37421), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n37422));
    SB_LUT4 add_145_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n37439), .O(n1083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_27 (.CI(n37439), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n37440));
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n37906), .I0(n2031), 
            .I1(VCC_net), .CO(n37907));
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n37905), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n37905), .I0(n2032), 
            .I1(GND_net), .CO(n37906));
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n37904), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n37904), .I0(n2033), 
            .I1(VCC_net), .CO(n37905));
    SB_LUT4 add_145_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n37438), .O(n1084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n37904));
    SB_CARRY add_145_26 (.CI(n37438), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n37439));
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n48038), .I1(n1917), 
            .I2(VCC_net), .I3(n37903), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n37902), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n37902), .I0(n1918), 
            .I1(VCC_net), .CO(n37903));
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n37901), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n37901), .I0(n1919), 
            .I1(VCC_net), .CO(n37902));
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n37900), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n37900), .I0(n1920), 
            .I1(VCC_net), .CO(n37901));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n37899), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n37899), .I0(n1921), 
            .I1(VCC_net), .CO(n37900));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n37898), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n37898), .I0(n1922), 
            .I1(VCC_net), .CO(n37899));
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n37897), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n37897), .I0(n1923), 
            .I1(VCC_net), .CO(n37898));
    SB_LUT4 add_145_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n37420), .O(n1102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n37896), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n37896), .I0(n1924), 
            .I1(VCC_net), .CO(n37897));
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n37895), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n37895), .I0(n1925), 
            .I1(VCC_net), .CO(n37896));
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n37894), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_5255), .I3(n38456), .O(n2_adj_5227)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n37894), .I0(n1926), 
            .I1(VCC_net), .CO(n37895));
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n37893), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n37893), .I0(n1927), 
            .I1(VCC_net), .CO(n37894));
    SB_LUT4 encoder0_position_31__I_0_i1858_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_5256), .I3(n38455), .O(n3_adj_5226)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n37437), .O(n1085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n37892), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n37892), .I0(n1928), 
            .I1(VCC_net), .CO(n37893));
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n37891), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n38455), 
            .I0(GND_net), .I1(n3_adj_5256), .CO(n38456));
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n37891), .I0(n1929), 
            .I1(GND_net), .CO(n37892));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_5257), .I3(n38454), .O(n4_adj_5225)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n38454), 
            .I0(GND_net), .I1(n4_adj_5257), .CO(n38455));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_5258), .I3(n38453), .O(n5_adj_5224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_25 (.CI(n37437), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n37438));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n38453), 
            .I0(GND_net), .I1(n5_adj_5258), .CO(n38454));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_5259), .I3(n38452), .O(n6_adj_5217)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n38452), 
            .I0(GND_net), .I1(n6_adj_5259), .CO(n38453));
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n37890), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n37890), .I0(n1930), 
            .I1(GND_net), .CO(n37891));
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n37889), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n37889), .I0(n1931), 
            .I1(VCC_net), .CO(n37890));
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n37888), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n37888), .I0(n1932), 
            .I1(GND_net), .CO(n37889));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5260), .I3(n38451), .O(n7_adj_5215)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_224_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n37451), .O(encoder1_position_scaled_23__N_75[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_224_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n37887), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n38451), 
            .I0(GND_net), .I1(n7_adj_5260), .CO(n38452));
    SB_LUT4 add_145_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n37436), .O(n1086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n37887), .I0(n1933), 
            .I1(VCC_net), .CO(n37888));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5261), .I3(n38450), .O(n8_adj_5214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_24 (.CI(n37436), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n37437));
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n37887));
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n48064), .I1(n1818), 
            .I2(VCC_net), .I3(n37886), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n37885), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n37885), .I0(n1819), 
            .I1(VCC_net), .CO(n37886));
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n37884), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n37435), .O(n1087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n37884), .I0(n1820), 
            .I1(VCC_net), .CO(n37885));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n38450), 
            .I0(GND_net), .I1(n8_adj_5261), .CO(n38451));
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n37883), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n37883), .I0(n1821), 
            .I1(VCC_net), .CO(n37884));
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n37882), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n37882), .I0(n1822), 
            .I1(VCC_net), .CO(n37883));
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n37881), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n37881), .I0(n1823), 
            .I1(VCC_net), .CO(n37882));
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n37880), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n37880), .I0(n1824), 
            .I1(VCC_net), .CO(n37881));
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n37879), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n37879), .I0(n1825), 
            .I1(VCC_net), .CO(n37880));
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n37878), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n37878), .I0(n1826), 
            .I1(VCC_net), .CO(n37879));
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n37877), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5262), .I3(n38449), .O(n9_adj_5205)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n37877), .I0(n1827), 
            .I1(VCC_net), .CO(n37878));
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n37876), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n38449), 
            .I0(GND_net), .I1(n9_adj_5262), .CO(n38450));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5263), .I3(n38448), .O(n10_adj_5204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n37876), .I0(n1828), 
            .I1(VCC_net), .CO(n37877));
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n37875), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n37875), .I0(n1829), 
            .I1(GND_net), .CO(n37876));
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n37874), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_23 (.CI(n37435), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n37436));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n38448), 
            .I0(GND_net), .I1(n10_adj_5263), .CO(n38449));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5264), .I3(n38447), .O(n11_adj_5203)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n37874), .I0(n1830), 
            .I1(GND_net), .CO(n37875));
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n37873), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n38447), 
            .I0(GND_net), .I1(n11_adj_5264), .CO(n38448));
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n37873), .I0(n1831), 
            .I1(VCC_net), .CO(n37874));
    SB_LUT4 add_145_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n37434), .O(n1088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n37872), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n37872), .I0(n1832), 
            .I1(GND_net), .CO(n37873));
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n37871), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n38431), 
            .I0(GND_net), .I1(n27_adj_5280), .CO(n38432));
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n37871), .I0(n1833), 
            .I1(VCC_net), .CO(n37872));
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n37871));
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n48088), .I1(n1719), 
            .I2(VCC_net), .I3(n37870), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n37869), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n37869), .I0(n1720), 
            .I1(VCC_net), .CO(n37870));
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n37868), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n37868), .I0(n1721), 
            .I1(VCC_net), .CO(n37869));
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n37867), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n37867), .I0(n1722), 
            .I1(VCC_net), .CO(n37868));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n37866), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n37866), .I0(n1723), 
            .I1(VCC_net), .CO(n37867));
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n37865), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n37865), .I0(n1724), 
            .I1(VCC_net), .CO(n37866));
    SB_CARRY add_145_8 (.CI(n37420), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n37421));
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n37864), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_22 (.CI(n37434), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n37435));
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n37864), .I0(n1725), 
            .I1(VCC_net), .CO(n37865));
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n37863), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n37863), .I0(n1726), 
            .I1(VCC_net), .CO(n37864));
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n37862), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n37862), .I0(n1727), 
            .I1(VCC_net), .CO(n37863));
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n37861), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n37861), .I0(n1728), 
            .I1(VCC_net), .CO(n37862));
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n37860), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n37860), .I0(n1729), 
            .I1(GND_net), .CO(n37861));
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n37859), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n37433), .O(n1089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n37859), .I0(n1730), 
            .I1(GND_net), .CO(n37860));
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n37858), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n37858), .I0(n1731), 
            .I1(VCC_net), .CO(n37859));
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n37857), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_21 (.CI(n37433), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n37434));
    SB_LUT4 add_145_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n37432), .O(n1090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_20 (.CI(n37432), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n37433));
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n37857), .I0(n1732), 
            .I1(GND_net), .CO(n37858));
    SB_LUT4 add_145_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n37431), .O(n1091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n37419), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n37856), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF commutation_state_i2 (.Q(commutation_state[2]), .C(CLK_c), .D(n43084));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n37856), .I0(n1733), 
            .I1(VCC_net), .CO(n37857));
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n37856));
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n48112), .I1(n1620), 
            .I2(VCC_net), .I3(n37855), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n37854), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n37854), .I0(n1621), 
            .I1(VCC_net), .CO(n37855));
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n37853), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n37853), .I0(n1622), 
            .I1(VCC_net), .CO(n37854));
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n37852), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n37852), .I0(n1623), 
            .I1(VCC_net), .CO(n37853));
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n37851), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n37851), .I0(n1624), 
            .I1(VCC_net), .CO(n37852));
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n37850), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n37850), .I0(n1625), 
            .I1(VCC_net), .CO(n37851));
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n37849), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n37849), .I0(n1626), 
            .I1(VCC_net), .CO(n37850));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n37848), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n37848), .I0(n1627), 
            .I1(VCC_net), .CO(n37849));
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n37847), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n37847), .I0(n1628), 
            .I1(VCC_net), .CO(n37848));
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n37846), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n37846), .I0(n1629), 
            .I1(GND_net), .CO(n37847));
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n28611));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n37845), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n28610));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n28609));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n28608));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n37845), .I0(n1630), 
            .I1(GND_net), .CO(n37846));
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n28607));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n28606));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n28605));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n37844), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n37844), .I0(n1631), 
            .I1(VCC_net), .CO(n37845));
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632_adj_5239), 
            .I2(GND_net), .I3(n37843), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5273), .I3(n38438), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n37843), .I0(n1632_adj_5239), 
            .I1(GND_net), .CO(n37844));
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n37842), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n37842), .I0(n1633), 
            .I1(VCC_net), .CO(n37843));
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n37842));
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n48130), .I1(n1521), 
            .I2(VCC_net), .I3(n37841), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n37840), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n37840), .I0(n1522), 
            .I1(VCC_net), .CO(n37841));
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n37839), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n37839), .I0(n1523), 
            .I1(VCC_net), .CO(n37840));
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n37838), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n37838), .I0(n1524), 
            .I1(VCC_net), .CO(n37839));
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n37837), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n37837), .I0(n1525), 
            .I1(VCC_net), .CO(n37838));
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n37836), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n37836), .I0(n1526), 
            .I1(VCC_net), .CO(n37837));
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n37835), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_7 (.CI(n37419), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n37420));
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n37835), .I0(n1527), 
            .I1(VCC_net), .CO(n37836));
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n37834), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n37834), .I0(n1528), 
            .I1(VCC_net), .CO(n37835));
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n37833), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n37833), .I0(n1529), 
            .I1(GND_net), .CO(n37834));
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n37832), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_238_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[6]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n37832), .I0(n1530), 
            .I1(GND_net), .CO(n37833));
    SB_CARRY add_145_19 (.CI(n37431), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n37432));
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n37831), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLB_183 (.Q(INLB_c_0), .C(CLK_c), .E(n27644), .D(GLB_N_398), 
            .R(n27973));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n37831), .I0(n1531), 
            .I1(VCC_net), .CO(n37832));
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n37830), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n37830), .I0(n1532), 
            .I1(GND_net), .CO(n37831));
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n37829), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n37829), .I0(n1533), 
            .I1(VCC_net), .CO(n37830));
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n37829));
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n37415));
    SB_LUT4 add_145_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n37430), .O(n1092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n37418), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(n48147), .I1(n1422), 
            .I2(VCC_net), .I3(n37828), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n37827), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14789_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n23622), .I3(GND_net), .O(n28303));   // verilog/coms.v(127[12] 300[6])
    defparam i14789_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n37827), .I0(n1423), 
            .I1(VCC_net), .CO(n37828));
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n37826), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n37826), .I0(n1424), 
            .I1(VCC_net), .CO(n37827));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5264));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5263));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5262));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n37825), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n37825), .I0(n1425), 
            .I1(VCC_net), .CO(n37826));
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n37824), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n37824), .I0(n1426), 
            .I1(VCC_net), .CO(n37825));
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n37823), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_18 (.CI(n37430), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n37431));
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n37823), .I0(n1427), 
            .I1(VCC_net), .CO(n37824));
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n37822), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n37822), .I0(n1428), 
            .I1(VCC_net), .CO(n37823));
    SB_LUT4 add_145_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n37429), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n37821), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n37821), .I0(n1429), 
            .I1(GND_net), .CO(n37822));
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n37820), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n37820), .I0(n1430), 
            .I1(GND_net), .CO(n37821));
    SB_CARRY add_145_17 (.CI(n37429), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n37430));
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n37819), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n37819), .I0(n1431), 
            .I1(VCC_net), .CO(n37820));
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n37818), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n37818), .I0(n1432), 
            .I1(GND_net), .CO(n37819));
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n37817), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n37817), .I0(n1433), 
            .I1(VCC_net), .CO(n37818));
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n37428), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n37817));
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n48162), .I1(n1323), 
            .I2(VCC_net), .I3(n37816), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n37815), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n37815), .I0(n1324), 
            .I1(VCC_net), .CO(n37816));
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n37814), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n28427));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n37814), .I0(n1325), 
            .I1(VCC_net), .CO(n37815));
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n37813), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n37813), .I0(n1326), 
            .I1(VCC_net), .CO(n37814));
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n37812), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n37812), .I0(n1327), 
            .I1(VCC_net), .CO(n37813));
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n37811), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n37811), .I0(n1328), 
            .I1(VCC_net), .CO(n37812));
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n37810), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n37810), .I0(n1329), 
            .I1(GND_net), .CO(n37811));
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n37809), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n37809), .I0(n1330), 
            .I1(GND_net), .CO(n37810));
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n37808), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n37808), .I0(n1331), 
            .I1(VCC_net), .CO(n37809));
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n37807), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n37807), .I0(n1332), 
            .I1(GND_net), .CO(n37808));
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n37806), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n37806), .I0(n1333), 
            .I1(VCC_net), .CO(n37807));
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n37806));
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n48177), .I1(n1224), 
            .I2(VCC_net), .I3(n37805), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n37804), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n37804), .I0(n1225), 
            .I1(VCC_net), .CO(n37805));
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n37803), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n37803), .I0(n1226), 
            .I1(VCC_net), .CO(n37804));
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n37802), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n37802), .I0(n1227), 
            .I1(VCC_net), .CO(n37803));
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n37801), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n37801), .I0(n1228), 
            .I1(VCC_net), .CO(n37802));
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n37800), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n37800), .I0(n1229), 
            .I1(GND_net), .CO(n37801));
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n37799), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15148_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n42264), .I3(GND_net), .O(n28662));   // verilog/coms.v(127[12] 300[6])
    defparam i15148_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_145_16 (.CI(n37428), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n37429));
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n37799), .I0(n1230), 
            .I1(GND_net), .CO(n37800));
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n37798), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n37798), .I0(n1231), 
            .I1(VCC_net), .CO(n37799));
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n37797), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n37797), .I0(n1232), 
            .I1(GND_net), .CO(n37798));
    SB_DFF read_189 (.Q(read), .C(CLK_c), .D(n44724));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n37796), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n37796), .I0(n1233), 
            .I1(VCC_net), .CO(n37797));
    SB_DFF dir_175 (.Q(dir), .C(CLK_c), .D(pwm_setpoint_23__N_215));   // verilog/TinyFPGA_B.v(104[9] 114[5])
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n37796));
    SB_LUT4 add_145_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n37427), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_15 (.CI(n37427), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n37428));
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n48191), .I1(n1125), 
            .I2(VCC_net), .I3(n37795), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n37794), .O(n1193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n37794), .I0(n1126), 
            .I1(VCC_net), .CO(n37795));
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n37793), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR GLC_185 (.Q(INLC_c_0), .C(CLK_c), .E(n27644), .D(GLC_N_412), 
            .R(n27973));   // verilog/TinyFPGA_B.v(128[9] 207[5])
    SB_CARRY add_145_6 (.CI(n37418), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n37419));
    motorControl control (.\Ki[15] (Ki[15]), .GND_net(GND_net), .PWMLimit({PWMLimit}), 
            .\Kp[6] (Kp[6]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), 
            .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[7] (Kp[7]), 
            .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), 
            .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), 
            .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), 
            .\Ki[4] (Ki[4]), .\Ki[10] (Ki[10]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .IntegralLimit({IntegralLimit}), 
            .\Ki[9] (Ki[9]), .setpoint({setpoint}), .motor_state({motor_state}), 
            .duty({duty}), .clk32MHz(clk32MHz), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(271[16] 283[4])
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n37793), .I0(n1127), 
            .I1(VCC_net), .CO(n37794));
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n37792), .O(n1195_adj_5238)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n37792), .I0(n1128), 
            .I1(VCC_net), .CO(n37793));
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n37791), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_145_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n37426), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_145_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n37791), .I0(n1129), 
            .I1(GND_net), .CO(n37792));
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n37790), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2625_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n37527), 
            .O(n7646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2625_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n37790), .I0(n1130), 
            .I1(GND_net), .CO(n37791));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n38438), 
            .I0(GND_net), .I1(n20_adj_5273), .CO(n38439));
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n37789), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n37789), .I0(n1131), 
            .I1(VCC_net), .CO(n37790));
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n37788), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_145_14 (.CI(n37426), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n37427));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n38439), 
            .I0(GND_net), .I1(n19_adj_5272), .CO(n38440));
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5272), .I3(n38439), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n37788), .I0(n1132), 
            .I1(GND_net), .CO(n37789));
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n37787), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n37787), .I0(n1133), 
            .I1(VCC_net), .CO(n37788));
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n37787));
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n37786), .O(n1093_adj_5229)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15149_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n42264), .I3(GND_net), .O(n28663));   // verilog/coms.v(127[12] 300[6])
    defparam i15149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15150_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n42264), .I3(GND_net), .O(n28664));   // verilog/coms.v(127[12] 300[6])
    defparam i15150_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5357_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHA_N_367));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i5357_3_lut_4_lut_4_lut.LUT_INIT = 16'h12c2;
    SB_LUT4 unary_minus_10_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5138));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1853_3_lut (.I0(n2722), .I1(n2789), 
            .I2(n2742), .I3(GND_net), .O(n2821));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1852_3_lut (.I0(n2721), .I1(n2788), 
            .I2(n2742), .I3(GND_net), .O(n2820));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5359_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLA_N_384));   // verilog/TinyFPGA_B.v(164[7] 183[15])
    defparam i5359_3_lut_4_lut_4_lut.LUT_INIT = 16'h212c;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n2826), .I1(n2824), .I2(n2827), .I3(n2825), 
            .O(n45412));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1701 (.I0(tx_active), .I1(r_SM_Main_2__N_3616[0]), 
            .I2(n34010), .I3(n19799), .O(n19_adj_5253));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1701.LUT_INIT = 16'heeef;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5261));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1702 (.I0(n45412), .I1(n2820), .I2(n2821), .I3(GND_net), 
            .O(n45414));
    defparam i1_3_lut_adj_1702.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5281));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5260));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut (.I0(dti_counter[0]), .I1(n14_adj_5245), .I2(n10_adj_5246), 
            .I3(dti_counter[3]), .O(n23805));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n2819), .I1(n2822), .I2(n2828), .I3(n2823), 
            .O(n45416));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 i20581_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n34092));
    defparam i20581_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i5361_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GHB_N_389));
    defparam i5361_3_lut_4_lut_4_lut.LUT_INIT = 16'hc121;
    SB_LUT4 i5363_3_lut_4_lut_4_lut (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(dir), .I3(commutation_state[0]), .O(GLB_N_398));
    defparam i5363_3_lut_4_lut_4_lut.LUT_INIT = 16'h1c12;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5259));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n2817), .I1(n2818), .I2(n45416), .I3(n45414), 
            .O(n45422));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5258));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5257));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5256));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n2829), .I1(n45422), .I2(n34092), .I3(n2830), 
            .O(n45424));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'heccc;
    SB_LUT4 mux_236_i21_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[20]), .I3(encoder0_position_scaled[20]), 
            .O(motor_state[20]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i22_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[21]), .I3(encoder0_position_scaled[21]), 
            .O(motor_state[21]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14777_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n23622), .I3(GND_net), .O(n28291));   // verilog/coms.v(127[12] 300[6])
    defparam i14777_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i23_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[22]), .I3(encoder0_position_scaled[22]), 
            .O(motor_state[22]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n45424), 
            .O(n45430));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n45430), 
            .O(n45436));
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5286));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i33267_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n45436), 
            .O(n2841));
    defparam i33267_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5285));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i24_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[23]), .I3(encoder0_position_scaled[23]), 
            .O(motor_state[23]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i1_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_5205), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n934));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27978_3_lut (.I0(n4_adj_5225), .I1(n7648), .I2(n42988), .I3(GND_net), 
            .O(n42997));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27979_3_lut (.I0(encoder0_position[29]), .I1(n42997), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1708 (.I0(n5_adj_5157), .I1(n3_adj_5226), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n45272));
    defparam i1_3_lut_adj_1708.LUT_INIT = 16'h8080;
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut (.I0(n2_adj_5227), .I1(n7646), 
            .I2(n45272), .I3(encoder0_position[31]), .O(n828));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 mux_236_i2_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i27980_3_lut (.I0(n3_adj_5226), .I1(n7647), .I2(n42988), .I3(GND_net), 
            .O(n42999));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i3_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15151_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n42264), .I3(GND_net), .O(n28665));   // verilog/coms.v(127[12] 300[6])
    defparam i15151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_236_i4_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i5_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i6_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i7_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i8_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i27981_3_lut (.I0(encoder0_position[30]), .I1(n42999), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7_adj_5215), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n4_adj_5225), .I1(n5_adj_5224), .I2(n731), 
            .I3(n6_adj_5217), .O(n5_adj_5157));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'heeea;
    SB_LUT4 encoder0_position_31__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1710 (.I0(n3_adj_5226), .I1(n2_adj_5227), .I2(n5_adj_5157), 
            .I3(GND_net), .O(n42988));
    defparam i1_3_lut_adj_1710.LUT_INIT = 16'h8080;
    SB_LUT4 i28046_2_lut (.I0(n26482), .I1(n3303), .I2(GND_net), .I3(GND_net), 
            .O(n43068));
    defparam i28046_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i27970_3_lut (.I0(n7_adj_5215), .I1(n7651), .I2(n42988), .I3(GND_net), 
            .O(n42989));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27971_3_lut (.I0(encoder0_position[26]), .I1(n42989), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i9_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), .I2(motor_state_23__N_123[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i27974_3_lut (.I0(n6_adj_5217), .I1(n7650), .I2(n42988), .I3(GND_net), 
            .O(n42993));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i27975_3_lut (.I0(encoder0_position[27]), .I1(n42993), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_5214), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n834));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20603_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n34114));
    defparam i20603_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 mux_236_i10_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[9]), .I3(encoder0_position_scaled[9]), 
            .O(motor_state[9]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i20711_4_lut (.I0(n829), .I1(n828), .I2(n34114), .I3(n830), 
            .O(n861));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i20711_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i27976_3_lut (.I0(n5_adj_5224), .I1(n7649), .I2(n42988), .I3(GND_net), 
            .O(n42995));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27976_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i11_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[10]), .I3(encoder0_position_scaled[10]), 
            .O(motor_state[10]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i12_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[11]), .I3(encoder0_position_scaled[11]), 
            .O(motor_state[11]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i13_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[12]), .I3(encoder0_position_scaled[12]), 
            .O(motor_state[12]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i14_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[13]), .I3(encoder0_position_scaled[13]), 
            .O(motor_state[13]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i27977_3_lut (.I0(encoder0_position[28]), .I1(n42995), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i27977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_236_i15_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[14]), .I3(encoder0_position_scaled[14]), 
            .O(motor_state[14]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i20623_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n34134));
    defparam i20623_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1711 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n45172));
    defparam i1_2_lut_adj_1711.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n927), .I1(n45172), .I2(n928), .I3(n34134), 
            .O(n960));
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'hfefa;
    SB_LUT4 mux_236_i16_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[15]), .I3(encoder0_position_scaled[15]), 
            .O(motor_state[15]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5270));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_236_i17_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[16]), .I3(encoder0_position_scaled[16]), 
            .O(motor_state[16]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14778_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n23622), .I3(GND_net), .O(n28292));   // verilog/coms.v(127[12] 300[6])
    defparam i14778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_238_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[7]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5284));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_236_i18_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[17]), .I3(encoder0_position_scaled[17]), 
            .O(motor_state[17]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i19_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[18]), .I3(encoder0_position_scaled[18]), 
            .O(motor_state[18]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_236_i20_3_lut_4_lut (.I0(n26277), .I1(control_mode[1]), 
            .I2(motor_state_23__N_123[19]), .I3(encoder0_position_scaled[19]), 
            .O(motor_state[19]));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam mux_236_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n27716), 
            .I3(rx_data_ready), .O(n41875));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 unary_minus_10_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n27716));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h2505;
    SB_LUT4 i1_2_lut_4_lut_adj_1713 (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_5150), .I3(control_mode[2]), .O(n26277));   // verilog/TinyFPGA_B.v(266[5:22])
    defparam i1_2_lut_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1714 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3542[2]), .O(n42166));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut_adj_1714.LUT_INIT = 16'h2000;
    SB_LUT4 mux_238_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[8]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28062_4_lut_4_lut_4_lut (.I0(h1), .I1(h3), .I2(h2), .I3(commutation_state[2]), 
            .O(n43084));   // verilog/TinyFPGA_B.v(151[7:23])
    defparam i28062_4_lut_4_lut_4_lut.LUT_INIT = 16'hc544;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5274));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5275));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19784_1_lut_2_lut (.I0(n23805), .I1(dti), .I2(GND_net), .I3(GND_net), 
            .O(n1964));
    defparam i19784_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5276));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1792_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5277));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1786_3_lut (.I0(n2623), .I1(n2690), 
            .I2(n2643), .I3(GND_net), .O(n2722));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_10_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1785_3_lut (.I0(n2622), .I1(n2689), 
            .I2(n2643), .I3(GND_net), .O(n2721));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14966_3_lut_4_lut (.I0(n1673), .I1(b_prev_adj_5194), .I2(a_new_adj_5325[1]), 
            .I3(direction_N_3907_adj_5195), .O(n28480));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14966_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 encoder0_position_31__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1715 (.I0(n2727), .I1(n2725), .I2(GND_net), .I3(GND_net), 
            .O(n45136));
    defparam i1_2_lut_adj_1715.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n2724), .I1(n2721), .I2(n2722), .I3(n2728), 
            .O(n45138));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_LUT4 i14947_3_lut_4_lut (.I0(n1632), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_3907), .O(n28461));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14947_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n2723), .I1(n2720), .I2(n45136), .I3(n2726), 
            .O(n45142));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 i20583_4_lut (.I0(n952), .I1(n2731), .I2(n2732), .I3(n2733), 
            .O(n34094));
    defparam i20583_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n2718), .I1(n2719), .I2(n45142), .I3(n45138), 
            .O(n45148));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_5225), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n2729), .I1(n45148), .I2(n34094), .I3(n2730), 
            .O(n45150));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n2715), .I1(n2716), .I2(n45150), .I3(n2717), 
            .O(n45156));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3_adj_5226), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n45156), 
            .O(n45162));
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'hfffe;
    SB_LUT4 i14779_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n23622), .I3(GND_net), .O(n28293));   // verilog/coms.v(127[12] 300[6])
    defparam i14779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_5249));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12_adj_5249), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n26299));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i33300_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n45162), 
            .O(n2742));
    defparam i33300_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1722 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n26296));
    defparam i2_3_lut_adj_1722.LUT_INIT = 16'hfefe;
    \grp_debouncer(3,1000)  debounce (.reg_B({reg_B}), .CLK_c(CLK_c), .GND_net(GND_net), 
            .VCC_net(VCC_net), .data_i({hall1, hall2, hall3}), .n28167(n28167), 
            .data_o({h1, h2, h3}), .n44732(n44732), .n28614(n28614), 
            .n28613(n28613));   // verilog/TinyFPGA_B.v(98[26] 102[3])
    SB_LUT4 i5_3_lut_adj_1723 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14));
    defparam i5_3_lut_adj_1723.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1724 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15));
    defparam i6_4_lut_adj_1724.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(delay_counter[2]), .I2(n14), .I3(delay_counter[6]), 
            .O(n26302));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4511_4_lut (.I0(n26302), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_5243));
    defparam i4511_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1725 (.I0(n24_adj_5243), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n44392));
    defparam i2_4_lut_adj_1725.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1726 (.I0(n44392), .I1(delay_counter[18]), .I2(n26296), 
            .I3(GND_net), .O(n44233));
    defparam i2_3_lut_adj_1726.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1727 (.I0(delay_counter[23]), .I1(n44233), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7_adj_5156));
    defparam i2_4_lut_adj_1727.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_1728 (.I0(n7_adj_5156), .I1(delay_counter[21]), 
            .I2(delay_counter[22]), .I3(n26299), .O(n62_adj_5244));
    defparam i4_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1729 (.I0(n62_adj_5244), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(delay_counter[31]), .I3(GND_net), .O(n4_adj_5216));
    defparam i1_3_lut_adj_1729.LUT_INIT = 16'hcece;
    SB_LUT4 i1_2_lut_adj_1730 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_5155));
    defparam i1_2_lut_adj_1730.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1731 (.I0(delay_counter[9]), .I1(n4_adj_5155), 
            .I2(delay_counter[10]), .I3(n26302), .O(n44389));
    defparam i2_4_lut_adj_1731.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1732 (.I0(n44389), .I1(n26296), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n44235));
    defparam i2_4_lut_adj_1732.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5152));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1733 (.I0(delay_counter[22]), .I1(n44235), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5154));
    defparam i2_4_lut_adj_1733.LUT_INIT = 16'ha8a0;
    SB_LUT4 i19910_4_lut (.I0(n7_adj_5154), .I1(delay_counter[31]), .I2(n26299), 
            .I3(n8_adj_5152), .O(n1195));   // verilog/TinyFPGA_B.v(378[14:38])
    defparam i19910_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5190));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1734 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_5185));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i6_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1735 (.I0(ID[3]), .I1(n14_adj_5185), .I2(n10_adj_5190), 
            .I3(ID[6]), .O(n26285));   // verilog/TinyFPGA_B.v(376[12:17])
    defparam i7_4_lut_adj_1735.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14599_4_lut (.I0(n7072), .I1(n1195), .I2(n4_adj_5216), .I3(n26286), 
            .O(n28084));   // verilog/TinyFPGA_B.v(357[10] 385[6])
    defparam i14599_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5364[2]), .I1(r_SM_Main_adj_5364[0]), 
            .I2(r_SM_Main_adj_5364[1]), .I3(r_SM_Main_2__N_3613[1]), .O(n48874));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 encoder0_position_31__I_0_i1723_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1723_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14780_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n23622), .I3(GND_net), .O(n28294));   // verilog/coms.v(127[12] 300[6])
    defparam i14780_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14781_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n23622), .I3(GND_net), .O(n28295));   // verilog/coms.v(127[12] 300[6])
    defparam i14781_3_lut.LUT_INIT = 16'hcaca;
    \quadrature_decoder(1,500000)  quad_counter1 (.a_new({a_new_adj_5325[1], 
            Open_0}), .ENCODER1_B_N_keep(ENCODER1_B_N), .n1668(CLK_c), 
            .ENCODER1_A_N_keep(ENCODER1_A_N), .encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .direction_N_3907(direction_N_3907_adj_5195), 
            .b_prev(b_prev_adj_5194), .n28480(n28480), .n1673(n1673)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(294[57] 301[6])
    SB_LUT4 encoder0_position_31__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32138_3_lut_4_lut (.I0(n2346), .I1(n2247), .I2(n2227), .I3(n45734), 
            .O(n2425));
    defparam i32138_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5282));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14652_3_lut_4_lut (.I0(\data_out_frame[27] [0]), .I1(n40583), 
            .I2(n42299), .I3(n27647), .O(n28166));   // verilog/coms.v(127[12] 300[6])
    defparam i14652_3_lut_4_lut.LUT_INIT = 16'hc3aa;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(commutation_state[2]), .I1(commutation_state[1]), 
            .I2(commutation_state_prev[2]), .I3(commutation_state_prev[1]), 
            .O(n4_adj_5247));   // verilog/TinyFPGA_B.v(131[7:48])
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'h7bde;
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_adj_1737 (.I0(dti_counter[1]), .I1(dti_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5246));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i2_2_lut_adj_1737.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i32375_3_lut (.I0(n2523), .I1(n2590), .I2(n2544), .I3(GND_net), 
            .O(n2622));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1720_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1720_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1724_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1724_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14757_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n44019), 
            .I3(GND_net), .O(n28271));   // verilog/coms.v(127[12] 300[6])
    defparam i14757_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1722_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_i1722_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_238_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[9]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14758_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n23622), .I3(GND_net), .O(n28272));   // verilog/coms.v(127[12] 300[6])
    defparam i14758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32561_3_lut (.I0(n2522), .I1(n2589), .I2(n2544), .I3(GND_net), 
            .O(n2621));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam i32561_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5278));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1738 (.I0(dti_counter[7]), .I1(dti_counter[4]), 
            .I2(dti_counter[5]), .I3(dti_counter[6]), .O(n14_adj_5245));   // verilog/TinyFPGA_B.v(156[9:23])
    defparam i6_4_lut_adj_1738.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n2623), .I1(n2628), .I2(n2624), .I3(n2622), 
            .O(n45374));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_238_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15_adj_5191), .I3(n15_adj_5158), .O(motor_state_23__N_123[10]));   // verilog/TinyFPGA_B.v(267[5] 269[10])
    defparam mux_238_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_3_lut_adj_1740 (.I0(n45374), .I1(n2621), .I2(n2626), .I3(GND_net), 
            .O(n45376));
    defparam i1_3_lut_adj_1740.LUT_INIT = 16'hfefe;
    SB_LUT4 i20585_4_lut (.I0(n951), .I1(n2631), .I2(n2632), .I3(n2633), 
            .O(n34096));
    defparam i20585_4_lut.LUT_INIT = 16'hfcec;
    EEPROM eeprom (.CLK_c(CLK_c), .read(read), .\state[0] (state_adj_5349[0]), 
           .enable_slow_N_4190(enable_slow_N_4190), .n5614({n5615}), .\state[1] (state_adj_5349[1]), 
           .n41883(n41883), .n41869(n41869), .n28229(n28229), .rw(rw), 
           .n41973(n41973), .data_ready(data_ready), .\state[3] (state_adj_5377[3]), 
           .n6(n6), .GND_net(GND_net), .\state[2] (state_adj_5377[2]), 
           .n7(n7_adj_5250), .n33881(n33881), .n43114(n43114), .n42289(n42289), 
           .scl_enable(scl_enable), .scl(scl), .\state_7__N_4103[3] (state_7__N_4103[3]), 
           .\state[0]_adj_13 (state_adj_5377[0]), .n33185(n33185), .n6692(n6692), 
           .\saved_addr[0] (saved_addr[0]), .VCC_net(VCC_net), .n4(n4_adj_5218), 
           .n4_adj_14(n4_adj_5192), .n33292(n33292), .sda_enable(sda_enable), 
           .\state_7__N_4087[0] (state_7__N_4087[0]), .n28193(n28193), .data({data}), 
           .n28192(n28192), .n28191(n28191), .n28190(n28190), .n28189(n28189), 
           .n28188(n28188), .n28187(n28187), .n10(n10_adj_5251), .n8(n8_adj_5241), 
           .n28330(n28330), .n28315(n28315), .n7233(n7233), .n26424(n26424), 
           .n26409(n26409), .sda_out(sda_out), .n46890(n46890)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(387[10] 398[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5280));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15152_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n42264), .I3(GND_net), .O(n28666));   // verilog/coms.v(127[12] 300[6])
    defparam i15152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15153_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n42264), .I3(GND_net), .O(n28667));   // verilog/coms.v(127[12] 300[6])
    defparam i15153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15154_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n42264), .I3(GND_net), .O(n28668));   // verilog/coms.v(127[12] 300[6])
    defparam i15154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1741 (.I0(n2618), .I1(n2619), .I2(n45376), .I3(n2620), 
            .O(n45382));
    defparam i1_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_3_lut (.I0(h2), .I1(h3), .I2(h1), .I3(GND_net), .O(n6_adj_5228));
    defparam i14_3_lut.LUT_INIT = 16'h7e7e;
    SB_LUT4 i1_3_lut_adj_1742 (.I0(h3), .I1(h2), .I2(h1), .I3(GND_net), 
            .O(commutation_state_7__N_216[0]));   // verilog/TinyFPGA_B.v(148[4] 150[7])
    defparam i1_3_lut_adj_1742.LUT_INIT = 16'h1414;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5279));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    TLI4970 tli (.GND_net(GND_net), .CS_c(CS_c), .CS_CLK_c(CS_CLK_c), 
            .n5(n5_adj_5186), .n5_adj_11(n5_adj_5196), .n33328(n33328), 
            .CLK_c(CLK_c), .VCC_net(VCC_net), .\data[15] (data_adj_5353[15]), 
            .n43722(n43722), .n28227(n28227), .current({current}), .n28692(n28692), 
            .n28691(n28691), .n28690(n28690), .n28689(n28689), .n28688(n28688), 
            .n28687(n28687), .n28686(n28686), .n28685(n28685), .n28684(n28684), 
            .n28683(n28683), .n28682(n28682), .n28681(n28681), .n28185(n28185), 
            .n28184(n28184), .\data[12] (data_adj_5353[12]), .n28183(n28183), 
            .\data[11] (data_adj_5353[11]), .n28182(n28182), .\data[10] (data_adj_5353[10]), 
            .n28181(n28181), .\data[9] (data_adj_5353[9]), .n28180(n28180), 
            .\data[8] (data_adj_5353[8]), .n28179(n28179), .\data[7] (data_adj_5353[7]), 
            .n28178(n28178), .\data[6] (data_adj_5353[6]), .n28177(n28177), 
            .\data[5] (data_adj_5353[5]), .n28176(n28176), .\data[4] (data_adj_5353[4]), 
            .n28175(n28175), .\data[3] (data_adj_5353[3]), .n28174(n28174), 
            .\data[2] (data_adj_5353[2]), .n28173(n28173), .\data[1] (data_adj_5353[1]), 
            .state_7__N_4293(state_7__N_4293), .n28458(n28458), .\data[0] (data_adj_5353[0]), 
            .n9(n9_adj_5198), .n11(n11_adj_5197), .n26432(n26432), .n26440(n26440), 
            .n26445(n26445), .n26435(n26435)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(400[11] 406[4])
    SB_LUT4 i1_2_lut_adj_1743 (.I0(n2625), .I1(n2627), .I2(GND_net), .I3(GND_net), 
            .O(n45534));
    defparam i1_2_lut_adj_1743.LUT_INIT = 16'heeee;
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.b_prev(b_prev), .a_new({a_new[1], 
            Open_1}), .encoder0_position({encoder0_position}), .GND_net(GND_net), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1668(CLK_c), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .VCC_net(VCC_net), .direction_N_3907(direction_N_3907), .n28461(n28461), 
            .n1632(n1632)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(285[57] 292[6])
    SB_LUT4 i14643_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n27617), .I3(GND_net), .O(n28157));   // verilog/coms.v(127[12] 300[6])
    defparam i14643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15155_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n42264), .I3(GND_net), .O(n28669));   // verilog/coms.v(127[12] 300[6])
    defparam i15155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5283));   // verilog/TinyFPGA_B.v(320[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n2629), .I1(n45382), .I2(n34096), .I3(n2630), 
            .O(n45384));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'heccc;
    pwm PWM (.pwm_out(pwm_out), .clk32MHz(clk32MHz), .GND_net(GND_net), 
        .VCC_net(VCC_net), .pwm_setpoint({pwm_setpoint})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    SB_LUT4 unary_minus_10_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5149));   // verilog/TinyFPGA_B.v(111[22:27])
    defparam unary_minus_10_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    coms neopxl_color_23__I_0 (.n28303(n28303), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .CLK_c(CLK_c), .\data_out_frame[20] ({\data_out_frame[20] }), .GND_net(GND_net), 
         .n28302(n28302), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n28301(n28301), .n28300(n28300), .n28299(n28299), .n28298(n28298), 
         .n28297(n28297), .n28296(n28296), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .n27647(n27647), 
         .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n40583(n40583), .n28295(n28295), .n28294(n28294), .n28293(n28293), 
         .n28292(n28292), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\data_out_frame[22] ({\data_out_frame[22] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .\data_out_frame[21][2] (\data_out_frame[21] [2]), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\FRAME_MATCHER.state ({Open_2, 
         Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, Open_9, 
         Open_10, Open_11, Open_12, Open_13, Open_14, Open_15, Open_16, 
         Open_17, Open_18, Open_19, Open_20, Open_21, Open_22, Open_23, 
         Open_24, Open_25, Open_26, Open_27, Open_28, Open_29, \FRAME_MATCHER.state [3], 
         Open_30, Open_31, \FRAME_MATCHER.state [0]}), .n28291(n28291), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .\data_out_frame[21][1] (\data_out_frame[21] [1]), 
         .n28290(n28290), .\data_in_frame[14] ({\data_in_frame[14] }), .\data_in_frame[19] ({\data_in_frame[19] }), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[10] ({\data_in_frame[10] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_in_frame[7] ({\data_in_frame[7] }), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .n28289(n28289), .\data_in_frame[8] ({\data_in_frame[8] }), .n27617(n27617), 
         .rx_data({rx_data}), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .\r_SM_Main_2__N_3616[0] (r_SM_Main_2__N_3616[0]), 
         .\data_out_frame[21][0] (\data_out_frame[21] [0]), .rx_data_ready(rx_data_ready), 
         .setpoint({setpoint}), .\data_out_frame[21][3] (\data_out_frame[21] [3]), 
         .n28288(n28288), .n28287(n28287), .n28286(n28286), .n28285(n28285), 
         .n28284(n28284), .n28283(n28283), .n28282(n28282), .\data_out_frame[21][4] (\data_out_frame[21] [4]), 
         .n28281(n28281), .n28280(n28280), .n28279(n28279), .n28278(n28278), 
         .n28277(n28277), .n28276(n28276), .n28275(n28275), .n28274(n28274), 
         .n28273(n28273), .\Kp[13] (Kp[13]), .n42276(n42276), .n42287(n42287), 
         .n42266(n42266), .n28272(n28272), .n28271(n28271), .\Ki[11] (Ki[11]), 
         .DE_c(DE_c), .n28270(n28270), .\Kp[12] (Kp[12]), .n28269(n28269), 
         .\Ki[12] (Ki[12]), .n28268(n28268), .\Ki[13] (Ki[13]), .n28267(n28267), 
         .\Ki[14] (Ki[14]), .n28266(n28266), .n28265(n28265), .\Kp[11] (Kp[11]), 
         .n28264(n28264), .\Ki[15] (Ki[15]), .n28263(n28263), .n28262(n28262), 
         .n28261(n28261), .n28260(n28260), .n28259(n28259), .n28258(n28258), 
         .n28257(n28257), .n28256(n28256), .n28255(n28255), .n28254(n28254), 
         .n28253(n28253), .\data_out_frame[27][0] (\data_out_frame[27] [0]), 
         .n28252(n28252), .ID({ID}), .n122(n122), .\FRAME_MATCHER.state_31__N_2660[2] (\FRAME_MATCHER.state_31__N_2660 [2]), 
         .n26494(n26494), .n4452(n4452), .n7(n7_adj_5248), .n3303(n3303), 
         .\FRAME_MATCHER.state_31__N_2788[2] (\FRAME_MATCHER.state_31__N_2788 [2]), 
         .n28251(n28251), .n28783(n28783), .neopxl_color({neopxl_color}), 
         .n28782(n28782), .n28781(n28781), .n28780(n28780), .n28779(n28779), 
         .n28778(n28778), .n28777(n28777), .n28776(n28776), .n28775(n28775), 
         .n28774(n28774), .n28773(n28773), .n28772(n28772), .n28771(n28771), 
         .n28770(n28770), .n28250(n28250), .n28249(n28249), .n28248(n28248), 
         .n28247(n28247), .n28246(n28246), .n28245(n28245), .n28244(n28244), 
         .n28243(n28243), .\Kp[14] (Kp[14]), .n28242(n28242), .n28241(n28241), 
         .\data_in[2] ({\data_in[2] }), .n28240(n28240), .n28239(n28239), 
         .n28238(n28238), .n28237(n28237), .n28236(n28236), .n28234(n28234), 
         .\Kp[10] (Kp[10]), .n28233(n28233), .\Kp[9] (Kp[9]), .n28232(n28232), 
         .n28226(n28226), .\Kp[8] (Kp[8]), .n28225(n28225), .\Kp[7] (Kp[7]), 
         .n28224(n28224), .\Kp[6] (Kp[6]), .n28223(n28223), .\Kp[5] (Kp[5]), 
         .n28222(n28222), .\Kp[4] (Kp[4]), .n28221(n28221), .n41665(n41665), 
         .n28219(n28219), .PWMLimit({PWMLimit}), .n28218(n28218), .\data_in[3] ({\data_in[3] }), 
         .LED_c(LED_c), .n28217(n28217), .control_mode({control_mode}), 
         .n28215(n28215), .n28214(n28214), .\Kp[3] (Kp[3]), .n28213(n28213), 
         .\Ki[0] (Ki[0]), .n28212(n28212), .\Kp[0] (Kp[0]), .n28211(n28211), 
         .\data_in[0] ({\data_in[0] }), .n28210(n28210), .\Kp[2] (Kp[2]), 
         .n28209(n28209), .\Kp[1] (Kp[1]), .n28208(n28208), .n28207(n28207), 
         .n28206(n28206), .n28205(n28205), .n28204(n28204), .n28202(n28202), 
         .n28746(n28746), .n28745(n28745), .n28744(n28744), .n28743(n28743), 
         .n28742(n28742), .n28741(n28741), .n28740(n28740), .n28739(n28739), 
         .n28730(n28730), .n28729(n28729), .n28728(n28728), .n28727(n28727), 
         .n28726(n28726), .n28725(n28725), .n28724(n28724), .n28723(n28723), 
         .n28714(n28714), .n28713(n28713), .n28712(n28712), .n28711(n28711), 
         .n28710(n28710), .n28709(n28709), .n28708(n28708), .n28707(n28707), 
         .n28169(n28169), .n28168(n28168), .IntegralLimit({IntegralLimit}), 
         .n28166(n28166), .n28164(n28164), .n28163(n28163), .n28162(n28162), 
         .n28161(n28161), .n28160(n28160), .n19799(n19799), .n34010(n34010), 
         .n23516(n23516), .n28159(n28159), .n28158(n28158), .\data_in[1] ({\data_in[1] }), 
         .n23622(n23622), .n42267(n42267), .n42288(n42288), .n28669(n28669), 
         .n28157(n28157), .n28668(n28668), .n28667(n28667), .n28666(n28666), 
         .n28665(n28665), .n42244(n42244), .n43094(n43094), .n26482(n26482), 
         .n62(n62), .n28664(n28664), .n28663(n28663), .n28662(n28662), 
         .n19(n19_adj_5253), .n28652(n28652), .n28651(n28651), .n28650(n28650), 
         .n28618(n28618), .n28617(n28617), .n28616(n28616), .n28615(n28615), 
         .n28612(n28612), .n28604(n28604), .n28603(n28603), .n28602(n28602), 
         .n28601(n28601), .n28600(n28600), .n28599(n28599), .n28598(n28598), 
         .n28597(n28597), .n28596(n28596), .n28595(n28595), .n28594(n28594), 
         .n28593(n28593), .n28592(n28592), .n28591(n28591), .n28590(n28590), 
         .n28589(n28589), .n28588(n28588), .n28587(n28587), .n28586(n28586), 
         .n28585(n28585), .n28584(n28584), .n28583(n28583), .n28582(n28582), 
         .n28581(n28581), .n28580(n28580), .n28579(n28579), .n28578(n28578), 
         .n28577(n28577), .n28576(n28576), .n28575(n28575), .n28574(n28574), 
         .n28573(n28573), .n28572(n28572), .n28571(n28571), .n20(n20_adj_5252), 
         .n28546(n28546), .n28545(n28545), .n28544(n28544), .n28543(n28543), 
         .n28542(n28542), .n28541(n28541), .n28540(n28540), .n28539(n28539), 
         .n28530(n28530), .n28529(n28529), .n28528(n28528), .n28527(n28527), 
         .n28526(n28526), .n28525(n28525), .n28524(n28524), .n28523(n28523), 
         .n28522(n28522), .n28521(n28521), .n28520(n28520), .n28519(n28519), 
         .n28518(n28518), .n28517(n28517), .n28516(n28516), .n28515(n28515), 
         .n28514(n28514), .n28510(n28510), .n28509(n28509), .n28508(n28508), 
         .n28507(n28507), .n28506(n28506), .n28505(n28505), .n28501(n28501), 
         .n28500(n28500), .n28499(n28499), .n28498(n28498), .n28497(n28497), 
         .n28496(n28496), .n28495(n28495), .n28494(n28494), .n28493(n28493), 
         .n28492(n28492), .n28491(n28491), .n28490(n28490), .n28489(n28489), 
         .n28488(n28488), .n28487(n28487), .n28483(n28483), .n28482(n28482), 
         .n28479(n28479), .n28478(n28478), .n28477(n28477), .n28476(n28476), 
         .n28475(n28475), .n28474(n28474), .n28473(n28473), .n28472(n28472), 
         .n28471(n28471), .n48873(n48873), .n28469(n28469), .n28468(n28468), 
         .n28467(n28467), .n28466(n28466), .n28465(n28465), .n28464(n28464), 
         .n28463(n28463), .n28462(n28462), .n28457(n28457), .n28456(n28456), 
         .n28455(n28455), .n28454(n28454), .n28453(n28453), .n28452(n28452), 
         .n28451(n28451), .n28450(n28450), .n28449(n28449), .n28448(n28448), 
         .n28447(n28447), .n28446(n28446), .n28445(n28445), .n28444(n28444), 
         .n28443(n28443), .n28442(n28442), .n28441(n28441), .n28440(n28440), 
         .n28439(n28439), .n28438(n28438), .n28433(n28433), .n28432(n28432), 
         .n28428(n28428), .n28426(n28426), .\Ki[1] (Ki[1]), .n28425(n28425), 
         .n28424(n28424), .\Ki[2] (Ki[2]), .n28423(n28423), .n28422(n28422), 
         .n28421(n28421), .n28420(n28420), .n28419(n28419), .n28418(n28418), 
         .n28417(n28417), .n28416(n28416), .n28415(n28415), .n28414(n28414), 
         .n28413(n28413), .n28412(n28412), .n28411(n28411), .n28410(n28410), 
         .n28409(n28409), .n28408(n28408), .n28407(n28407), .n28406(n28406), 
         .n28405(n28405), .n28404(n28404), .n28403(n28403), .n28402(n28402), 
         .n28401(n28401), .n28400(n28400), .n28399(n28399), .n28398(n28398), 
         .n28397(n28397), .n28396(n28396), .n28395(n28395), .n28394(n28394), 
         .n28393(n28393), .n28392(n28392), .n28391(n28391), .n28390(n28390), 
         .n28389(n28389), .n28384(n28384), .n28383(n28383), .\Ki[3] (Ki[3]), 
         .n28382(n28382), .\Ki[4] (Ki[4]), .n28381(n28381), .n28380(n28380), 
         .n28379(n28379), .\Ki[5] (Ki[5]), .n28378(n28378), .n28377(n28377), 
         .n28376(n28376), .n28375(n28375), .n28374(n28374), .n28373(n28373), 
         .n28372(n28372), .n28371(n28371), .n28370(n28370), .n28369(n28369), 
         .n28368(n28368), .n28367(n28367), .n28366(n28366), .n28365(n28365), 
         .n28364(n28364), .n28363(n28363), .n28362(n28362), .n28361(n28361), 
         .n28360(n28360), .n28359(n28359), .n28358(n28358), .n28357(n28357), 
         .n28356(n28356), .n28355(n28355), .n28354(n28354), .n28353(n28353), 
         .n28352(n28352), .n28351(n28351), .n28350(n28350), .n28349(n28349), 
         .n28348(n28348), .n28347(n28347), .n28346(n28346), .n28345(n28345), 
         .n28344(n28344), .n28343(n28343), .n28342(n28342), .n28341(n28341), 
         .n28340(n28340), .n28335(n28335), .n28331(n28331), .n28329(n28329), 
         .n28328(n28328), .n28327(n28327), .n28326(n28326), .n28325(n28325), 
         .n28324(n28324), .n28323(n28323), .n28322(n28322), .n28321(n28321), 
         .n28320(n28320), .n28319(n28319), .\Ki[6] (Ki[6]), .n28317(n28317), 
         .n28316(n28316), .n28314(n28314), .\Kp[15] (Kp[15]), .n28313(n28313), 
         .n28312(n28312), .n28311(n28311), .\Ki[7] (Ki[7]), .n28310(n28310), 
         .\Ki[8] (Ki[8]), .n28309(n28309), .\Ki[9] (Ki[9]), .n28308(n28308), 
         .n28156(n28156), .n28307(n28307), .\Ki[10] (Ki[10]), .n28306(n28306), 
         .n28305(n28305), .n28304(n28304), .n60(n60), .n6(n6_adj_5159), 
         .tx_active(tx_active), .\state[0] (state_adj_5377[0]), .\state[2] (state_adj_5377[2]), 
         .\state[3] (state_adj_5377[3]), .n7233(n7233), .n43068(n43068), 
         .n42251(n42251), .n42255(n42255), .n42299(n42299), .n32652(n32652), 
         .n42277(n42277), .n42264(n42264), .n42285(n42285), .n44019(n44019), 
         .\r_Bit_Index[0] (r_Bit_Index_adj_5366[0]), .n27840(n27840), .r_SM_Main({r_SM_Main_adj_5364}), 
         .n28123(n28123), .\r_SM_Main_2__N_3613[1] (r_SM_Main_2__N_3613[1]), 
         .tx_o(tx_o), .VCC_net(VCC_net), .n28387(n28387), .n28235(n28235), 
         .n18934(n18934), .n4(n4_adj_5153), .n48874(n48874), .tx_enable(tx_enable), 
         .\r_Bit_Index[0]_adj_3 (r_Bit_Index[0]), .n27844(n27844), .r_SM_Main_adj_10({r_SM_Main}), 
         .n28125(n28125), .\r_SM_Main_2__N_3542[2] (r_SM_Main_2__N_3542[2]), 
         .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), .n4_adj_7(n4_adj_5200), 
         .n4_adj_8(n4_adj_5184), .n4_adj_9(n4_adj_5199), .n26398(n26398), 
         .n26390(n26390), .n33332(n33332), .n28431(n28431), .n41875(n41875), 
         .n28203(n28203), .n28201(n28201), .n28200(n28200), .n28199(n28199), 
         .n28198(n28198), .n28197(n28197), .n28196(n28196), .n42166(n42166), 
         .n28437(n28437)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(238[8] 261[4])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (\neo_pixel_transmitter.t0 , GND_net, 
            CLK_c, \state[1] , n41203, VCC_net, timer, neopxl_color, 
            n43011, \state_3__N_528[1] , n27791, n28195, n28165, LED_c, 
            n28649, n28648, n28647, n28646, n28645, n28644, n28643, 
            n28642, n28641, n28640, n28639, n28638, n28637, n28636, 
            n28635, n28634, n28633, n28632, n28631, n28630, n28629, 
            n28628, n28627, n28626, n28625, n28624, n28623, n28622, 
            n28621, n28620, n28619, NEOPXL_c) /* synthesis syn_module_defined=1 */ ;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input GND_net;
    input CLK_c;
    output \state[1] ;
    output n41203;
    input VCC_net;
    output [31:0]timer;
    input [23:0]neopxl_color;
    output n43011;
    output \state_3__N_528[1] ;
    output n27791;
    input n28195;
    input n28165;
    input LED_c;
    input n28649;
    input n28648;
    input n28647;
    input n28646;
    input n28645;
    input n28644;
    input n28643;
    input n28642;
    input n28641;
    input n28640;
    input n28639;
    input n28638;
    input n28637;
    input n28636;
    input n28635;
    input n28634;
    input n28633;
    input n28632;
    input n28631;
    input n28630;
    input n28629;
    input n28628;
    input n28627;
    input n28626;
    input n28625;
    input n28624;
    input n28623;
    input n28622;
    input n28621;
    input n28620;
    input n28619;
    output NEOPXL_c;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [31:0]n1;
    
    wire n37471;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n37472, n33857;
    wire [31:0]color_bit_N_722;
    
    wire \neo_pixel_transmitter.done_N_736 , n48855, \neo_pixel_transmitter.done , 
        start_N_727, n7, start;
    wire [31:0]n282;
    
    wire n27646, n28039, n37470, n26283, n43104, n39092;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire n43208, n7_adj_5134, n26417, n34074, n37469, n47200, n46811, 
        n34008, n43212, n47201, n43230, \neo_pixel_transmitter.done_N_742 ;
    wire [31:0]n133;
    
    wire n38277, n38276, n38275, n38274, n38273, n38272, n38271, 
        n38270, n38269, n38268, n38267, n38266, n38265, n38264, 
        n38263, n38262, n38261, n38260, n38259, n38258, n38257, 
        n38256, n38255, n38254, n38253, n38252, n38251, n38250, 
        n38249, n38248, n38247, n48784, n48787, n26449, n37657, 
        n45586, n37656, n45584, n37655, n45582, n37654, n45580, 
        n37653, n45578, n37652, n45576, n37651, n45574, n37650, 
        n45572, n48724, n48727, n48712, n48715, n48706, n48709, 
        n1991, n46813, n45968, n48601, n47450, n49107, n39590, 
        n47528, n48619, n46833;
    wire [3:0]state_3__N_528;
    
    wire n37649, n45570, n37648, n45568, n37647, n45566, n37646, 
        n45564, n37645, n45562, n37644, n45560, n37643, n45558, 
        n37642, n45556, n37641, n45554, n37640, n45552, n37639, 
        n45550, n37638;
    wire [31:0]one_wire_N_679;
    
    wire n48616, n37637, n37636, n37635, n37634, n37633, n37632, 
        n37499, n37631, n37630, n37498, n30, n48, n46, n47, 
        n45, n37629, n37628, n43001, n37627, n37497, n37496, n37495, 
        n37494, n37493, n37492, n37491, n44, n37490, n43, n37489, 
        n54, n37488, n49, n37487, n37486, n37485, n37484, n37483, 
        n1977, n37482, n37481, n37480, n37479, n37478, n37477, 
        n37476, n33935, n6921, n46884, n37475, n37474, n48598, 
        n37473, n44844, n42982, n45588, n45594, n46823, n43181, 
        n43100, n42246, n103, n16_adj_5136, n6_adj_5137;
    
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_5 (.CI(n37471), .I0(bit_ctr[3]), .I1(GND_net), .CO(n37472));
    SB_LUT4 i20354_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n33857));
    defparam i20354_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(color_bit_N_722[2]));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h1e1e;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n48855), .D(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE start_103 (.Q(start), .C(CLK_c), .E(n7), .D(start_N_727));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n27646), .D(n282[1]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n27646), .D(n282[2]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n27646), .D(n282[3]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n27646), .D(n282[4]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n27646), .D(n282[5]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n27646), .D(n282[6]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n27646), .D(n282[7]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n27646), .D(n282[8]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n27646), .D(n282[9]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n27646), 
            .D(n282[10]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n27646), 
            .D(n282[11]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n27646), 
            .D(n282[12]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n27646), 
            .D(n282[13]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n27646), 
            .D(n282[14]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n27646), 
            .D(n282[15]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n27646), 
            .D(n282[16]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n27646), 
            .D(n282[17]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n27646), 
            .D(n282[18]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n27646), 
            .D(n282[19]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n27646), 
            .D(n282[20]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n27646), 
            .D(n282[21]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n27646), 
            .D(n282[22]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n27646), 
            .D(n282[23]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n27646), 
            .D(n282[24]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n27646), 
            .D(n282[25]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n27646), 
            .D(n282[26]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n27646), 
            .D(n282[27]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n27646), 
            .D(n282[28]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n27646), 
            .D(n282[29]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n27646), 
            .D(n282[30]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n27646), 
            .D(n282[31]), .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n37470), .O(n282[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28180_4_lut (.I0(n26283), .I1(n43104), .I2(n39092), .I3(state[0]), 
            .O(n43208));
    defparam i28180_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[1] ), 
            .I2(start), .I3(n43208), .O(n7_adj_5134));
    defparam i20_4_lut.LUT_INIT = 16'hcecf;
    SB_LUT4 i1_4_lut (.I0(n26417), .I1(n7_adj_5134), .I2(n34074), .I3(\state[1] ), 
            .O(n41203));
    defparam i1_4_lut.LUT_INIT = 16'hcc8c;
    SB_CARRY add_21_4 (.CI(n37470), .I0(bit_ctr[2]), .I1(GND_net), .CO(n37471));
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n37469), .O(n282[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_3 (.CI(n37469), .I0(bit_ctr[1]), .I1(GND_net), .CO(n37470));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n282[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n37469));
    SB_LUT4 i32307_4_lut (.I0(n39092), .I1(n43104), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n47200));
    defparam i32307_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n46811), .I1(n34008), .I2(\state[1] ), .I3(n26283), 
            .O(n43212));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n43212), .I1(n47201), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n43230));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i3_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(\neo_pixel_transmitter.done_N_742 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_2189_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n38277), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_2189_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n38276), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_32 (.CI(n38276), .I0(GND_net), .I1(timer[30]), 
            .CO(n38277));
    SB_LUT4 timer_2189_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n38275), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_31 (.CI(n38275), .I0(GND_net), .I1(timer[29]), 
            .CO(n38276));
    SB_LUT4 timer_2189_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n38274), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_30 (.CI(n38274), .I0(GND_net), .I1(timer[28]), 
            .CO(n38275));
    SB_LUT4 timer_2189_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n38273), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_29 (.CI(n38273), .I0(GND_net), .I1(timer[27]), 
            .CO(n38274));
    SB_LUT4 timer_2189_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n38272), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_28 (.CI(n38272), .I0(GND_net), .I1(timer[26]), 
            .CO(n38273));
    SB_LUT4 timer_2189_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n38271), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_27 (.CI(n38271), .I0(GND_net), .I1(timer[25]), 
            .CO(n38272));
    SB_LUT4 timer_2189_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n38270), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_26 (.CI(n38270), .I0(GND_net), .I1(timer[24]), 
            .CO(n38271));
    SB_LUT4 timer_2189_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n38269), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_25 (.CI(n38269), .I0(GND_net), .I1(timer[23]), 
            .CO(n38270));
    SB_LUT4 timer_2189_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n38268), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_24 (.CI(n38268), .I0(GND_net), .I1(timer[22]), 
            .CO(n38269));
    SB_LUT4 timer_2189_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n38267), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_23 (.CI(n38267), .I0(GND_net), .I1(timer[21]), 
            .CO(n38268));
    SB_LUT4 timer_2189_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n38266), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_22 (.CI(n38266), .I0(GND_net), .I1(timer[20]), 
            .CO(n38267));
    SB_LUT4 timer_2189_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n38265), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_21 (.CI(n38265), .I0(GND_net), .I1(timer[19]), 
            .CO(n38266));
    SB_LUT4 timer_2189_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n38264), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_20 (.CI(n38264), .I0(GND_net), .I1(timer[18]), 
            .CO(n38265));
    SB_LUT4 timer_2189_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n38263), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_19 (.CI(n38263), .I0(GND_net), .I1(timer[17]), 
            .CO(n38264));
    SB_LUT4 timer_2189_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n38262), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_18 (.CI(n38262), .I0(GND_net), .I1(timer[16]), 
            .CO(n38263));
    SB_LUT4 timer_2189_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n38261), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_17 (.CI(n38261), .I0(GND_net), .I1(timer[15]), 
            .CO(n38262));
    SB_LUT4 timer_2189_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n38260), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_16 (.CI(n38260), .I0(GND_net), .I1(timer[14]), 
            .CO(n38261));
    SB_LUT4 timer_2189_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n38259), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_15 (.CI(n38259), .I0(GND_net), .I1(timer[13]), 
            .CO(n38260));
    SB_LUT4 timer_2189_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n38258), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_14 (.CI(n38258), .I0(GND_net), .I1(timer[12]), 
            .CO(n38259));
    SB_LUT4 timer_2189_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n38257), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_13 (.CI(n38257), .I0(GND_net), .I1(timer[11]), 
            .CO(n38258));
    SB_LUT4 timer_2189_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n38256), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_12 (.CI(n38256), .I0(GND_net), .I1(timer[10]), 
            .CO(n38257));
    SB_LUT4 timer_2189_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n38255), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_11 (.CI(n38255), .I0(GND_net), .I1(timer[9]), 
            .CO(n38256));
    SB_LUT4 timer_2189_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n38254), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_10 (.CI(n38254), .I0(GND_net), .I1(timer[8]), 
            .CO(n38255));
    SB_LUT4 timer_2189_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n38253), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_9 (.CI(n38253), .I0(GND_net), .I1(timer[7]), 
            .CO(n38254));
    SB_LUT4 timer_2189_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n38252), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_8 (.CI(n38252), .I0(GND_net), .I1(timer[6]), 
            .CO(n38253));
    SB_LUT4 timer_2189_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n38251), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_7 (.CI(n38251), .I0(GND_net), .I1(timer[5]), 
            .CO(n38252));
    SB_LUT4 timer_2189_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n38250), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_6 (.CI(n38250), .I0(GND_net), .I1(timer[4]), 
            .CO(n38251));
    SB_LUT4 timer_2189_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n38249), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_5 (.CI(n38249), .I0(GND_net), .I1(timer[3]), 
            .CO(n38250));
    SB_LUT4 timer_2189_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n38248), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_4 (.CI(n38248), .I0(GND_net), .I1(timer[2]), 
            .CO(n38249));
    SB_LUT4 timer_2189_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n38247), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_3 (.CI(n38247), .I0(GND_net), .I1(timer[1]), 
            .CO(n38248));
    SB_LUT4 timer_2189_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_2189_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_2189_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n38247));
    SB_DFF timer_2189__i31 (.Q(timer[31]), .C(CLK_c), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i30 (.Q(timer[30]), .C(CLK_c), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i29 (.Q(timer[29]), .C(CLK_c), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i28 (.Q(timer[28]), .C(CLK_c), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i27 (.Q(timer[27]), .C(CLK_c), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i26 (.Q(timer[26]), .C(CLK_c), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i25 (.Q(timer[25]), .C(CLK_c), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i24 (.Q(timer[24]), .C(CLK_c), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i23 (.Q(timer[23]), .C(CLK_c), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i22 (.Q(timer[22]), .C(CLK_c), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i21 (.Q(timer[21]), .C(CLK_c), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i20 (.Q(timer[20]), .C(CLK_c), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i19 (.Q(timer[19]), .C(CLK_c), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i18 (.Q(timer[18]), .C(CLK_c), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i17 (.Q(timer[17]), .C(CLK_c), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i16 (.Q(timer[16]), .C(CLK_c), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i15 (.Q(timer[15]), .C(CLK_c), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i14 (.Q(timer[14]), .C(CLK_c), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i13 (.Q(timer[13]), .C(CLK_c), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i12 (.Q(timer[12]), .C(CLK_c), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i11 (.Q(timer[11]), .C(CLK_c), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i10 (.Q(timer[10]), .C(CLK_c), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i9 (.Q(timer[9]), .C(CLK_c), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i8 (.Q(timer[8]), .C(CLK_c), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i7 (.Q(timer[7]), .C(CLK_c), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i6 (.Q(timer[6]), .C(CLK_c), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i5 (.Q(timer[5]), .C(CLK_c), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i4 (.Q(timer[4]), .C(CLK_c), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i3 (.Q(timer[3]), .C(CLK_c), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i2 (.Q(timer[2]), .C(CLK_c), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_2189__i1 (.Q(timer[1]), .C(CLK_c), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 n48784_bdd_4_lut (.I0(n48784), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(color_bit_N_722[1]), .O(n48787));
    defparam n48784_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_add_2_33_lut (.I0(n45586), .I1(timer[31]), .I2(n1[31]), 
            .I3(n37657), .O(n26449)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n45584), .I1(timer[30]), .I2(n1[30]), 
            .I3(n37656), .O(n45586)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n37656), .I0(timer[30]), .I1(n1[30]), 
            .CO(n37657));
    SB_LUT4 sub_14_add_2_31_lut (.I0(n45582), .I1(timer[29]), .I2(n1[29]), 
            .I3(n37655), .O(n45584)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n37655), .I0(timer[29]), .I1(n1[29]), 
            .CO(n37656));
    SB_LUT4 sub_14_add_2_30_lut (.I0(n45580), .I1(timer[28]), .I2(n1[28]), 
            .I3(n37654), .O(n45582)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_30 (.CI(n37654), .I0(timer[28]), .I1(n1[28]), 
            .CO(n37655));
    SB_LUT4 sub_14_add_2_29_lut (.I0(n45578), .I1(timer[27]), .I2(n1[27]), 
            .I3(n37653), .O(n45580)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n37653), .I0(timer[27]), .I1(n1[27]), 
            .CO(n37654));
    SB_LUT4 sub_14_add_2_28_lut (.I0(n45576), .I1(timer[26]), .I2(n1[26]), 
            .I3(n37652), .O(n45578)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_28 (.CI(n37652), .I0(timer[26]), .I1(n1[26]), 
            .CO(n37653));
    SB_LUT4 sub_14_add_2_27_lut (.I0(n45574), .I1(timer[25]), .I2(n1[25]), 
            .I3(n37651), .O(n45576)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_27 (.CI(n37651), .I0(timer[25]), .I1(n1[25]), 
            .CO(n37652));
    SB_LUT4 sub_14_add_2_26_lut (.I0(n45572), .I1(timer[24]), .I2(n1[24]), 
            .I3(n37650), .O(n45574)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_26 (.CI(n37650), .I0(timer[24]), .I1(n1[24]), 
            .CO(n37651));
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 n48724_bdd_4_lut (.I0(n48724), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(color_bit_N_722[1]), .O(n48727));
    defparam n48724_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n48712_bdd_4_lut (.I0(n48712), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(color_bit_N_722[1]), .O(n48715));
    defparam n48712_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 n48706_bdd_4_lut (.I0(n48706), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(color_bit_N_722[1]), .O(n48709));
    defparam n48706_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i509_2_lut (.I0(n34008), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1991));   // verilog/neopixel.v(103[9] 111[12])
    defparam i509_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut (.I0(n34074), .I1(n46813), .I2(\state[1] ), .I3(n26417), 
            .O(n43011));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i30837_3_lut (.I0(n48727), .I1(n48715), .I2(color_bit_N_722[2]), 
            .I3(GND_net), .O(n45968));
    defparam i30837_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32318_3_lut (.I0(n48601), .I1(n48709), .I2(color_bit_N_722[2]), 
            .I3(GND_net), .O(n47450));
    defparam i32318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_rep_335_2_lut (.I0(bit_ctr[3]), .I1(n33857), .I2(GND_net), 
            .I3(GND_net), .O(n49107));
    defparam i1_rep_335_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[4]), .I1(bit_ctr[3]), .I2(n33857), .I3(GND_net), 
            .O(n39590));
    defparam i1_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i32396_4_lut (.I0(n47450), .I1(n45968), .I2(bit_ctr[3]), .I3(n33857), 
            .O(n47528));   // verilog/neopixel.v(22[26:38])
    defparam i32396_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i31841_4_lut (.I0(n48619), .I1(n49107), .I2(n48787), .I3(color_bit_N_722[2]), 
            .O(n46833));
    defparam i31841_4_lut.LUT_INIT = 16'hc088;
    SB_LUT4 i19786_4_lut (.I0(n46833), .I1(\state_3__N_528[1] ), .I2(n47528), 
            .I3(n39590), .O(state_3__N_528[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i19786_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_25_lut (.I0(n45570), .I1(timer[23]), .I2(n1[23]), 
            .I3(n37649), .O(n45572)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n37649), .I0(timer[23]), .I1(n1[23]), 
            .CO(n37650));
    SB_LUT4 sub_14_add_2_24_lut (.I0(n45568), .I1(timer[22]), .I2(n1[22]), 
            .I3(n37648), .O(n45570)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n37648), .I0(timer[22]), .I1(n1[22]), 
            .CO(n37649));
    SB_LUT4 sub_14_add_2_23_lut (.I0(n45566), .I1(timer[21]), .I2(n1[21]), 
            .I3(n37647), .O(n45568)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n37647), .I0(timer[21]), .I1(n1[21]), 
            .CO(n37648));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n45564), .I1(timer[20]), .I2(n1[20]), 
            .I3(n37646), .O(n45566)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n37646), .I0(timer[20]), .I1(n1[20]), 
            .CO(n37647));
    SB_LUT4 sub_14_add_2_21_lut (.I0(n45562), .I1(timer[19]), .I2(n1[19]), 
            .I3(n37645), .O(n45564)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_21 (.CI(n37645), .I0(timer[19]), .I1(n1[19]), 
            .CO(n37646));
    SB_LUT4 sub_14_add_2_20_lut (.I0(n45560), .I1(timer[18]), .I2(n1[18]), 
            .I3(n37644), .O(n45562)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_20 (.CI(n37644), .I0(timer[18]), .I1(n1[18]), 
            .CO(n37645));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n45558), .I1(timer[17]), .I2(n1[17]), 
            .I3(n37643), .O(n45560)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n37643), .I0(timer[17]), .I1(n1[17]), 
            .CO(n37644));
    SB_DFFESS state_i0 (.Q(state[0]), .C(CLK_c), .E(n27791), .D(state_3__N_528[0]), 
            .S(n43011));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_18_lut (.I0(n45556), .I1(timer[16]), .I2(n1[16]), 
            .I3(n37642), .O(n45558)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_18 (.CI(n37642), .I0(timer[16]), .I1(n1[16]), 
            .CO(n37643));
    SB_LUT4 sub_14_add_2_17_lut (.I0(n45554), .I1(timer[15]), .I2(n1[15]), 
            .I3(n37641), .O(n45556)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_DFF timer_2189__i0 (.Q(timer[0]), .C(CLK_c), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n27646), .D(n282[0]), 
            .R(n28039));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(color_bit_N_722[1]));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY sub_14_add_2_17 (.CI(n37641), .I0(timer[15]), .I1(n1[15]), 
            .CO(n37642));
    SB_DFFE state_i1 (.Q(\state[1] ), .C(CLK_c), .E(VCC_net), .D(n28195));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n28165));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_16_lut (.I0(n45552), .I1(timer[14]), .I2(n1[14]), 
            .I3(n37640), .O(n45554)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n37640), .I0(timer[14]), .I1(n1[14]), 
            .CO(n37641));
    SB_LUT4 sub_14_add_2_15_lut (.I0(n45550), .I1(timer[13]), .I2(n1[13]), 
            .I3(n37639), .O(n45552)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_15 (.CI(n37639), .I0(timer[13]), .I1(n1[13]), 
            .CO(n37640));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_679[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n37638), .O(n45550)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 n48616_bdd_4_lut (.I0(n48616), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(color_bit_N_722[1]), .O(n48619));
    defparam n48616_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_14 (.CI(n37638), .I0(timer[12]), .I1(n1[12]), 
            .CO(n37639));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n37637), .O(one_wire_N_679[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n37637), .I0(timer[11]), .I1(n1[11]), 
            .CO(n37638));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n37636), .O(one_wire_N_679[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n37636), .I0(timer[10]), .I1(n1[10]), 
            .CO(n37637));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n37635), .O(one_wire_N_679[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n37635), .I0(timer[9]), .I1(n1[9]), 
            .CO(n37636));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n37634), .O(one_wire_N_679[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n37634), .I0(timer[8]), .I1(n1[8]), 
            .CO(n37635));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n37633), .O(one_wire_N_679[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n37633), .I0(timer[7]), .I1(n1[7]), .CO(n37634));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n37632), .O(one_wire_N_679[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n37632), .I0(timer[6]), .I1(n1[6]), .CO(n37633));
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n37499), .O(n282[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n37631), .O(one_wire_N_679[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n37631), .I0(timer[5]), .I1(n1[5]), .CO(n37632));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n37630), .O(one_wire_N_679[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n37498), .O(n282[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n37630), .I0(timer[4]), .I1(n1[4]), .CO(n37631));
    SB_LUT4 i2_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_1560 (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48));
    defparam i20_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n37629), .O(one_wire_N_679[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n37629), .I0(timer[3]), .I1(n1[3]), .CO(n37630));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n37628), .O(one_wire_N_679[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n37628), .I0(timer[2]), .I1(n1[2]), .CO(n37629));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_679[3]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n37627), .O(n43001)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_3 (.CI(n37627), .I0(timer[1]), .I1(n1[1]), .CO(n37628));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n37627));
    SB_CARRY add_21_32 (.CI(n37498), .I0(bit_ctr[30]), .I1(GND_net), .CO(n37499));
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n37497), .O(n282[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_31 (.CI(n37497), .I0(bit_ctr[29]), .I1(GND_net), .CO(n37498));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n37496), .O(n282[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n37496), .I0(bit_ctr[28]), .I1(GND_net), .CO(n37497));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n37495), .O(n282[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n37495), .I0(bit_ctr[27]), .I1(GND_net), .CO(n37496));
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n37494), .O(n282[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_28 (.CI(n37494), .I0(bit_ctr[26]), .I1(GND_net), .CO(n37495));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n37493), .O(n282[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_27 (.CI(n37493), .I0(bit_ctr[25]), .I1(GND_net), .CO(n37494));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n37492), .O(n282[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_26 (.CI(n37492), .I0(bit_ctr[24]), .I1(GND_net), .CO(n37493));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n37491), .O(n282[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_25 (.CI(n37491), .I0(bit_ctr[23]), .I1(GND_net), .CO(n37492));
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n37490), .O(n282[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_24 (.CI(n37490), .I0(bit_ctr[22]), .I1(GND_net), .CO(n37491));
    SB_LUT4 i15_4_lut_adj_1561 (.I0(bit_ctr[3]), .I1(n30), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43));
    defparam i15_4_lut_adj_1561.LUT_INIT = 16'hfefc;
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n37489), .O(n282[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n37489), .I0(bit_ctr[21]), .I1(GND_net), .CO(n37490));
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n37488), .O(n282[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_22 (.CI(n37488), .I0(bit_ctr[20]), .I1(GND_net), .CO(n37489));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n37487), .O(n282[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_528[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n26417));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'hbbbb;
    SB_CARRY add_21_21 (.CI(n37487), .I0(bit_ctr[19]), .I1(GND_net), .CO(n37488));
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n37486), .O(n282[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_20 (.CI(n37486), .I0(bit_ctr[18]), .I1(GND_net), .CO(n37487));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n37485), .O(n282[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_19 (.CI(n37485), .I0(bit_ctr[17]), .I1(GND_net), .CO(n37486));
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n37484), .O(n282[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_18 (.CI(n37484), .I0(bit_ctr[16]), .I1(GND_net), .CO(n37485));
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n37483), .O(n282[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i495_2_lut (.I0(LED_c), .I1(\state_3__N_528[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1977));   // verilog/neopixel.v(40[18] 45[12])
    defparam i495_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_21_17 (.CI(n37483), .I0(bit_ctr[15]), .I1(GND_net), .CO(n37484));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n37482), .O(n282[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_16 (.CI(n37482), .I0(bit_ctr[14]), .I1(GND_net), .CO(n37483));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n37481), .O(n282[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_15 (.CI(n37481), .I0(bit_ctr[13]), .I1(GND_net), .CO(n37482));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n37480), .O(n282[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_14 (.CI(n37480), .I0(bit_ctr[12]), .I1(GND_net), .CO(n37481));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n37479), .O(n282[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_13 (.CI(n37479), .I0(bit_ctr[11]), .I1(GND_net), .CO(n37480));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n37478), .O(n282[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n28649));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n28648));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n28647));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n28646));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n28645));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n28644));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_12 (.CI(n37478), .I0(bit_ctr[10]), .I1(GND_net), .CO(n37479));
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n28643));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n28642));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n28641));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n28640));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n28639));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n28638));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n28637));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n28636));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n28635));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n28634));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n28633));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n28632));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n28631));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n28630));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n28629));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n28628));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n28627));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n28626));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n28625));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n28624));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n28623));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n28622));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n37477), .O(n282[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n28621));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n28620));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n28619));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_11 (.CI(n37477), .I0(bit_ctr[9]), .I1(GND_net), .CO(n37478));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n37476), .O(n282[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4559_4_lut (.I0(n33935), .I1(n1977), .I2(\state[1] ), .I3(n26417), 
            .O(n6921));
    defparam i4559_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i31907_3_lut (.I0(n39092), .I1(n26417), .I2(n26283), .I3(GND_net), 
            .O(n46884));
    defparam i31907_3_lut.LUT_INIT = 16'hcdcd;
    SB_CARRY add_21_10 (.CI(n37476), .I0(bit_ctr[8]), .I1(GND_net), .CO(n37477));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n37475), .O(n282[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_9 (.CI(n37475), .I0(bit_ctr[7]), .I1(GND_net), .CO(n37476));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n37474), .O(n282[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_ctr_0__bdd_4_lut_33477_4_lut_4_lut (.I0(bit_ctr[1]), .I1(bit_ctr[0]), 
            .I2(neopxl_color[13]), .I3(neopxl_color[12]), .O(n48598));   // verilog/neopixel.v(19[6:15])
    defparam bit_ctr_0__bdd_4_lut_33477_4_lut_4_lut.LUT_INIT = 16'hd5c4;
    SB_CARRY add_21_8 (.CI(n37474), .I0(bit_ctr[6]), .I1(GND_net), .CO(n37475));
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n37473), .O(n282[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_7 (.CI(n37473), .I0(bit_ctr[5]), .I1(GND_net), .CO(n37474));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n37472), .O(n282[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_6 (.CI(n37472), .I0(bit_ctr[4]), .I1(GND_net), .CO(n37473));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n43230), .D(\neo_pixel_transmitter.done_N_742 ), 
            .R(n44844));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n37471), .O(n282[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[1] ), .I1(state[0]), .I2(n1991), 
            .I3(n42982), .O(n27791));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hdf8a;
    SB_LUT4 i32702_4_lut_4_lut (.I0(\state[1] ), .I1(state[0]), .I2(n6921), 
            .I3(n46884), .O(n27646));
    defparam i32702_4_lut_4_lut.LUT_INIT = 16'h0c1d;
    SB_LUT4 i2_2_lut_3_lut (.I0(n26283), .I1(one_wire_N_679[3]), .I2(one_wire_N_679[2]), 
            .I3(GND_net), .O(n33935));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut (.I0(state[0]), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_528[1] ), .O(n28039));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 bit_ctr_0__bdd_4_lut_33550_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n48616));
    defparam bit_ctr_0__bdd_4_lut_33550_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i1_2_lut_3_lut_adj_1563 (.I0(n34074), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n42982));
    defparam i1_2_lut_3_lut_adj_1563.LUT_INIT = 16'h2020;
    SB_LUT4 i31771_2_lut_3_lut (.I0(n34008), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n46813));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31771_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 bit_ctr_0__bdd_4_lut_33555_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n48706));
    defparam bit_ctr_0__bdd_4_lut_33555_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_33564_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n48712));
    defparam bit_ctr_0__bdd_4_lut_33564_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_33614_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n48724));
    defparam bit_ctr_0__bdd_4_lut_33614_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 bit_ctr_0__bdd_4_lut_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n48784));
    defparam bit_ctr_0__bdd_4_lut_4_lut.LUT_INIT = 16'heea0;
    SB_LUT4 i20499_4_lut (.I0(one_wire_N_679[8]), .I1(n26449), .I2(one_wire_N_679[10]), 
            .I3(one_wire_N_679[9]), .O(n34008));
    defparam i20499_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i28081_2_lut (.I0(one_wire_N_679[3]), .I1(one_wire_N_679[2]), 
            .I2(GND_net), .I3(GND_net), .O(n43104));
    defparam i28081_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1564 (.I0(one_wire_N_679[2]), .I1(n43001), .I2(GND_net), 
            .I3(GND_net), .O(n39092));
    defparam i2_2_lut_adj_1564.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1565 (.I0(one_wire_N_679[5]), .I1(one_wire_N_679[4]), 
            .I2(GND_net), .I3(GND_net), .O(n45588));   // verilog/neopixel.v(55[15:42])
    defparam i1_2_lut_adj_1565.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1566 (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[7]), 
            .I2(one_wire_N_679[6]), .I3(n45588), .O(n45594));   // verilog/neopixel.v(55[15:42])
    defparam i1_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1567 (.I0(one_wire_N_679[10]), .I1(n26449), .I2(one_wire_N_679[9]), 
            .I3(n45594), .O(n26283));   // verilog/neopixel.v(55[15:42])
    defparam i1_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 i28128_4_lut (.I0(n26283), .I1(n39092), .I2(n43104), .I3(state[0]), 
            .O(n34074));
    defparam i28128_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i31951_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n46823));
    defparam i31951_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i28154_3_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(n34074), .I3(GND_net), .O(n43181));
    defparam i28154_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i15_4_lut_adj_1568 (.I0(n43181), .I1(n46823), .I2(\state[1] ), 
            .I3(n34008), .O(n7));
    defparam i15_4_lut_adj_1568.LUT_INIT = 16'h3a0a;
    SB_LUT4 i33079_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(start_N_727));   // verilog/neopixel.v(36[4] 116[11])
    defparam i33079_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i28077_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n43100));
    defparam i28077_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i32675_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42246));
    defparam i32675_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1569 (.I0(one_wire_N_679[2]), .I1(n42246), .I2(one_wire_N_679[3]), 
            .I3(n43001), .O(n103));
    defparam i1_4_lut_adj_1569.LUT_INIT = 16'h45cd;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_679[7]), .I1(one_wire_N_679[9]), .I2(n43100), 
            .I3(n103), .O(n16_adj_5136));
    defparam i6_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1570 (.I0(one_wire_N_679[8]), .I1(one_wire_N_679[4]), 
            .I2(n16_adj_5136), .I3(n26449), .O(n6_adj_5137));
    defparam i1_4_lut_adj_1570.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_679[10]), .I1(one_wire_N_679[6]), .I2(one_wire_N_679[5]), 
            .I3(n6_adj_5137), .O(n48855));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1255_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_736 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_1255_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i32069_3_lut_4_lut (.I0(n26283), .I1(n47200), .I2(start), 
            .I3(\state[1] ), .O(n47201));
    defparam i32069_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31953_2_lut_3_lut (.I0(one_wire_N_679[3]), .I1(one_wire_N_679[2]), 
            .I2(start), .I3(GND_net), .O(n46811));
    defparam i31953_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n34008), .I1(\state[1] ), .I2(state[0]), 
            .I3(\neo_pixel_transmitter.done ), .O(n44844));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 n48598_bdd_4_lut_4_lut (.I0(color_bit_N_722[1]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(n48598), .O(n48601));   // verilog/neopixel.v(19[6:15])
    defparam n48598_bdd_4_lut_4_lut.LUT_INIT = 16'hf588;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=52, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Ki[15] , GND_net, PWMLimit, \Kp[6] , \Kp[1] , 
            \Kp[0] , \Kp[2] , \Kp[3] , \Kp[4] , \Kp[5] , \Kp[7] , 
            \Kp[8] , \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , 
            \Kp[14] , \Kp[15] , \Ki[1] , \Ki[0] , \Ki[2] , \Ki[3] , 
            \Ki[4] , \Ki[10] , \Ki[5] , \Ki[6] , \Ki[7] , \Ki[8] , 
            \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , IntegralLimit, 
            \Ki[9] , setpoint, motor_state, duty, clk32MHz, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input \Ki[15] ;
    input GND_net;
    input [23:0]PWMLimit;
    input \Kp[6] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[10] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input [23:0]IntegralLimit;
    input \Ki[9] ;
    input [23:0]setpoint;
    input [23:0]motor_state;
    output [23:0]duty;
    input clk32MHz;
    input VCC_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]\PID_CONTROLLER.integral_23__N_3672 ;
    
    wire n1117, n38548;
    wire [15:0]n15425;
    
    wire n749, n38549;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    wire [23:0]n4236;
    
    wire n37591;
    wire [23:0]n1;
    wire [23:0]n28;
    
    wire n487, n95, n26, n37592, n168, n241, n314, n387, n460, 
        n533, n560, n606, n679, n752, n825, n898, n37590, n971, 
        n1044;
    wire [16:0]n14813;
    
    wire n676, n38547, n1117_adj_4709, n119, n50, n192, n265, 
        n338, n101, n32, n174, n755, n411, n484, n557, n630, 
        n92, n828, n23, n165, n238;
    wire [23:0]duty_23__N_3772;
    
    wire n47011, n247, n311, n901, n384, n457, n530, n603, n974, 
        n676_adj_4710, n749_adj_4711, n822, n895, n968, n1041, n1114, 
        n6, n89, n20_adj_4712, n162;
    wire [10:0]n17545;
    wire [9:0]n17809;
    
    wire n840, n38425, n235, n308, n381, n454, n527, n600;
    wire [47:0]n155;
    wire [47:0]n106;
    
    wire n673, n746, n819, n892, n965, n1047, n1038, n1111, 
        n92_adj_4714, n23_adj_4715, n47311, n47520, n48879, n47101, 
        n47698, n320, \PID_CONTROLLER.integral_23__N_3720 , n393, n466, 
        n116, n165_adj_4717, n47, n189, n47759, n47319, n1120, 
        n262, n335, n119_adj_4719, n767, n38424, n694, n38423, 
        n621, n38422, n47702;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3723 ;
    
    wire \PID_CONTROLLER.integral_23__N_3722 , n408, n50_adj_4720, n548, 
        n38421, n475, n38420, n481, n554, n627, n700, n86, n17, 
        n159, n192_adj_4721, n232, n305, n378, n451, n603_adj_4722, 
        n38546, n402, n38419, n524, n329, n38418, n597, n670, 
        n743, n816, n889, n962, n1035, n1108, n539, n83, n256, 
        n38417, n37589, n14, n156, n229, n302, n530_adj_4724, 
        n38545, n183, n38416, n41, n110, n375, n448, n521, n594, 
        n47103, n47750, n667, n740, n813, n886, n959, n1032, 
        n1105, n80, n11_adj_4725, n153, n226, n299, n372, n445, 
        n518, n457_adj_4726, n38544, n591, n664, n737, n810, n883, 
        n956, n1029, n1102, n384_adj_4727, n38543, n612, n113, 
        n44, n265_adj_4728, n186, n259;
    wire [23:0]n257;
    
    wire n256_adj_4729;
    wire [23:0]duty_23__N_3747;
    
    wire n332, duty_23__N_3771;
    wire [23:0]duty_23__N_3648;
    
    wire n405, n478, n311_adj_4730, n38542, n77, n8_adj_4734, n150, 
        n223, n296, n369, n442, n37676, n37677, n238_adj_4736, 
        n38541, n37675, n38540, n515, n37674, n588, n661, n37673, 
        n734, n807, n37672, n880, n37671, n37670, n953, n47133, 
        n1026, n1099, n37669, n11_adj_4740, n9_adj_4741, n47131, 
        n37668;
    wire [14:0]n15969;
    
    wire n38539, n38538, n48927, n47570, n17_adj_4742, n47384, n48909, 
        n47382, n1044_adj_4743, n38537, n822_adj_4744, n895_adj_4745, 
        n968_adj_4746, n47380, n971_adj_4747, n38536, n1041_adj_4748, 
        n37667, n898_adj_4749, n38535;
    wire [0:0]n10614;
    wire [0:0]n10083;
    
    wire n37588, n37587, n48903, n1114_adj_4750, n825_adj_4751, n38534, 
        n37586, n37666, n752_adj_4753, n38533, n679_adj_4754, n38532, 
        n116_adj_4755, n27, n15_adj_4756, n13_adj_4757, n11_adj_4758, 
        n47071, n47_adj_4759, n606_adj_4760, n38531, n37585, n533_adj_4762, 
        n38530, n37665, n460_adj_4763, n38529, n387_adj_4764, n38528, 
        n189_adj_4765, n262_adj_4766, n37664, n37584, n335_adj_4767, 
        n408_adj_4768, n481_adj_4769, n314_adj_4770, n38527, n241_adj_4771, 
        n38526, n37583, n21_adj_4772, n19_adj_4773, n17_adj_4774, 
        n9_adj_4775, n47080, n37663, n37582, n37662;
    wire [23:0]n1_adj_5132;
    
    wire n168_adj_4778, n38525, n551, n43, n16_adj_4779, n37661, 
        n26_adj_4781, n95_adj_4782, n37660, n37581;
    wire [7:0]n18289;
    wire [6:0]n18416;
    
    wire n630_adj_4783, n38524, n554_adj_4784, n47013, n8_adj_4785, 
        n74, n5_adj_4786, n147, n220, n293, n366, n439, n624, 
        n512, n585, n658, n731, n804, n877, n557_adj_4787, n38523, 
        n950, n37659;
    wire [8:0]n18029;
    
    wire n770, n37758, n1023, n697, n37757, n484_adj_4789, n38522, 
        n37658, n1096, n411_adj_4790, n38521, n37580, n45, n24_adj_4791, 
        n7_adj_4792, n5_adj_4793, n47097, n37756, n47356, n37755, 
        n47352, n25_adj_4794, n23_adj_4795, n47720, n31, n29, n47536, 
        n37, n35, n33, n47752, n338_adj_4796, n38520, n37754, 
        n37753, n47386, n37752, n48896, n37751, n37750, n47374, 
        n48891, n12_adj_4797, n47109, n48914, n10_adj_4798, n30, 
        n47654, n37579, n38519, n39, n41_adj_4800, n37578, n45_adj_4801, 
        n43_adj_4802, n29_adj_4803, n31_adj_4804, n37577, n37_adj_4805, 
        n23_adj_4806, n25_adj_4807, n37576, n35_adj_4809, n38518, 
        n47117, n11_adj_4811, n13_adj_4812, n15_adj_4813, n27_adj_4814, 
        n33_adj_4815, n9_adj_4816, n17_adj_4817, n37575, n19_adj_4818, 
        n627_adj_4819, n37574, n37573;
    wire [13:0]n16449;
    
    wire n38517, n21_adj_4820, n46988, n46982, n12_adj_4821, n48894, 
        n38516, n37572, n10_adj_4823, n30_adj_4824, n37571, n47302, 
        n47562, n48920, n47724, n48885, n38515, n37570, n47780, 
        n47286, n47690, n48882, n47490, n16_adj_4826, n37569, n38514, 
        n47746, n38513, n47099, n16_adj_4828, n47696, n47697, n685, 
        n38512, n8_adj_4830, n24_adj_4831, n24_adj_4832, n6_adj_4833, 
        n47646, n47647, n46965, n46962, n47524, n47617, n700_adj_4834, 
        n89_adj_4836, n4_adj_4837, n20_adj_4838, n47662, n162_adj_4839, 
        n47663, n46977, n46975, n47762, n235_adj_4840, n47619, n47802, 
        n47803, n47791, n8_adj_4841, n308_adj_4842, n46967, n47706, 
        n40, n47708, n381_adj_4843, n41_adj_4844, n682, n38511, 
        n39_adj_4845, n454_adj_4846, n609, n38510, n45_adj_4847, n536, 
        n38509, n463, n38508, n390, n38507, n37568, n317, n38506, 
        n244, n38505, n171, n38504, n29_adj_4848, n98;
    wire [12:0]n16869;
    
    wire n1050, n38503, n977, n38502, n527_adj_4849, n904, n38501, 
        n831, n38500, n3_adj_4850, n4_adj_4851, n758, n38499, n47554, 
        n600_adj_4852, n673_adj_4853, n43_adj_4854, n746_adj_4855, n37_adj_4856, 
        n29_adj_4857, n31_adj_4858;
    wire [21:0]n11121;
    
    wire n38923, n38922, n819_adj_4860, n38921, n38920, n38919, 
        n38918, n38917, n37567, n892_adj_4861, n38498, n38916, n37726, 
        n965_adj_4862, n1038_adj_4863, n47555, n23_adj_4864, n25_adj_4865, 
        n35_adj_4866, n12_adj_4867, n38915, n38914, n33_adj_4868, 
        n11_adj_4869, n38913, n38912, n38911, n38910, n38909, n38908, 
        n38907, n13_adj_4870, n15_adj_4871, n38906, n38905, n38904, 
        n38903, n38902;
    wire [20:0]n12088;
    
    wire n38901, n38900, n27_adj_4873, n9_adj_4874, n17_adj_4875, 
        n19_adj_4876, n21_adj_4877, n46947, n47065, n10_adj_4878, 
        n46941, n12_adj_4879, n30_adj_4880, n47067, n10_adj_4881, 
        n30_adj_4882, n46960, n47242, n47238, n47682, n47470, n1111_adj_4883, 
        n38899, n38898, n38897, n38896, n38895, n37566, n38894, 
        n37725, n38893, n38892, n38891, n38890, n38889, n38888, 
        n38887, n38886, n47744, n16_adj_4884, n6_adj_4885, n47678, 
        n38885, n38884, n38883, n38882, n38881;
    wire [19:0]n12969;
    
    wire n38880, n38879, n38878, n38877, n38876, n37724, n47670, 
        n47679, n86_adj_4886, n17_adj_4887, n8_adj_4888, n24_adj_4889, 
        n46922, n46920, n47526, n47623, n159_adj_4890, n232_adj_4891, 
        n4_adj_4892, n38497, n305_adj_4893, n38875, n38874, n38873, 
        n47323, n38872, n38871, n47778, n38870, n38869, n38868, 
        n38867, n38866, n38865, n38864, n38863, n38862, n378_adj_4894, 
        n47676, n47677, n38861, n46937;
    wire [18:0]n13768;
    
    wire n38860, n38859, n38858, n38857, n38856, n46935, n47764, 
        n38855, n38854, n38853, n38852, n38851, n38850, n38849, 
        n37723, n47779, n451_adj_4895, n524_adj_4896, n597_adj_4897, 
        n38848, n38847, n38846, n38845, n38844, n38843, n38842;
    wire [17:0]n14489;
    
    wire n38841, n38840, n38839, n38496, n38838, n38837, n47625, 
        n38836, n47804, n38835, n47805, n38834, n38833, n670_adj_4898, 
        n47789, n38832, n38831, n38830, n38829, n38828, n46924, 
        n743_adj_4899, n47712, n38827, n40_adj_4900, n38826, n47714, 
        n38825, n38824, n816_adj_4901, n889_adj_4902;
    wire [7:0]n18209;
    
    wire n38823, n38822, n39_adj_4903, n47757, n38821, n38820, n6_adj_4904, 
        n47556, n38819, n47557, n38818, n47015, n38817, n38816, 
        n47522, n47321, n41_adj_4905, n47025, n38495, n47700, n38494, 
        n37722;
    wire [16:0]n15136;
    
    wire n38815, n47329, n38493, n38814, n38813, n38812, n38811, 
        n38810, n38809, n38808, n38807, n38806, n38805, n962_adj_4907, 
        n38804, n38803, n38802, n38801, n38800, n38799;
    wire [15:0]n15713;
    
    wire n38798, n38797, n38796, n38795, n38794, n38793, n4_adj_4908, 
        n38792, n38791, n38790, n1035_adj_4909, n38789, n38788, 
        n38787, n1108_adj_4910, n38786, n38785, n38492, n37160;
    wire [1:0]n18673;
    
    wire n4_adj_4911;
    wire [2:0]n18649;
    
    wire n37721, n4_adj_4912;
    wire [3:0]n18609;
    
    wire n6_adj_4913, n38784, n38783;
    wire [4:0]n18549;
    
    wire n37242;
    wire [6:0]n18353;
    
    wire n38782, n38781, n38780, n38779, n38491, n47564, n38778, 
        n38777, n47565, n113_adj_4914, n44_adj_4915, n47111, n62, 
        n131, n204, n38776, n4_adj_4916, n47668, n47313;
    wire [14:0]n16224;
    
    wire n38775, n38774, n38773, n38772, n38771, n38770, n38769, 
        n4_adj_4917;
    wire [3:0]n18633;
    
    wire n6_adj_4918, n37720, n38768, n38767;
    wire [5:0]n18513;
    
    wire n38490, n38766, n38765, n38764, n37719, n38763;
    wire [4:0]n18584;
    
    wire n38762, n38761, n37718, n38489, n37717, n37716;
    wire [13:0]n16673;
    
    wire n1120_adj_4920, n38760, n37715, n414, n38488, n37714, n1047_adj_4923, 
        n38759, n341, n38487, n37374, n974_adj_4924, n38758, n37713, 
        n901_adj_4926, n38757, n828_adj_4927, n38756, n755_adj_4928, 
        n38755, n682_adj_4929, n38754, n268_adj_4930, n38486, n186_adj_4931, 
        n259_adj_4932, n37292;
    wire [1:0]n18681;
    
    wire n4_adj_4934;
    wire [2:0]n18664;
    
    wire n609_adj_4935, n38753, n536_adj_4936, n38752, n332_adj_4937, 
        n463_adj_4938, n38751, n390_adj_4939, n38750, n62_adj_4940, 
        n131_adj_4941, n204_adj_4942, n317_adj_4943, n38749, n244_adj_4944, 
        n38748, n171_adj_4946, n38747, n405_adj_4947, n29_adj_4948, 
        n98_adj_4949, n478_adj_4950, n551_adj_4951;
    wire [5:0]n18465;
    
    wire n560_adj_4952, n38746, n624_adj_4953, n697_adj_4954, n195_adj_4955, 
        n38485, n487_adj_4956, n38745, n414_adj_4957, n38744, n341_adj_4958, 
        n38743, n53, n122, n268_adj_4959, n38742;
    wire [11:0]n17233;
    
    wire n980, n38484, n195_adj_4960, n38741, n907, n38483, n53_adj_4961, 
        n122_adj_4962;
    wire [12:0]n17064;
    
    wire n1050_adj_4963, n38740, n977_adj_4964, n38739, n904_adj_4965, 
        n38738, n831_adj_4966, n38737, n758_adj_4967, n38736, n770_adj_4968, 
        n685_adj_4969, n38735, n612_adj_4970, n38734, n539_adj_4971, 
        n38733, n466_adj_4972, n38732, n393_adj_4973, n38731, n320_adj_4974, 
        n38730, n247_adj_4975, n38729, n174_adj_4976, n38728, n32_adj_4977, 
        n101_adj_4978;
    wire [11:0]n17401;
    
    wire n980_adj_4979, n38727, n834, n38482, n907_adj_4980, n38726, 
        n834_adj_4981, n38725, n761, n38724, n37712, n761_adj_4983, 
        n38481, n688, n38480, n615, n38479, n688_adj_4985, n38723, 
        n37711, n615_adj_4987, n38722, n47766, n4_adj_4988, n83_adj_4989, 
        n542, n38478, n469, n38477, n396, n38476, n37710, n14_adj_4991, 
        n542_adj_4992, n38721, n469_adj_4993, n38720, n323, n38475, 
        n396_adj_4994, n38719, n323_adj_4995, n38718, n250, n38474, 
        n250_adj_4996, n38717, n177, n38473, n35_adj_4997, n104, 
        n177_adj_4999, n38716, n35_adj_5000, n104_adj_5001, n910, 
        n38472, n43796, n490, n38715, n837, n38471, n417, n38714, 
        n344, n38713, n156_adj_5002, n271_adj_5003, n38712, n198_adj_5004, 
        n38711, n764, n38470, n691, n38469, n618, n38468, n37709, 
        n56, n125, n545, n38467;
    wire [10:0]n17688;
    
    wire n910_adj_5006, n38710, n837_adj_5007, n38709, n472, n38466, 
        n399, n38465, n37708, n326, n38464, n253, n38463, n180, 
        n38462, n37707, n38, n107, n764_adj_5010, n38708, n691_adj_5011, 
        n38707, n44030, n490_adj_5012, n38461, n618_adj_5013, n38706, 
        n417_adj_5014, n38460, n545_adj_5015, n38705, n472_adj_5016, 
        n38704, n399_adj_5017, n38703, n326_adj_5018, n38702, n253_adj_5019, 
        n38701, n180_adj_5020, n38700, n38_adj_5021, n107_adj_5022;
    wire [9:0]n17929;
    
    wire n840_adj_5023, n38699, n37706, n37705, n767_adj_5026, n38698, 
        n344_adj_5027, n38459, n229_adj_5028, n694_adj_5029, n38697, 
        n37704, n621_adj_5031, n38696, n548_adj_5032, n38695, n475_adj_5033, 
        n38694, n402_adj_5034, n38693, n329_adj_5035, n38692, n256_adj_5036, 
        n38691, n183_adj_5037, n38690, n41_adj_5038, n110_adj_5039;
    wire [21:0]n10590;
    
    wire n38689, n38688, n38687, n38686, n37703, n37702, n38685, 
        n38684, n271_adj_5043, n38458, n38683, n198_adj_5044, n38457, 
        n38682, n1096_adj_5045, n38681, n1023_adj_5046, n38680, n950_adj_5047, 
        n38679, n56_adj_5048, n125_adj_5049, n877_adj_5050, n38678, 
        n804_adj_5051, n38677, n731_adj_5052, n38676, n658_adj_5053, 
        n38675, n585_adj_5054, n38674, n512_adj_5055, n38673, n439_adj_5056, 
        n38672, n366_adj_5057, n38671, n293_adj_5058, n38670, n220_adj_5059, 
        n38669, n147_adj_5060, n38668, n5_adj_5061, n74_adj_5062;
    wire [20:0]n11605;
    
    wire n38667, n38666, n37701, n38665, n38664, n38663, n38662, 
        n38661, n1099_adj_5064, n38660, n1026_adj_5065, n38659, n953_adj_5066, 
        n38658, n880_adj_5067, n38657, n807_adj_5068, n38656, n734_adj_5069, 
        n38655, n661_adj_5070, n38654, n588_adj_5071, n38653, n515_adj_5072, 
        n38652, n442_adj_5073, n38651, n369_adj_5074, n38650, n296_adj_5075, 
        n38649, n37700, n223_adj_5077, n38648, n150_adj_5078, n38647, 
        n8_adj_5079, n77_adj_5080, n37699;
    wire [19:0]n12529;
    
    wire n38646, n38645, n37698, n37697, n38644, n37696, n38643, 
        n38642, n38641, n1102_adj_5085, n38640, n37695, n1029_adj_5087, 
        n38639, n956_adj_5088, n38638, n883_adj_5089, n38637, n810_adj_5090, 
        n38636, n737_adj_5091, n38635, n664_adj_5092, n38634, n591_adj_5093, 
        n38633, n518_adj_5094, n38632, n445_adj_5095, n38631, n37694, 
        n372_adj_5097, n38630, n37611, n37693, n37610, n299_adj_5099, 
        n38629, n226_adj_5100, n38628, n153_adj_5101, n38627, n11_adj_5102, 
        n80_adj_5103;
    wire [18:0]n13369;
    
    wire n38626, n38625, n37692, n37609, n37691, n37608, n38624, 
        n38623, n38622, n1105_adj_5106, n38621, n1032_adj_5107, n38620, 
        n959_adj_5108, n38619, n886_adj_5109, n38618, n813_adj_5110, 
        n38617, n740_adj_5111, n38616, n667_adj_5112, n38615, n37607, 
        n37690, n594_adj_5114, n38614, n521_adj_5115, n38613, n448_adj_5116, 
        n38612, n375_adj_5117, n38611, n302_adj_5118, n38610, n38609, 
        n38608, n37606, n37689;
    wire [8:0]n18128;
    
    wire n38607, n38606, n38605, n38604, n38603, n38602, n37688, 
        n38601, n38600, n38599;
    wire [17:0]n14129;
    
    wire n38598, n38597, n38596, n38595, n38594, n38593, n38592, 
        n37605, n37687, n37604, n37603, n38591, n38590, n38589, 
        n38588, n38587, n38586, n38585, n38584, n38583, n38582, 
        n38581, n38580, n38579, n38578, n38577, n47767, n38576, 
        n38575, n38574, n38573, n38572, n38571, n38570, n38569, 
        n38568, n38567, n38566, n38565, n38564, n37602, n37686, 
        n38563, n37685, n37684, n38562, n37683, n37601, n37600, 
        n37682, n37599, n37598, n38561, n37597, n37681, n37596, 
        n37595, n37594, n38560, n38559, n38558, n38557, n38556, 
        n37593, n37680, n38555, n38554, n37679, n38553, n37678, 
        n38552, n38551, n38550, n12_adj_5120, n8_adj_5121, n11_adj_5122, 
        n6_adj_5123, n37185, n18_adj_5124, n13_adj_5125, n12_adj_5126, 
        n8_adj_5127, n11_adj_5128, n6_adj_5129, n37358, n18_adj_5130, 
        n13_adj_5131;
    
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_11 (.CI(n38548), .I0(n15425[8]), .I1(n749), .CO(n38549));
    SB_LUT4 add_958_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n4236[3]), .I3(n37591), .O(\PID_CONTROLLER.integral_23__N_3672 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_958_5 (.CI(n37591), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n4236[3]), .CO(n37592));
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_958_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n4236[2]), .I3(n37590), .O(\PID_CONTROLLER.integral_23__N_3672 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5019_10_lut (.I0(GND_net), .I1(n15425[7]), .I2(n676), 
            .I3(n38547), .O(n14813[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4709));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31880_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(PWMLimit[2]), .O(n47011));   // verilog/motorControl.v(36[10:25])
    defparam i31880_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4710));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4711));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3772[3]), 
            .I2(duty_23__N_3772[2]), .I3(GND_net), .O(n6));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4712));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_10 (.CI(n38547), .I0(n15425[7]), .I1(n676), .CO(n38548));
    SB_LUT4 add_5187_12_lut (.I0(GND_net), .I1(n17809[9]), .I2(n840), 
            .I3(n38425), .O(n17545[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4714));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4715));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32566_4_lut (.I0(n47311), .I1(n47520), .I2(n48879), .I3(n47101), 
            .O(n47698));   // verilog/motorControl.v(31[10:34])
    defparam i32566_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19752_2_lut (.I0(n28[0]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19752_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4717));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32187_3_lut (.I0(n47759), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n47319));   // verilog/motorControl.v(31[10:34])
    defparam i32187_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4719));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5187_11_lut (.I0(GND_net), .I1(n17809[8]), .I2(n767), 
            .I3(n38424), .O(n17545[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5187_11 (.CI(n38424), .I0(n17809[8]), .I1(n767), .CO(n38425));
    SB_LUT4 add_5187_10_lut (.I0(GND_net), .I1(n17809[7]), .I2(n694), 
            .I3(n38423), .O(n17545[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5187_10 (.CI(n38423), .I0(n17809[7]), .I1(n694), .CO(n38424));
    SB_LUT4 add_5187_9_lut (.I0(GND_net), .I1(n17809[6]), .I2(n621), .I3(n38422), 
            .O(n17545[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32571_3_lut (.I0(n47702), .I1(\PID_CONTROLLER.integral_23__N_3723 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3722 ));   // verilog/motorControl.v(31[38:63])
    defparam i32571_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4720));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5187_9 (.CI(n38422), .I0(n17809[6]), .I1(n621), .CO(n38423));
    SB_LUT4 add_5187_8_lut (.I0(GND_net), .I1(n17809[5]), .I2(n548), .I3(n38421), 
            .O(n17545[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5187_8 (.CI(n38421), .I0(n17809[5]), .I1(n548), .CO(n38422));
    SB_LUT4 add_5187_7_lut (.I0(GND_net), .I1(n17809[4]), .I2(n475), .I3(n38420), 
            .O(n17545[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4721));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5187_7 (.CI(n38420), .I0(n17809[4]), .I1(n475), .CO(n38421));
    SB_LUT4 add_5019_9_lut (.I0(GND_net), .I1(n15425[6]), .I2(n603_adj_4722), 
            .I3(n38546), .O(n14813[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5187_6_lut (.I0(GND_net), .I1(n17809[3]), .I2(n402), .I3(n38419), 
            .O(n17545[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5187_6 (.CI(n38419), .I0(n17809[3]), .I1(n402), .CO(n38420));
    SB_LUT4 add_5187_5_lut (.I0(GND_net), .I1(n17809[2]), .I2(n329), .I3(n38418), 
            .O(n17545[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5187_5 (.CI(n38418), .I0(n17809[2]), .I1(n329), .CO(n38419));
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5187_4_lut (.I0(GND_net), .I1(n17809[1]), .I2(n256), .I3(n38417), 
            .O(n17545[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5187_4 (.CI(n38417), .I0(n17809[1]), .I1(n256), .CO(n38418));
    SB_CARRY add_958_4 (.CI(n37590), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n4236[2]), .CO(n37591));
    SB_LUT4 add_958_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n4236[1]), .I3(n37589), .O(\PID_CONTROLLER.integral_23__N_3672 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_9 (.CI(n38546), .I0(n15425[6]), .I1(n603_adj_4722), 
            .CO(n38547));
    SB_LUT4 add_5019_8_lut (.I0(GND_net), .I1(n15425[5]), .I2(n530_adj_4724), 
            .I3(n38545), .O(n14813[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5187_3_lut (.I0(GND_net), .I1(n17809[0]), .I2(n183), .I3(n38416), 
            .O(n17545[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5187_3 (.CI(n38416), .I0(n17809[0]), .I1(n183), .CO(n38417));
    SB_LUT4 add_5187_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n17545[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5187_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5187_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n38416));
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32618_4_lut (.I0(n47319), .I1(n47698), .I2(n48879), .I3(n47103), 
            .O(n47750));   // verilog/motorControl.v(31[10:34])
    defparam i32618_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4725));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_958_3 (.CI(n37589), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n4236[1]), .CO(n37590));
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_8 (.CI(n38545), .I0(n15425[5]), .I1(n530_adj_4724), 
            .CO(n38546));
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5019_7_lut (.I0(GND_net), .I1(n15425[4]), .I2(n457_adj_4726), 
            .I3(n38544), .O(n14813[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_7 (.CI(n38544), .I0(n15425[4]), .I1(n457_adj_4726), 
            .CO(n38545));
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5019_6_lut (.I0(GND_net), .I1(n15425[3]), .I2(n384_adj_4727), 
            .I3(n38543), .O(n14813[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4728));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_6 (.CI(n38543), .I0(n15425[3]), .I1(n384_adj_4727), 
            .CO(n38544));
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3772[1]), .I1(n257[1]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3747[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3772[2]), .I1(n257[2]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3747[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3747[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3747[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5019_5_lut (.I0(GND_net), .I1(n15425[2]), .I2(n311_adj_4730), 
            .I3(n38542), .O(n14813[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3747[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3747[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3747[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3747[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3747[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3747[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5019_5 (.CI(n38542), .I0(n15425[2]), .I1(n311_adj_4730), 
            .CO(n38543));
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3747[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3747[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3747[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3747[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3747[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3747[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3747[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3747[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3747[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3747[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3747[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3747[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3772[23]), .I1(n257[23]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3747[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_850_4_lut  (.I0(n47750), .I1(\PID_CONTROLLER.integral_23__N_3722 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3720 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_850_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n37676), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n37676), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n37677));
    SB_LUT4 add_5019_4_lut (.I0(GND_net), .I1(n15425[1]), .I2(n238_adj_4736), 
            .I3(n38541), .O(n14813[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3648[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5019_4 (.CI(n38541), .I0(n15425[1]), .I1(n238_adj_4736), 
            .CO(n38542));
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n37675), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_3_lut (.I0(GND_net), .I1(n15425[0]), .I2(n165_adj_4717), 
            .I3(n38540), .O(n14813[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n37675), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n37676));
    SB_LUT4 add_958_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n4236[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3672 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_3 (.CI(n38540), .I0(n15425[0]), .I1(n165_adj_4717), 
            .CO(n38541));
    SB_LUT4 add_5019_2_lut (.I0(GND_net), .I1(n23_adj_4715), .I2(n92_adj_4714), 
            .I3(GND_net), .O(n14813[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n37674), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_19 (.CI(n37674), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n37675));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n37673), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n37673), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n37674));
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n37672), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_17 (.CI(n37672), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n37673));
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n37671), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n37671), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n37672));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n37670), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32002_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n47133));
    defparam i32002_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_2 (.CI(GND_net), .I0(n23_adj_4715), .I1(n92_adj_4714), 
            .CO(n38540));
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_15 (.CI(n37670), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n37671));
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n37669), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_14 (.CI(n37669), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n37670));
    SB_LUT4 i32000_3_lut (.I0(n11_adj_4740), .I1(n9_adj_4741), .I2(n47133), 
            .I3(GND_net), .O(n47131));
    defparam i32000_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n37668), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n4236[0]), .CO(n37589));
    SB_LUT4 add_5052_17_lut (.I0(GND_net), .I1(n15969[14]), .I2(GND_net), 
            .I3(n38539), .O(n15425[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5052_16_lut (.I0(GND_net), .I1(n15969[13]), .I2(n1117), 
            .I3(n38538), .O(n15425[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_16 (.CI(n38538), .I0(n15969[13]), .I1(n1117), .CO(n38539));
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_155_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n48927));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_155_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32438_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n48927), 
            .I2(IntegralLimit[7]), .I3(n47131), .O(n47570));
    defparam i32438_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32252_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4742), 
            .I2(IntegralLimit[9]), .I3(n47570), .O(n47384));
    defparam i32252_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_137_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n48909));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_137_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32250_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4742), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4741), .O(n47382));
    defparam i32250_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4741));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4740));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4742));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5052_15_lut (.I0(GND_net), .I1(n15969[12]), .I2(n1044_adj_4743), 
            .I3(n38537), .O(n15425[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4744));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_13 (.CI(n37668), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n37669));
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4745));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4746));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32248_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n48909), 
            .I2(IntegralLimit[11]), .I3(n47382), .O(n47380));
    defparam i32248_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_5052_15 (.CI(n38537), .I0(n15969[12]), .I1(n1044_adj_4743), 
            .CO(n38538));
    SB_LUT4 add_5052_14_lut (.I0(GND_net), .I1(n15969[11]), .I2(n971_adj_4747), 
            .I3(n38536), .O(n15425[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4748));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5052_14 (.CI(n38536), .I0(n15969[11]), .I1(n971_adj_4747), 
            .CO(n38537));
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n37667), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_12 (.CI(n37667), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n37668));
    SB_LUT4 i20012_2_lut (.I0(n28[4]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20012_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5052_13_lut (.I0(GND_net), .I1(n15969[10]), .I2(n898_adj_4749), 
            .I3(n38535), .O(n15425[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n10614[0]), .I2(n10083[0]), 
            .I3(n37588), .O(duty_23__N_3772[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_13 (.CI(n38535), .I0(n15969[10]), .I1(n898_adj_4749), 
            .CO(n38536));
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n37587), .O(duty_23__N_3772[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_24 (.CI(n37587), .I0(n106[22]), .I1(n155[22]), .CO(n37588));
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_131_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n48903));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_131_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4750));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5052_12_lut (.I0(GND_net), .I1(n15969[9]), .I2(n825_adj_4751), 
            .I3(n38534), .O(n15425[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n37586), .O(duty_23__N_3772[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n37666), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_12 (.CI(n38534), .I0(n15969[9]), .I1(n825_adj_4751), 
            .CO(n38535));
    SB_LUT4 add_5052_11_lut (.I0(GND_net), .I1(n15969[8]), .I2(n752_adj_4753), 
            .I3(n38533), .O(n15425[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_11 (.CI(n38533), .I0(n15969[8]), .I1(n752_adj_4753), 
            .CO(n38534));
    SB_LUT4 add_5052_10_lut (.I0(GND_net), .I1(n15969[7]), .I2(n679_adj_4754), 
            .I3(n38532), .O(n15425[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_10 (.CI(n38532), .I0(n15969[7]), .I1(n679_adj_4754), 
            .CO(n38533));
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4755));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31940_4_lut (.I0(n27), .I1(n15_adj_4756), .I2(n13_adj_4757), 
            .I3(n11_adj_4758), .O(n47071));
    defparam i31940_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4759));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_23 (.CI(n37586), .I0(n106[21]), .I1(n155[21]), .CO(n37587));
    SB_LUT4 add_5052_9_lut (.I0(GND_net), .I1(n15969[6]), .I2(n606_adj_4760), 
            .I3(n38531), .O(n15425[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_9 (.CI(n38531), .I0(n15969[6]), .I1(n606_adj_4760), 
            .CO(n38532));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n37585), .O(duty_23__N_3772[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5052_8_lut (.I0(GND_net), .I1(n15969[5]), .I2(n533_adj_4762), 
            .I3(n38530), .O(n15425[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_11 (.CI(n37666), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n37667));
    SB_LUT4 i20011_2_lut (.I0(n28[5]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20011_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_22 (.CI(n37585), .I0(n106[20]), .I1(n155[20]), .CO(n37586));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n37665), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_8 (.CI(n38530), .I0(n15969[5]), .I1(n533_adj_4762), 
            .CO(n38531));
    SB_LUT4 add_5052_7_lut (.I0(GND_net), .I1(n15969[4]), .I2(n460_adj_4763), 
            .I3(n38529), .O(n15425[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n37665), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n37666));
    SB_CARRY add_5052_7 (.CI(n38529), .I0(n15969[4]), .I1(n460_adj_4763), 
            .CO(n38530));
    SB_LUT4 add_5052_6_lut (.I0(GND_net), .I1(n15969[3]), .I2(n387_adj_4764), 
            .I3(n38528), .O(n15425[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4765));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4766));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n37664), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n37584), .O(duty_23__N_3772[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_6 (.CI(n38528), .I0(n15969[3]), .I1(n387_adj_4764), 
            .CO(n38529));
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4767));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4768));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4769));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5052_5_lut (.I0(GND_net), .I1(n15969[2]), .I2(n314_adj_4770), 
            .I3(n38527), .O(n15425[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20010_2_lut (.I0(n28[6]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20010_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5052_5 (.CI(n38527), .I0(n15969[2]), .I1(n314_adj_4770), 
            .CO(n38528));
    SB_CARRY add_12_21 (.CI(n37584), .I0(n106[19]), .I1(n155[19]), .CO(n37585));
    SB_LUT4 add_5052_4_lut (.I0(GND_net), .I1(n15969[1]), .I2(n241_adj_4771), 
            .I3(n38526), .O(n15425[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20009_2_lut (.I0(n28[7]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20009_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n37583), .O(duty_23__N_3772[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_9 (.CI(n37664), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n37665));
    SB_LUT4 i20008_2_lut (.I0(n28[8]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20008_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31949_4_lut (.I0(n21_adj_4772), .I1(n19_adj_4773), .I2(n17_adj_4774), 
            .I3(n9_adj_4775), .O(n47080));
    defparam i31949_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n37663), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_20 (.CI(n37583), .I0(n106[18]), .I1(n155[18]), .CO(n37584));
    SB_CARRY sub_3_add_2_8 (.CI(n37663), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n37664));
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n37582), .O(duty_23__N_3772[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n37662), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5052_4 (.CI(n38526), .I0(n15969[1]), .I1(n241_adj_4771), 
            .CO(n38527));
    SB_LUT4 add_5052_3_lut (.I0(GND_net), .I1(n15969[0]), .I2(n168_adj_4778), 
            .I3(n38525), .O(n15425[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n37582), .I0(n106[17]), .I1(n155[17]), .CO(n37583));
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4779));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_7 (.CI(n37662), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n37663));
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n37661), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5052_3 (.CI(n38525), .I0(n15969[0]), .I1(n168_adj_4778), 
            .CO(n38526));
    SB_LUT4 add_5052_2_lut (.I0(GND_net), .I1(n26_adj_4781), .I2(n95_adj_4782), 
            .I3(GND_net), .O(n15425[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5052_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5052_2 (.CI(GND_net), .I0(n26_adj_4781), .I1(n95_adj_4782), 
            .CO(n38525));
    SB_CARRY sub_3_add_2_6 (.CI(n37661), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n37662));
    SB_LUT4 i20007_2_lut (.I0(n28[9]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20007_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n37660), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_5 (.CI(n37660), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n37661));
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n37581), .O(duty_23__N_3772[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5252_9_lut (.I0(GND_net), .I1(n18416[6]), .I2(n630_adj_4783), 
            .I3(n38524), .O(n18289[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4784));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31882_2_lut (.I0(n43), .I1(n19_adj_4773), .I2(GND_net), .I3(GND_net), 
            .O(n47013));
    defparam i31882_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4774), .I3(GND_net), 
            .O(n8_adj_4785));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4786));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5252_8_lut (.I0(GND_net), .I1(n18416[5]), .I2(n557_adj_4787), 
            .I3(n38523), .O(n18289[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_18 (.CI(n37581), .I0(n106[16]), .I1(n155[16]), .CO(n37582));
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n37659), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_8 (.CI(n38523), .I0(n18416[5]), .I1(n557_adj_4787), 
            .CO(n38524));
    SB_LUT4 i20006_2_lut (.I0(n28[10]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20006_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5208_11_lut (.I0(GND_net), .I1(n18029[8]), .I2(n770), 
            .I3(n37758), .O(n17809[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_4 (.CI(n37659), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n37660));
    SB_LUT4 i20005_2_lut (.I0(n28[11]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20005_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5208_10_lut (.I0(GND_net), .I1(n18029[7]), .I2(n697), 
            .I3(n37757), .O(n17809[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5252_7_lut (.I0(GND_net), .I1(n18416[4]), .I2(n484_adj_4789), 
            .I3(n38522), .O(n18289[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n37658), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_7 (.CI(n38522), .I0(n18416[4]), .I1(n484_adj_4789), 
            .CO(n38523));
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5252_6_lut (.I0(GND_net), .I1(n18416[3]), .I2(n411_adj_4790), 
            .I3(n38521), .O(n18289[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n37658), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n37659));
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20004_2_lut (.I0(n28[12]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20004_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n37580), .O(duty_23__N_3772[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_10 (.CI(n37757), .I0(n18029[7]), .I1(n697), .CO(n37758));
    SB_CARRY add_5252_6 (.CI(n38521), .I0(n18416[3]), .I1(n411_adj_4790), 
            .CO(n38522));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4779), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4791));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i31966_2_lut (.I0(n7_adj_4792), .I1(n5_adj_4793), .I2(GND_net), 
            .I3(GND_net), .O(n47097));
    defparam i31966_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_5208_9_lut (.I0(GND_net), .I1(n18029[6]), .I2(n624), .I3(n37756), 
            .O(n17809[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32224_4_lut (.I0(n13_adj_4757), .I1(n11_adj_4758), .I2(n9_adj_4775), 
            .I3(n47097), .O(n47356));
    defparam i32224_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5208_9 (.CI(n37756), .I0(n18029[6]), .I1(n624), .CO(n37757));
    SB_LUT4 add_5208_8_lut (.I0(GND_net), .I1(n18029[5]), .I2(n551), .I3(n37755), 
            .O(n17809[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_8 (.CI(n37755), .I0(n18029[5]), .I1(n551), .CO(n37756));
    SB_LUT4 i32220_4_lut (.I0(n19_adj_4773), .I1(n17_adj_4774), .I2(n15_adj_4756), 
            .I3(n47356), .O(n47352));
    defparam i32220_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32588_4_lut (.I0(n25_adj_4794), .I1(n23_adj_4795), .I2(n21_adj_4772), 
            .I3(n47352), .O(n47720));
    defparam i32588_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32404_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n47720), 
            .O(n47536));
    defparam i32404_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32620_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n47536), 
            .O(n47752));
    defparam i32620_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5252_5_lut (.I0(GND_net), .I1(n18416[2]), .I2(n338_adj_4796), 
            .I3(n38520), .O(n18289[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5208_7_lut (.I0(GND_net), .I1(n18029[4]), .I2(n478), .I3(n37754), 
            .O(n17809[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20013_2_lut (.I0(n28[3]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20013_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5208_7 (.CI(n37754), .I0(n18029[4]), .I1(n478), .CO(n37755));
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5208_6_lut (.I0(GND_net), .I1(n18029[3]), .I2(n405), .I3(n37753), 
            .O(n17809[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20003_2_lut (.I0(n28[13]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20003_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32254_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n48927), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4740), .O(n47386));
    defparam i32254_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n37658));
    SB_CARRY add_5208_6 (.CI(n37753), .I0(n18029[3]), .I1(n405), .CO(n37754));
    SB_LUT4 add_5208_5_lut (.I0(GND_net), .I1(n18029[2]), .I2(n332), .I3(n37752), 
            .O(n17809[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_124_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n48896));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_124_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5208_5 (.CI(n37752), .I0(n18029[2]), .I1(n332), .CO(n37753));
    SB_LUT4 add_5208_4_lut (.I0(GND_net), .I1(n18029[1]), .I2(n259), .I3(n37751), 
            .O(n17809[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_4 (.CI(n37751), .I0(n18029[1]), .I1(n259), .CO(n37752));
    SB_LUT4 add_5208_3_lut (.I0(GND_net), .I1(n18029[0]), .I2(n186), .I3(n37750), 
            .O(n17809[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_5 (.CI(n38520), .I0(n18416[2]), .I1(n338_adj_4796), 
            .CO(n38521));
    SB_CARRY add_12_17 (.CI(n37580), .I0(n106[15]), .I1(n155[15]), .CO(n37581));
    SB_LUT4 i32242_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n48896), 
            .I2(IntegralLimit[14]), .I3(n47386), .O(n47374));
    defparam i32242_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_119_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n48891));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_119_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4797));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31978_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n47109));
    defparam i31978_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_142_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n48914));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_142_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4798));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4797), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32522_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n48909), 
            .I2(IntegralLimit[11]), .I3(n47384), .O(n47654));
    defparam i32522_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n37579), .O(duty_23__N_3772[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_3 (.CI(n37750), .I0(n18029[0]), .I1(n186), .CO(n37751));
    SB_LUT4 add_5252_4_lut (.I0(GND_net), .I1(n18416[1]), .I2(n265_adj_4728), 
            .I3(n38519), .O(n18289[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3772[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_16 (.CI(n37579), .I0(n106[14]), .I1(n155[14]), .CO(n37580));
    SB_LUT4 duty_23__I_851_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3772[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4800));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5208_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n17809[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n37578), .O(duty_23__N_3772[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3772[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4801));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4802));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3772[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4803));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_15 (.CI(n37578), .I0(n106[13]), .I1(n155[13]), .CO(n37579));
    SB_LUT4 duty_23__I_851_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3772[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4804));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5208_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n37750));
    SB_CARRY add_5252_4 (.CI(n38519), .I0(n18416[1]), .I1(n265_adj_4728), 
            .CO(n38520));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n37577), .O(duty_23__N_3772[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n37577), .I0(n106[12]), .I1(n155[12]), .CO(n37578));
    SB_LUT4 duty_23__I_851_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3772[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4805));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3772[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4806));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3772[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4807));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n37576), .O(duty_23__N_3772[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3772[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4809));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5252_3_lut (.I0(GND_net), .I1(n18416[0]), .I2(n192_adj_4721), 
            .I3(n38518), .O(n18289[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31986_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n48903), 
            .I2(IntegralLimit[13]), .I3(n47654), .O(n47117));
    defparam i31986_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 duty_23__I_851_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3772[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4811));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3772[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4812));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3772[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4813));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3772[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4814));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4815));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3772[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4816));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_851_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3772[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4817));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5252_3 (.CI(n38518), .I0(n18416[0]), .I1(n192_adj_4721), 
            .CO(n38519));
    SB_CARRY add_12_13 (.CI(n37576), .I0(n106[11]), .I1(n155[11]), .CO(n37577));
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n37575), .O(duty_23__N_3772[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3772[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4818));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_12 (.CI(n37575), .I0(n106[10]), .I1(n155[10]), .CO(n37576));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n37574), 
            .O(duty_23__N_3772[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n37574), .I0(n106[9]), .I1(n155[9]), .CO(n37575));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n37573), 
            .O(duty_23__N_3772[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5252_2_lut (.I0(GND_net), .I1(n50_adj_4720), .I2(n119_adj_4719), 
            .I3(GND_net), .O(n18289[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_2 (.CI(GND_net), .I0(n50_adj_4720), .I1(n119_adj_4719), 
            .CO(n38518));
    SB_CARRY add_12_10 (.CI(n37573), .I0(n106[8]), .I1(n155[8]), .CO(n37574));
    SB_LUT4 add_5083_16_lut (.I0(GND_net), .I1(n16449[13]), .I2(n1120), 
            .I3(n38517), .O(n15969[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3772[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4820));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31857_4_lut (.I0(n21_adj_4820), .I1(n19_adj_4818), .I2(n17_adj_4817), 
            .I3(n9_adj_4816), .O(n46988));
    defparam i31857_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31851_4_lut (.I0(n27_adj_4814), .I1(n15_adj_4813), .I2(n13_adj_4812), 
            .I3(n11_adj_4811), .O(n46982));
    defparam i31851_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_851_i12_3_lut (.I0(duty_23__N_3772[7]), .I1(duty_23__N_3772[16]), 
            .I2(n33_adj_4815), .I3(GND_net), .O(n12_adj_4821));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_122_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n48894));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_122_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5083_15_lut (.I0(GND_net), .I1(n16449[12]), .I2(n1047), 
            .I3(n38516), .O(n15969[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n37572), 
            .O(duty_23__N_3772[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_851_i10_3_lut (.I0(duty_23__N_3772[5]), .I1(duty_23__N_3772[6]), 
            .I2(n13_adj_4812), .I3(GND_net), .O(n10_adj_4823));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5083_15 (.CI(n38516), .I0(n16449[12]), .I1(n1047), .CO(n38517));
    SB_LUT4 duty_23__I_851_i30_3_lut (.I0(n12_adj_4821), .I1(duty_23__N_3772[17]), 
            .I2(n35_adj_4809), .I3(GND_net), .O(n30_adj_4824));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_12_9 (.CI(n37572), .I0(n106[7]), .I1(n155[7]), .CO(n37573));
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n37571), 
            .O(duty_23__N_3772[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32170_4_lut (.I0(n13_adj_4812), .I1(n11_adj_4811), .I2(n9_adj_4816), 
            .I3(n47011), .O(n47302));
    defparam i32170_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32430_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n48894), 
            .I2(IntegralLimit[15]), .I3(n47117), .O(n47562));
    defparam i32430_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_12_8 (.CI(n37571), .I0(n106[6]), .I1(n155[6]), .CO(n37572));
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_148_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n48920));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_148_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32592_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n48920), 
            .I2(IntegralLimit[17]), .I3(n47562), .O(n47724));
    defparam i32592_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_113_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n48885));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_113_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5083_14_lut (.I0(GND_net), .I1(n16449[11]), .I2(n974), 
            .I3(n38515), .O(n15969[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n37570), 
            .O(duty_23__N_3772[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_12_7 (.CI(n37570), .I0(n106[5]), .I1(n155[5]), .CO(n37571));
    SB_CARRY add_5083_14 (.CI(n38515), .I0(n16449[11]), .I1(n974), .CO(n38516));
    SB_LUT4 i32648_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n48885), 
            .I2(IntegralLimit[19]), .I3(n47724), .O(n47780));
    defparam i32648_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i32154_4_lut (.I0(n19_adj_4818), .I1(n17_adj_4817), .I2(n15_adj_4813), 
            .I3(n47302), .O(n47286));
    defparam i32154_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32558_4_lut (.I0(n25_adj_4807), .I1(n23_adj_4806), .I2(n21_adj_4820), 
            .I3(n47286), .O(n47690));
    defparam i32558_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_110_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n48882));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_110_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32358_4_lut (.I0(n31_adj_4804), .I1(n29_adj_4803), .I2(n27_adj_4814), 
            .I3(n47690), .O(n47490));
    defparam i32358_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4826));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n37569), 
            .O(duty_23__N_3772[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_13_lut (.I0(GND_net), .I1(n16449[10]), .I2(n901), 
            .I3(n38514), .O(n15969[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32614_4_lut (.I0(n37_adj_4805), .I1(n35_adj_4809), .I2(n33_adj_4815), 
            .I3(n47490), .O(n47746));
    defparam i32614_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_5083_13 (.CI(n38514), .I0(n16449[10]), .I1(n901), .CO(n38515));
    SB_LUT4 add_5083_12_lut (.I0(GND_net), .I1(n16449[9]), .I2(n828), 
            .I3(n38513), .O(n15969[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31968_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n47099));
    defparam i31968_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 duty_23__I_851_i16_3_lut (.I0(duty_23__N_3772[9]), .I1(duty_23__N_3772[21]), 
            .I2(n43_adj_4802), .I3(GND_net), .O(n16_adj_4828));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32564_3_lut (.I0(n6), .I1(duty_23__N_3772[10]), .I2(n21_adj_4820), 
            .I3(GND_net), .O(n47696));   // verilog/motorControl.v(36[10:25])
    defparam i32564_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i32565_3_lut (.I0(n47696), .I1(duty_23__N_3772[11]), .I2(n23_adj_4806), 
            .I3(GND_net), .O(n47697));   // verilog/motorControl.v(36[10:25])
    defparam i32565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5083_12 (.CI(n38513), .I0(n16449[9]), .I1(n828), .CO(n38514));
    SB_LUT4 add_5083_11_lut (.I0(GND_net), .I1(n16449[8]), .I2(n755), 
            .I3(n38512), .O(n15969[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_11 (.CI(n38512), .I0(n16449[8]), .I1(n755), .CO(n38513));
    SB_LUT4 duty_23__I_851_i8_3_lut (.I0(duty_23__N_3772[4]), .I1(duty_23__N_3772[8]), 
            .I2(n17_adj_4817), .I3(GND_net), .O(n8_adj_4830));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_851_i24_3_lut (.I0(n16_adj_4828), .I1(duty_23__N_3772[22]), 
            .I2(n45_adj_4801), .I3(GND_net), .O(n24_adj_4831));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4826), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4832));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4833));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32514_3_lut (.I0(n6_adj_4833), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n47646));   // verilog/motorControl.v(31[10:34])
    defparam i32514_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32515_3_lut (.I0(n47646), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n47647));   // verilog/motorControl.v(31[10:34])
    defparam i32515_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i31970_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n48903), 
            .I2(IntegralLimit[21]), .I3(n47380), .O(n47101));
    defparam i31970_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i31834_4_lut (.I0(n43_adj_4802), .I1(n25_adj_4807), .I2(n23_adj_4806), 
            .I3(n46988), .O(n46965));
    defparam i31834_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32392_4_lut (.I0(n24_adj_4831), .I1(n8_adj_4830), .I2(n45_adj_4801), 
            .I3(n46962), .O(n47524));   // verilog/motorControl.v(36[10:25])
    defparam i32392_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32485_3_lut (.I0(n47697), .I1(duty_23__N_3772[12]), .I2(n25_adj_4807), 
            .I3(GND_net), .O(n47617));   // verilog/motorControl.v(36[10:25])
    defparam i32485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20002_2_lut (.I0(n28[14]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20002_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4836));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_851_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(duty_23__N_3772[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4837));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_851_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4838));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32530_3_lut (.I0(n4_adj_4837), .I1(duty_23__N_3772[13]), .I2(n27_adj_4814), 
            .I3(GND_net), .O(n47662));   // verilog/motorControl.v(36[10:25])
    defparam i32530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4839));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_107_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n48879));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_107_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32531_3_lut (.I0(n47662), .I1(duty_23__N_3772[14]), .I2(n29_adj_4803), 
            .I3(GND_net), .O(n47663));   // verilog/motorControl.v(36[10:25])
    defparam i32531_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31846_4_lut (.I0(n33_adj_4815), .I1(n31_adj_4804), .I2(n29_adj_4803), 
            .I3(n46982), .O(n46977));
    defparam i31846_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32630_4_lut (.I0(n30_adj_4824), .I1(n10_adj_4823), .I2(n35_adj_4809), 
            .I3(n46975), .O(n47762));   // verilog/motorControl.v(36[10:25])
    defparam i32630_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32487_3_lut (.I0(n47663), .I1(duty_23__N_3772[15]), .I2(n31_adj_4804), 
            .I3(GND_net), .O(n47619));   // verilog/motorControl.v(36[10:25])
    defparam i32487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32670_4_lut (.I0(n47619), .I1(n47762), .I2(n35_adj_4809), 
            .I3(n46977), .O(n47802));   // verilog/motorControl.v(36[10:25])
    defparam i32670_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32671_3_lut (.I0(n47802), .I1(duty_23__N_3772[18]), .I2(n37_adj_4805), 
            .I3(GND_net), .O(n47803));   // verilog/motorControl.v(36[10:25])
    defparam i32671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32659_3_lut (.I0(n47803), .I1(duty_23__N_3772[19]), .I2(n39), 
            .I3(GND_net), .O(n47791));   // verilog/motorControl.v(36[10:25])
    defparam i32659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32388_4_lut (.I0(n24_adj_4832), .I1(n8_adj_4841), .I2(n48879), 
            .I3(n47099), .O(n47520));   // verilog/motorControl.v(31[10:34])
    defparam i32388_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4842));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31836_4_lut (.I0(n43_adj_4802), .I1(n41_adj_4800), .I2(n39), 
            .I3(n47746), .O(n46967));
    defparam i31836_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32179_3_lut (.I0(n47647), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n47311));   // verilog/motorControl.v(31[10:34])
    defparam i32179_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32574_4_lut (.I0(n47617), .I1(n47524), .I2(n45_adj_4801), 
            .I3(n46965), .O(n47706));   // verilog/motorControl.v(36[10:25])
    defparam i32574_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32641_3_lut (.I0(n47791), .I1(duty_23__N_3772[20]), .I2(n41_adj_4800), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(36[10:25])
    defparam i32641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32576_4_lut (.I0(n40), .I1(n47706), .I2(n45_adj_4801), .I3(n46967), 
            .O(n47708));   // verilog/motorControl.v(36[10:25])
    defparam i32576_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32577_3_lut (.I0(n47708), .I1(PWMLimit[23]), .I2(duty_23__N_3772[23]), 
            .I3(GND_net), .O(duty_23__N_3771));   // verilog/motorControl.v(36[10:25])
    defparam i32577_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4843));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3772[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4844));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5083_10_lut (.I0(GND_net), .I1(n16449[7]), .I2(n682), 
            .I3(n38511), .O(n15969[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_10 (.CI(n38511), .I0(n16449[7]), .I1(n682), .CO(n38512));
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3772[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4845));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4846));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5083_9_lut (.I0(GND_net), .I1(n16449[6]), .I2(n609), .I3(n38510), 
            .O(n15969[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_9 (.CI(n38510), .I0(n16449[6]), .I1(n609), .CO(n38511));
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3772[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4847));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5083_8_lut (.I0(GND_net), .I1(n16449[5]), .I2(n536), .I3(n38509), 
            .O(n15969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_8 (.CI(n38509), .I0(n16449[5]), .I1(n536), .CO(n38510));
    SB_LUT4 add_5083_7_lut (.I0(GND_net), .I1(n16449[4]), .I2(n463), .I3(n38508), 
            .O(n15969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_7 (.CI(n38508), .I0(n16449[4]), .I1(n463), .CO(n38509));
    SB_LUT4 add_5083_6_lut (.I0(GND_net), .I1(n16449[3]), .I2(n390), .I3(n38507), 
            .O(n15969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_6 (.CI(n37569), .I0(n106[4]), .I1(n155[4]), .CO(n37570));
    SB_CARRY add_5083_6 (.CI(n38507), .I0(n16449[3]), .I1(n390), .CO(n38508));
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n37568), 
            .O(duty_23__N_3772[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5083_5_lut (.I0(GND_net), .I1(n16449[2]), .I2(n317), .I3(n38506), 
            .O(n15969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_5 (.CI(n38506), .I0(n16449[2]), .I1(n317), .CO(n38507));
    SB_LUT4 add_5083_4_lut (.I0(GND_net), .I1(n16449[1]), .I2(n244), .I3(n38505), 
            .O(n15969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_4 (.CI(n38505), .I0(n16449[1]), .I1(n244), .CO(n38506));
    SB_LUT4 add_5083_3_lut (.I0(GND_net), .I1(n16449[0]), .I2(n171), .I3(n38504), 
            .O(n15969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5083_3 (.CI(n38504), .I0(n16449[0]), .I1(n171), .CO(n38505));
    SB_LUT4 add_5083_2_lut (.I0(GND_net), .I1(n29_adj_4848), .I2(n98), 
            .I3(GND_net), .O(n15969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5083_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_5 (.CI(n37568), .I0(n106[3]), .I1(n155[3]), .CO(n37569));
    SB_CARRY add_5083_2 (.CI(GND_net), .I0(n29_adj_4848), .I1(n98), .CO(n38504));
    SB_LUT4 add_5112_15_lut (.I0(GND_net), .I1(n16869[12]), .I2(n1050), 
            .I3(n38503), .O(n16449[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5112_14_lut (.I0(GND_net), .I1(n16869[11]), .I2(n977), 
            .I3(n38502), .O(n16449[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4849));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5112_14 (.CI(n38502), .I0(n16869[11]), .I1(n977), .CO(n38503));
    SB_LUT4 add_5112_13_lut (.I0(GND_net), .I1(n16869[10]), .I2(n904), 
            .I3(n38501), .O(n16449[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5112_13 (.CI(n38501), .I0(n16869[10]), .I1(n904), .CO(n38502));
    SB_LUT4 add_5112_12_lut (.I0(GND_net), .I1(n16869[9]), .I2(n831), 
            .I3(n38500), .O(n16449[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3723 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4850), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4851));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_CARRY add_5112_12 (.CI(n38500), .I0(n16869[9]), .I1(n831), .CO(n38501));
    SB_LUT4 add_5112_11_lut (.I0(GND_net), .I1(n16869[8]), .I2(n758), 
            .I3(n38499), .O(n16449[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32422_3_lut (.I0(n4_adj_4851), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n47554));   // verilog/motorControl.v(31[38:63])
    defparam i32422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4852));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4853));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4796));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4854));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4855));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3772[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4856));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3772[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4857));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3772[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4858));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5112_11 (.CI(n38499), .I0(n16869[8]), .I1(n758), .CO(n38500));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n28[23]), .I1(n11121[21]), .I2(GND_net), 
            .I3(n38923), .O(n10614[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n11121[20]), .I2(GND_net), 
            .I3(n38922), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4860));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_23 (.CI(n38922), .I0(n11121[20]), .I1(GND_net), 
            .CO(n38923));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n11121[19]), .I2(GND_net), 
            .I3(n38921), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n38921), .I0(n11121[19]), .I1(GND_net), 
            .CO(n38922));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n11121[18]), .I2(GND_net), 
            .I3(n38920), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n38920), .I0(n11121[18]), .I1(GND_net), 
            .CO(n38921));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n11121[17]), .I2(GND_net), 
            .I3(n38919), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n38919), .I0(n11121[17]), .I1(GND_net), 
            .CO(n38920));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n11121[16]), .I2(GND_net), 
            .I3(n38918), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n38918), .I0(n11121[16]), .I1(GND_net), 
            .CO(n38919));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n11121[15]), .I2(GND_net), 
            .I3(n38917), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n38917), .I0(n11121[15]), .I1(GND_net), 
            .CO(n38918));
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n37567), 
            .O(duty_23__N_3772[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4861));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5112_10_lut (.I0(GND_net), .I1(n16869[7]), .I2(n685), 
            .I3(n38498), .O(n16449[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n11121[14]), .I2(GND_net), 
            .I3(n38916), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n37726), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n38916), .I0(n11121[14]), .I1(GND_net), 
            .CO(n38917));
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4862));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4863));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32423_3_lut (.I0(n47554), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n47555));   // verilog/motorControl.v(31[38:63])
    defparam i32423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3772[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4864));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3772[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4865));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3772[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4866));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4867));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n11121[13]), .I2(n1096), 
            .I3(n38915), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n38915), .I0(n11121[13]), .I1(n1096), 
            .CO(n38916));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n11121[12]), .I2(n1023), 
            .I3(n38914), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4868));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3772[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4869));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_15 (.CI(n38914), .I0(n11121[12]), .I1(n1023), 
            .CO(n38915));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n11121[11]), .I2(n950), 
            .I3(n38913), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n38913), .I0(n11121[11]), .I1(n950), 
            .CO(n38914));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n11121[10]), .I2(n877), 
            .I3(n38912), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n38912), .I0(n11121[10]), .I1(n877), 
            .CO(n38913));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n11121[9]), .I2(n804), 
            .I3(n38911), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n38911), .I0(n11121[9]), .I1(n804), 
            .CO(n38912));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n11121[8]), .I2(n731), 
            .I3(n38910), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n38910), .I0(n11121[8]), .I1(n731), 
            .CO(n38911));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n11121[7]), .I2(n658), 
            .I3(n38909), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n38909), .I0(n11121[7]), .I1(n658), 
            .CO(n38910));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n11121[6]), .I2(n585), 
            .I3(n38908), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n38908), .I0(n11121[6]), .I1(n585), 
            .CO(n38909));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n11121[5]), .I2(n512), 
            .I3(n38907), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3772[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4870));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_12_4 (.CI(n37567), .I0(n106[2]), .I1(n155[2]), .CO(n37568));
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3772[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4871));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY mult_10_add_1225_8 (.CI(n38907), .I0(n11121[5]), .I1(n512), 
            .CO(n38908));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n11121[4]), .I2(n439), 
            .I3(n38906), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n38906), .I0(n11121[4]), .I1(n439), 
            .CO(n38907));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n11121[3]), .I2(n366), 
            .I3(n38905), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n38905), .I0(n11121[3]), .I1(n366), 
            .CO(n38906));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n11121[2]), .I2(n293), 
            .I3(n38904), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n38904), .I0(n11121[2]), .I1(n293), 
            .CO(n38905));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n11121[1]), .I2(n220), 
            .I3(n38903), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n38903), .I0(n11121[1]), .I1(n220), 
            .CO(n38904));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n11121[0]), .I2(n147), 
            .I3(n38902), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n38902), .I0(n11121[0]), .I1(n147), 
            .CO(n38903));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4786), .I2(n74), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4786), .I1(n74), 
            .CO(n38902));
    SB_LUT4 add_4846_23_lut (.I0(GND_net), .I1(n12088[20]), .I2(GND_net), 
            .I3(n38901), .O(n11121[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4846_22_lut (.I0(GND_net), .I1(n12088[19]), .I2(GND_net), 
            .I3(n38900), .O(n11121[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3772[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4873));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3772[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4874));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3772[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4875));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3772[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4876));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3772[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4877));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i31816_4_lut (.I0(n21_adj_4877), .I1(n19_adj_4876), .I2(n17_adj_4875), 
            .I3(n9_adj_4874), .O(n46947));
    defparam i31816_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i31934_2_lut (.I0(n33), .I1(n15_adj_4756), .I2(GND_net), .I3(GND_net), 
            .O(n47065));
    defparam i31934_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4757), .I3(GND_net), 
            .O(n10_adj_4878));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i31810_4_lut (.I0(n27_adj_4873), .I1(n15_adj_4871), .I2(n13_adj_4870), 
            .I3(n11_adj_4869), .O(n46941));
    defparam i31810_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4868), 
            .I3(GND_net), .O(n12_adj_4879));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4867), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_4880));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i31936_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n47071), 
            .O(n47067));
    defparam i31936_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4870), 
            .I3(GND_net), .O(n10_adj_4881));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4879), .I1(n257[17]), .I2(n35_adj_4866), 
            .I3(GND_net), .O(n30_adj_4882));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4846_22 (.CI(n38900), .I0(n12088[19]), .I1(GND_net), 
            .CO(n38901));
    SB_LUT4 i32110_4_lut (.I0(n13_adj_4870), .I1(n11_adj_4869), .I2(n9_adj_4874), 
            .I3(n46960), .O(n47242));
    defparam i32110_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32106_4_lut (.I0(n19_adj_4876), .I1(n17_adj_4875), .I2(n15_adj_4871), 
            .I3(n47242), .O(n47238));
    defparam i32106_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32550_4_lut (.I0(n25_adj_4865), .I1(n23_adj_4864), .I2(n21_adj_4877), 
            .I3(n47238), .O(n47682));
    defparam i32550_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32338_4_lut (.I0(n31_adj_4858), .I1(n29_adj_4857), .I2(n27_adj_4873), 
            .I3(n47682), .O(n47470));
    defparam i32338_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4846_21_lut (.I0(GND_net), .I1(n12088[18]), .I2(GND_net), 
            .I3(n38899), .O(n11121[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_21 (.CI(n38899), .I0(n12088[18]), .I1(GND_net), 
            .CO(n38900));
    SB_LUT4 add_4846_20_lut (.I0(GND_net), .I1(n12088[17]), .I2(GND_net), 
            .I3(n38898), .O(n11121[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_20 (.CI(n38898), .I0(n12088[17]), .I1(GND_net), 
            .CO(n38899));
    SB_LUT4 add_4846_19_lut (.I0(GND_net), .I1(n12088[16]), .I2(GND_net), 
            .I3(n38897), .O(n11121[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_19 (.CI(n38897), .I0(n12088[16]), .I1(GND_net), 
            .CO(n38898));
    SB_LUT4 add_4846_18_lut (.I0(GND_net), .I1(n12088[15]), .I2(GND_net), 
            .I3(n38896), .O(n11121[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_18 (.CI(n38896), .I0(n12088[15]), .I1(GND_net), 
            .CO(n38897));
    SB_LUT4 add_4846_17_lut (.I0(GND_net), .I1(n12088[14]), .I2(GND_net), 
            .I3(n38895), .O(n11121[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n37566), 
            .O(duty_23__N_3772[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_17 (.CI(n38895), .I0(n12088[14]), .I1(GND_net), 
            .CO(n38896));
    SB_LUT4 add_4846_16_lut (.I0(GND_net), .I1(n12088[13]), .I2(n1099), 
            .I3(n38894), .O(n11121[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_16 (.CI(n38894), .I0(n12088[13]), .I1(n1099), .CO(n38895));
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n37725), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4846_15_lut (.I0(GND_net), .I1(n12088[12]), .I2(n1026), 
            .I3(n38893), .O(n11121[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_15 (.CI(n38893), .I0(n12088[12]), .I1(n1026), .CO(n38894));
    SB_CARRY add_5112_10 (.CI(n38498), .I0(n16869[7]), .I1(n685), .CO(n38499));
    SB_LUT4 add_4846_14_lut (.I0(GND_net), .I1(n12088[11]), .I2(n953), 
            .I3(n38892), .O(n11121[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_14 (.CI(n38892), .I0(n12088[11]), .I1(n953), .CO(n38893));
    SB_LUT4 add_4846_13_lut (.I0(GND_net), .I1(n12088[10]), .I2(n880), 
            .I3(n38891), .O(n11121[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_13 (.CI(n38891), .I0(n12088[10]), .I1(n880), .CO(n38892));
    SB_LUT4 add_4846_12_lut (.I0(GND_net), .I1(n12088[9]), .I2(n807), 
            .I3(n38890), .O(n11121[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_12 (.CI(n38890), .I0(n12088[9]), .I1(n807), .CO(n38891));
    SB_LUT4 add_4846_11_lut (.I0(GND_net), .I1(n12088[8]), .I2(n734), 
            .I3(n38889), .O(n11121[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_11 (.CI(n38889), .I0(n12088[8]), .I1(n734), .CO(n38890));
    SB_LUT4 add_4846_10_lut (.I0(GND_net), .I1(n12088[7]), .I2(n661), 
            .I3(n38888), .O(n11121[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_10 (.CI(n38888), .I0(n12088[7]), .I1(n661), .CO(n38889));
    SB_LUT4 add_4846_9_lut (.I0(GND_net), .I1(n12088[6]), .I2(n588), .I3(n38887), 
            .O(n11121[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_9 (.CI(n38887), .I0(n12088[6]), .I1(n588), .CO(n38888));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n37725), .I0(GND_net), .I1(n1[22]), 
            .CO(n37726));
    SB_LUT4 add_4846_8_lut (.I0(GND_net), .I1(n12088[5]), .I2(n515), .I3(n38886), 
            .O(n11121[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_8 (.CI(n38886), .I0(n12088[5]), .I1(n515), .CO(n38887));
    SB_LUT4 i32612_4_lut (.I0(n37_adj_4856), .I1(n35_adj_4866), .I2(n33_adj_4868), 
            .I3(n47470), .O(n47744));
    defparam i32612_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4854), 
            .I3(GND_net), .O(n16_adj_4884));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32546_3_lut (.I0(n6_adj_4885), .I1(n257[10]), .I2(n21_adj_4877), 
            .I3(GND_net), .O(n47678));   // verilog/motorControl.v(38[19:35])
    defparam i32546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4846_7_lut (.I0(GND_net), .I1(n12088[4]), .I2(n442), .I3(n38885), 
            .O(n11121[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_7 (.CI(n38885), .I0(n12088[4]), .I1(n442), .CO(n38886));
    SB_LUT4 add_4846_6_lut (.I0(GND_net), .I1(n12088[3]), .I2(n369), .I3(n38884), 
            .O(n11121[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_6 (.CI(n38884), .I0(n12088[3]), .I1(n369), .CO(n38885));
    SB_LUT4 add_4846_5_lut (.I0(GND_net), .I1(n12088[2]), .I2(n296), .I3(n38883), 
            .O(n11121[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_5 (.CI(n38883), .I0(n12088[2]), .I1(n296), .CO(n38884));
    SB_LUT4 add_4846_4_lut (.I0(GND_net), .I1(n12088[1]), .I2(n223), .I3(n38882), 
            .O(n11121[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_4 (.CI(n38882), .I0(n12088[1]), .I1(n223), .CO(n38883));
    SB_LUT4 add_4846_3_lut (.I0(GND_net), .I1(n12088[0]), .I2(n150), .I3(n38881), 
            .O(n11121[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_3 (.CI(n38881), .I0(n12088[0]), .I1(n150), .CO(n38882));
    SB_LUT4 add_4846_2_lut (.I0(GND_net), .I1(n8_adj_4734), .I2(n77), 
            .I3(GND_net), .O(n11121[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4846_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4846_2 (.CI(GND_net), .I0(n8_adj_4734), .I1(n77), .CO(n38881));
    SB_LUT4 add_4888_22_lut (.I0(GND_net), .I1(n12969[19]), .I2(GND_net), 
            .I3(n38880), .O(n12088[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4888_21_lut (.I0(GND_net), .I1(n12969[18]), .I2(GND_net), 
            .I3(n38879), .O(n12088[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_21 (.CI(n38879), .I0(n12969[18]), .I1(GND_net), 
            .CO(n38880));
    SB_LUT4 add_4888_20_lut (.I0(GND_net), .I1(n12969[17]), .I2(GND_net), 
            .I3(n38878), .O(n12088[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_20 (.CI(n38878), .I0(n12969[17]), .I1(GND_net), 
            .CO(n38879));
    SB_LUT4 add_4888_19_lut (.I0(GND_net), .I1(n12969[16]), .I2(GND_net), 
            .I3(n38877), .O(n12088[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_19 (.CI(n38877), .I0(n12969[16]), .I1(GND_net), 
            .CO(n38878));
    SB_LUT4 add_4888_18_lut (.I0(GND_net), .I1(n12969[15]), .I2(GND_net), 
            .I3(n38876), .O(n12088[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n37724), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32538_4_lut (.I0(n30_adj_4880), .I1(n10_adj_4878), .I2(n35), 
            .I3(n47065), .O(n47670));   // verilog/motorControl.v(31[38:63])
    defparam i32538_4_lut.LUT_INIT = 16'haaac;
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3672 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3648[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3648[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3648[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3648[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3648[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3648[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3648[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3648[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3648[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3648[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3648[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3648[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3648[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3648[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3648[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3648[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3648[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i32547_3_lut (.I0(n47678), .I1(n257[11]), .I2(n23_adj_4864), 
            .I3(GND_net), .O(n47679));   // verilog/motorControl.v(38[19:35])
    defparam i32547_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3648[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3648[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3648[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3648[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3648[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3648[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4886));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n37724), .I0(GND_net), .I1(n1[21]), 
            .CO(n37725));
    SB_CARRY add_4888_18 (.CI(n38876), .I0(n12969[15]), .I1(GND_net), 
            .CO(n38877));
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4887));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4875), 
            .I3(GND_net), .O(n8_adj_4888));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4884), .I1(n257[22]), .I2(n45_adj_4847), 
            .I3(GND_net), .O(n24_adj_4889));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31791_4_lut (.I0(n43_adj_4854), .I1(n25_adj_4865), .I2(n23_adj_4864), 
            .I3(n46947), .O(n46922));
    defparam i31791_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32394_4_lut (.I0(n24_adj_4889), .I1(n8_adj_4888), .I2(n45_adj_4847), 
            .I3(n46920), .O(n47526));   // verilog/motorControl.v(38[19:35])
    defparam i32394_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32491_3_lut (.I0(n47679), .I1(n257[12]), .I2(n25_adj_4865), 
            .I3(GND_net), .O(n47623));   // verilog/motorControl.v(38[19:35])
    defparam i32491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4890));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4891));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3772[0]), .I1(n257[1]), 
            .I2(duty_23__N_3772[1]), .I3(n257[0]), .O(n4_adj_4892));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_5112_9_lut (.I0(GND_net), .I1(n16869[6]), .I2(n612), .I3(n38497), 
            .O(n16449[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4893));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4888_17_lut (.I0(GND_net), .I1(n12969[14]), .I2(GND_net), 
            .I3(n38875), .O(n12088[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_17 (.CI(n38875), .I0(n12969[14]), .I1(GND_net), 
            .CO(n38876));
    SB_LUT4 add_4888_16_lut (.I0(GND_net), .I1(n12969[13]), .I2(n1102), 
            .I3(n38874), .O(n12088[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_16 (.CI(n38874), .I0(n12969[13]), .I1(n1102), .CO(n38875));
    SB_LUT4 add_4888_15_lut (.I0(GND_net), .I1(n12969[12]), .I2(n1029), 
            .I3(n38873), .O(n12088[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_15 (.CI(n38873), .I0(n12969[12]), .I1(n1029), .CO(n38874));
    SB_LUT4 i32191_3_lut (.I0(n47555), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n47323));   // verilog/motorControl.v(31[38:63])
    defparam i32191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4888_14_lut (.I0(GND_net), .I1(n12969[11]), .I2(n956), 
            .I3(n38872), .O(n12088[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_14 (.CI(n38872), .I0(n12969[11]), .I1(n956), .CO(n38873));
    SB_LUT4 add_4888_13_lut (.I0(GND_net), .I1(n12969[10]), .I2(n883), 
            .I3(n38871), .O(n12088[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32646_4_lut (.I0(n47323), .I1(n47670), .I2(n35), .I3(n47067), 
            .O(n47778));   // verilog/motorControl.v(31[38:63])
    defparam i32646_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4888_13 (.CI(n38871), .I0(n12969[10]), .I1(n883), .CO(n38872));
    SB_LUT4 add_4888_12_lut (.I0(GND_net), .I1(n12969[9]), .I2(n810), 
            .I3(n38870), .O(n12088[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_12 (.CI(n38870), .I0(n12969[9]), .I1(n810), .CO(n38871));
    SB_LUT4 add_4888_11_lut (.I0(GND_net), .I1(n12969[8]), .I2(n737), 
            .I3(n38869), .O(n12088[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_11 (.CI(n38869), .I0(n12969[8]), .I1(n737), .CO(n38870));
    SB_LUT4 add_4888_10_lut (.I0(GND_net), .I1(n12969[7]), .I2(n664), 
            .I3(n38868), .O(n12088[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_10 (.CI(n38868), .I0(n12969[7]), .I1(n664), .CO(n38869));
    SB_LUT4 add_4888_9_lut (.I0(GND_net), .I1(n12969[6]), .I2(n591), .I3(n38867), 
            .O(n12088[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_9 (.CI(n38867), .I0(n12969[6]), .I1(n591), .CO(n38868));
    SB_LUT4 add_4888_8_lut (.I0(GND_net), .I1(n12969[5]), .I2(n518), .I3(n38866), 
            .O(n12088[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_8 (.CI(n38866), .I0(n12969[5]), .I1(n518), .CO(n38867));
    SB_LUT4 add_4888_7_lut (.I0(GND_net), .I1(n12969[4]), .I2(n445), .I3(n38865), 
            .O(n12088[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_7 (.CI(n38865), .I0(n12969[4]), .I1(n445), .CO(n38866));
    SB_LUT4 add_4888_6_lut (.I0(GND_net), .I1(n12969[3]), .I2(n372), .I3(n38864), 
            .O(n12088[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_6 (.CI(n38864), .I0(n12969[3]), .I1(n372), .CO(n38865));
    SB_LUT4 add_4888_5_lut (.I0(GND_net), .I1(n12969[2]), .I2(n299), .I3(n38863), 
            .O(n12088[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_5 (.CI(n38863), .I0(n12969[2]), .I1(n299), .CO(n38864));
    SB_LUT4 add_4888_4_lut (.I0(GND_net), .I1(n12969[1]), .I2(n226), .I3(n38862), 
            .O(n12088[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4894));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4888_4 (.CI(n38862), .I0(n12969[1]), .I1(n226), .CO(n38863));
    SB_LUT4 i32544_3_lut (.I0(n4_adj_4892), .I1(n257[13]), .I2(n27_adj_4873), 
            .I3(GND_net), .O(n47676));   // verilog/motorControl.v(38[19:35])
    defparam i32544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32545_3_lut (.I0(n47676), .I1(n257[14]), .I2(n29_adj_4857), 
            .I3(GND_net), .O(n47677));   // verilog/motorControl.v(38[19:35])
    defparam i32545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4888_3_lut (.I0(GND_net), .I1(n12969[0]), .I2(n153), .I3(n38861), 
            .O(n12088[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_3 (.CI(n38861), .I0(n12969[0]), .I1(n153), .CO(n38862));
    SB_LUT4 i31806_4_lut (.I0(n33_adj_4868), .I1(n31_adj_4858), .I2(n29_adj_4857), 
            .I3(n46941), .O(n46937));
    defparam i31806_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_4888_2_lut (.I0(GND_net), .I1(n11_adj_4725), .I2(n80), 
            .I3(GND_net), .O(n12088[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4888_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4888_2 (.CI(GND_net), .I0(n11_adj_4725), .I1(n80), .CO(n38861));
    SB_LUT4 add_4928_21_lut (.I0(GND_net), .I1(n13768[18]), .I2(GND_net), 
            .I3(n38860), .O(n12969[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4928_20_lut (.I0(GND_net), .I1(n13768[17]), .I2(GND_net), 
            .I3(n38859), .O(n12969[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_20 (.CI(n38859), .I0(n13768[17]), .I1(GND_net), 
            .CO(n38860));
    SB_LUT4 add_4928_19_lut (.I0(GND_net), .I1(n13768[16]), .I2(GND_net), 
            .I3(n38858), .O(n12969[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_19 (.CI(n38858), .I0(n13768[16]), .I1(GND_net), 
            .CO(n38859));
    SB_LUT4 add_4928_18_lut (.I0(GND_net), .I1(n13768[15]), .I2(GND_net), 
            .I3(n38857), .O(n12969[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_18 (.CI(n38857), .I0(n13768[15]), .I1(GND_net), 
            .CO(n38858));
    SB_LUT4 add_4928_17_lut (.I0(GND_net), .I1(n13768[14]), .I2(GND_net), 
            .I3(n38856), .O(n12969[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_17 (.CI(n38856), .I0(n13768[14]), .I1(GND_net), 
            .CO(n38857));
    SB_LUT4 i32632_4_lut (.I0(n30_adj_4882), .I1(n10_adj_4881), .I2(n35_adj_4866), 
            .I3(n46935), .O(n47764));   // verilog/motorControl.v(38[19:35])
    defparam i32632_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_4928_16_lut (.I0(GND_net), .I1(n13768[13]), .I2(n1105), 
            .I3(n38855), .O(n12969[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_16 (.CI(n38855), .I0(n13768[13]), .I1(n1105), .CO(n38856));
    SB_LUT4 add_4928_15_lut (.I0(GND_net), .I1(n13768[12]), .I2(n1032), 
            .I3(n38854), .O(n12969[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_15 (.CI(n38854), .I0(n13768[12]), .I1(n1032), .CO(n38855));
    SB_LUT4 add_4928_14_lut (.I0(GND_net), .I1(n13768[11]), .I2(n959), 
            .I3(n38853), .O(n12969[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_14 (.CI(n38853), .I0(n13768[11]), .I1(n959), .CO(n38854));
    SB_LUT4 add_4928_13_lut (.I0(GND_net), .I1(n13768[10]), .I2(n886), 
            .I3(n38852), .O(n12969[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_13 (.CI(n38852), .I0(n13768[10]), .I1(n886), .CO(n38853));
    SB_LUT4 add_4928_12_lut (.I0(GND_net), .I1(n13768[9]), .I2(n813), 
            .I3(n38851), .O(n12969[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_12 (.CI(n38851), .I0(n13768[9]), .I1(n813), .CO(n38852));
    SB_LUT4 add_4928_11_lut (.I0(GND_net), .I1(n13768[8]), .I2(n740), 
            .I3(n38850), .O(n12969[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_11 (.CI(n38850), .I0(n13768[8]), .I1(n740), .CO(n38851));
    SB_LUT4 add_4928_10_lut (.I0(GND_net), .I1(n13768[7]), .I2(n667), 
            .I3(n38849), .O(n12969[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n37723), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32647_3_lut (.I0(n47778), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n47779));   // verilog/motorControl.v(31[38:63])
    defparam i32647_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4896));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4897));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4928_10 (.CI(n38849), .I0(n13768[7]), .I1(n667), .CO(n38850));
    SB_LUT4 add_4928_9_lut (.I0(GND_net), .I1(n13768[6]), .I2(n594), .I3(n38848), 
            .O(n12969[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_9 (.CI(n38848), .I0(n13768[6]), .I1(n594), .CO(n38849));
    SB_LUT4 add_4928_8_lut (.I0(GND_net), .I1(n13768[5]), .I2(n521), .I3(n38847), 
            .O(n12969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_8 (.CI(n38847), .I0(n13768[5]), .I1(n521), .CO(n38848));
    SB_LUT4 add_4928_7_lut (.I0(GND_net), .I1(n13768[4]), .I2(n448), .I3(n38846), 
            .O(n12969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_7 (.CI(n38846), .I0(n13768[4]), .I1(n448), .CO(n38847));
    SB_LUT4 add_4928_6_lut (.I0(GND_net), .I1(n13768[3]), .I2(n375), .I3(n38845), 
            .O(n12969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_6 (.CI(n38845), .I0(n13768[3]), .I1(n375), .CO(n38846));
    SB_LUT4 add_4928_5_lut (.I0(GND_net), .I1(n13768[2]), .I2(n302), .I3(n38844), 
            .O(n12969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_5 (.CI(n38844), .I0(n13768[2]), .I1(n302), .CO(n38845));
    SB_LUT4 add_4928_4_lut (.I0(GND_net), .I1(n13768[1]), .I2(n229), .I3(n38843), 
            .O(n12969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_4 (.CI(n38843), .I0(n13768[1]), .I1(n229), .CO(n38844));
    SB_LUT4 add_4928_3_lut (.I0(GND_net), .I1(n13768[0]), .I2(n156), .I3(n38842), 
            .O(n12969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5112_9 (.CI(n38497), .I0(n16869[6]), .I1(n612), .CO(n38498));
    SB_CARRY add_4928_3 (.CI(n38842), .I0(n13768[0]), .I1(n156), .CO(n38843));
    SB_LUT4 add_4928_2_lut (.I0(GND_net), .I1(n14), .I2(n83), .I3(GND_net), 
            .O(n12969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4928_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4928_2 (.CI(GND_net), .I0(n14), .I1(n83), .CO(n38842));
    SB_LUT4 add_4966_20_lut (.I0(GND_net), .I1(n14489[17]), .I2(GND_net), 
            .I3(n38841), .O(n13768[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4966_19_lut (.I0(GND_net), .I1(n14489[16]), .I2(GND_net), 
            .I3(n38840), .O(n13768[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_19 (.CI(n38840), .I0(n14489[16]), .I1(GND_net), 
            .CO(n38841));
    SB_LUT4 add_4966_18_lut (.I0(GND_net), .I1(n14489[15]), .I2(GND_net), 
            .I3(n38839), .O(n13768[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_18 (.CI(n38839), .I0(n14489[15]), .I1(GND_net), 
            .CO(n38840));
    SB_LUT4 add_5112_8_lut (.I0(GND_net), .I1(n16869[5]), .I2(n539), .I3(n38496), 
            .O(n16449[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4966_17_lut (.I0(GND_net), .I1(n14489[14]), .I2(GND_net), 
            .I3(n38838), .O(n13768[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_17 (.CI(n38838), .I0(n14489[14]), .I1(GND_net), 
            .CO(n38839));
    SB_LUT4 add_4966_16_lut (.I0(GND_net), .I1(n14489[13]), .I2(n1108), 
            .I3(n38837), .O(n13768[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_16 (.CI(n38837), .I0(n14489[13]), .I1(n1108), .CO(n38838));
    SB_LUT4 i32493_3_lut (.I0(n47677), .I1(n257[15]), .I2(n31_adj_4858), 
            .I3(GND_net), .O(n47625));   // verilog/motorControl.v(38[19:35])
    defparam i32493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4966_15_lut (.I0(GND_net), .I1(n14489[12]), .I2(n1035), 
            .I3(n38836), .O(n13768[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32672_4_lut (.I0(n47625), .I1(n47764), .I2(n35_adj_4866), 
            .I3(n46937), .O(n47804));   // verilog/motorControl.v(38[19:35])
    defparam i32672_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4966_15 (.CI(n38836), .I0(n14489[12]), .I1(n1035), .CO(n38837));
    SB_LUT4 add_4966_14_lut (.I0(GND_net), .I1(n14489[11]), .I2(n962), 
            .I3(n38835), .O(n13768[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_14 (.CI(n38835), .I0(n14489[11]), .I1(n962), .CO(n38836));
    SB_LUT4 i32673_3_lut (.I0(n47804), .I1(n257[18]), .I2(n37_adj_4856), 
            .I3(GND_net), .O(n47805));   // verilog/motorControl.v(38[19:35])
    defparam i32673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4966_13_lut (.I0(GND_net), .I1(n14489[10]), .I2(n889), 
            .I3(n38834), .O(n13768[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_13 (.CI(n38834), .I0(n14489[10]), .I1(n889), .CO(n38835));
    SB_LUT4 add_4966_12_lut (.I0(GND_net), .I1(n14489[9]), .I2(n816), 
            .I3(n38833), .O(n13768[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_12 (.CI(n38833), .I0(n14489[9]), .I1(n816), .CO(n38834));
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32657_3_lut (.I0(n47805), .I1(n257[19]), .I2(n39_adj_4845), 
            .I3(GND_net), .O(n47789));   // verilog/motorControl.v(38[19:35])
    defparam i32657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4966_11_lut (.I0(GND_net), .I1(n14489[8]), .I2(n743), 
            .I3(n38832), .O(n13768[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n37723), .I0(GND_net), .I1(n1[20]), 
            .CO(n37724));
    SB_CARRY add_4966_11 (.CI(n38832), .I0(n14489[8]), .I1(n743), .CO(n38833));
    SB_CARRY add_12_3 (.CI(n37566), .I0(n106[1]), .I1(n155[1]), .CO(n37567));
    SB_LUT4 add_4966_10_lut (.I0(GND_net), .I1(n14489[7]), .I2(n670), 
            .I3(n38831), .O(n13768[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_10 (.CI(n38831), .I0(n14489[7]), .I1(n670), .CO(n38832));
    SB_LUT4 add_4966_9_lut (.I0(GND_net), .I1(n14489[6]), .I2(n597), .I3(n38830), 
            .O(n13768[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_9 (.CI(n38830), .I0(n14489[6]), .I1(n597), .CO(n38831));
    SB_LUT4 add_4966_8_lut (.I0(GND_net), .I1(n14489[5]), .I2(n524), .I3(n38829), 
            .O(n13768[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_8 (.CI(n38829), .I0(n14489[5]), .I1(n524), .CO(n38830));
    SB_LUT4 add_4966_7_lut (.I0(GND_net), .I1(n14489[4]), .I2(n451), .I3(n38828), 
            .O(n13768[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31793_4_lut (.I0(n43_adj_4854), .I1(n41_adj_4844), .I2(n39_adj_4845), 
            .I3(n47744), .O(n46924));
    defparam i31793_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4966_7 (.CI(n38828), .I0(n14489[4]), .I1(n451), .CO(n38829));
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4899));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32580_4_lut (.I0(n47623), .I1(n47526), .I2(n45_adj_4847), 
            .I3(n46922), .O(n47712));   // verilog/motorControl.v(38[19:35])
    defparam i32580_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4966_6_lut (.I0(GND_net), .I1(n14489[3]), .I2(n378), .I3(n38827), 
            .O(n13768[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_6 (.CI(n38827), .I0(n14489[3]), .I1(n378), .CO(n38828));
    SB_LUT4 i32643_3_lut (.I0(n47789), .I1(n257[20]), .I2(n41_adj_4844), 
            .I3(GND_net), .O(n40_adj_4900));   // verilog/motorControl.v(38[19:35])
    defparam i32643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4966_5_lut (.I0(GND_net), .I1(n14489[2]), .I2(n305), .I3(n38826), 
            .O(n13768[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_5 (.CI(n38826), .I0(n14489[2]), .I1(n305), .CO(n38827));
    SB_LUT4 i32582_4_lut (.I0(n40_adj_4900), .I1(n47712), .I2(n45_adj_4847), 
            .I3(n46924), .O(n47714));   // verilog/motorControl.v(38[19:35])
    defparam i32582_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_4966_4_lut (.I0(GND_net), .I1(n14489[1]), .I2(n232), .I3(n38825), 
            .O(n13768[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_4 (.CI(n38825), .I0(n14489[1]), .I1(n232), .CO(n38826));
    SB_LUT4 add_4966_3_lut (.I0(GND_net), .I1(n14489[0]), .I2(n159), .I3(n38824), 
            .O(n13768[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4966_3 (.CI(n38824), .I0(n14489[0]), .I1(n159), .CO(n38825));
    SB_LUT4 add_4966_2_lut (.I0(GND_net), .I1(n17), .I2(n86), .I3(GND_net), 
            .O(n13768[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4966_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32583_3_lut (.I0(n47714), .I1(duty_23__N_3772[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4729));   // verilog/motorControl.v(38[19:35])
    defparam i32583_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3772[0]), .I1(n257[0]), .I2(n256_adj_4729), 
            .I3(GND_net), .O(duty_23__N_3747[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4966_2 (.CI(GND_net), .I0(n17), .I1(n86), .CO(n38824));
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4902));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3747[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3771), .I3(GND_net), .O(duty_23__N_3648[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5227_10_lut (.I0(GND_net), .I1(n18209[7]), .I2(n700), 
            .I3(n38823), .O(n18029[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5227_9_lut (.I0(GND_net), .I1(n18209[6]), .I2(n627), .I3(n38822), 
            .O(n18029[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32625_3_lut (.I0(n47779), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_4903), .I3(GND_net), .O(n47757));   // verilog/motorControl.v(31[38:63])
    defparam i32625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4736));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5227_9 (.CI(n38822), .I0(n18209[6]), .I1(n627), .CO(n38823));
    SB_LUT4 add_5227_8_lut (.I0(GND_net), .I1(n18209[5]), .I2(n554), .I3(n38821), 
            .O(n18029[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4848));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5227_8 (.CI(n38821), .I0(n18209[5]), .I1(n554), .CO(n38822));
    SB_LUT4 add_5227_7_lut (.I0(GND_net), .I1(n18209[4]), .I2(n481), .I3(n38820), 
            .O(n18029[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4792), .I3(GND_net), 
            .O(n6_adj_4904));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_5227_7 (.CI(n38820), .I0(n18209[4]), .I1(n481), .CO(n38821));
    SB_LUT4 i32424_3_lut (.I0(n6_adj_4904), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4772), .I3(GND_net), .O(n47556));   // verilog/motorControl.v(31[38:63])
    defparam i32424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5227_6_lut (.I0(GND_net), .I1(n18209[3]), .I2(n408), .I3(n38819), 
            .O(n18029[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20001_2_lut (.I0(n28[15]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20001_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32425_3_lut (.I0(n47556), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4795), .I3(GND_net), .O(n47557));   // verilog/motorControl.v(31[38:63])
    defparam i32425_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5227_6 (.CI(n38819), .I0(n18209[3]), .I1(n408), .CO(n38820));
    SB_LUT4 add_5227_5_lut (.I0(GND_net), .I1(n18209[2]), .I2(n335), .I3(n38818), 
            .O(n18029[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i31884_4_lut (.I0(n43), .I1(n25_adj_4794), .I2(n23_adj_4795), 
            .I3(n47080), .O(n47015));
    defparam i31884_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5227_5 (.CI(n38818), .I0(n18209[2]), .I1(n335), .CO(n38819));
    SB_LUT4 add_5227_4_lut (.I0(GND_net), .I1(n18209[1]), .I2(n262), .I3(n38817), 
            .O(n18029[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_4 (.CI(n38817), .I0(n18209[1]), .I1(n262), .CO(n38818));
    SB_LUT4 add_5227_3_lut (.I0(GND_net), .I1(n18209[0]), .I2(n189), .I3(n38816), 
            .O(n18029[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32390_4_lut (.I0(n24_adj_4791), .I1(n8_adj_4785), .I2(n45), 
            .I3(n47013), .O(n47522));   // verilog/motorControl.v(31[38:63])
    defparam i32390_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32189_3_lut (.I0(n47557), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4794), .I3(GND_net), .O(n47321));   // verilog/motorControl.v(31[38:63])
    defparam i32189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31894_4_lut (.I0(n43), .I1(n41_adj_4905), .I2(n39_adj_4903), 
            .I3(n47752), .O(n47025));
    defparam i31894_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5227_3 (.CI(n38816), .I0(n18209[0]), .I1(n189), .CO(n38817));
    SB_LUT4 add_5227_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n18029[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n38816));
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5112_8 (.CI(n38496), .I0(n16869[5]), .I1(n539), .CO(n38497));
    SB_LUT4 add_5112_7_lut (.I0(GND_net), .I1(n16869[4]), .I2(n466), .I3(n38495), 
            .O(n16449[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32568_4_lut (.I0(n47321), .I1(n47522), .I2(n45), .I3(n47015), 
            .O(n47700));   // verilog/motorControl.v(31[38:63])
    defparam i32568_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5112_7 (.CI(n38495), .I0(n16869[4]), .I1(n466), .CO(n38496));
    SB_LUT4 add_5112_6_lut (.I0(GND_net), .I1(n16869[3]), .I2(n393), .I3(n38494), 
            .O(n16449[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20000_2_lut (.I0(n28[16]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20000_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n37722), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5112_6 (.CI(n38494), .I0(n16869[3]), .I1(n393), .CO(n38495));
    SB_LUT4 add_5002_19_lut (.I0(GND_net), .I1(n15136[16]), .I2(GND_net), 
            .I3(n38815), .O(n14489[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32197_3_lut (.I0(n47757), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4905), .I3(GND_net), .O(n47329));   // verilog/motorControl.v(31[38:63])
    defparam i32197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5112_5_lut (.I0(GND_net), .I1(n16869[2]), .I2(n320), .I3(n38493), 
            .O(n16449[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5002_18_lut (.I0(GND_net), .I1(n15136[15]), .I2(GND_net), 
            .I3(n38814), .O(n14489[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_18 (.CI(n38814), .I0(n15136[15]), .I1(GND_net), 
            .CO(n38815));
    SB_LUT4 add_5002_17_lut (.I0(GND_net), .I1(n15136[14]), .I2(GND_net), 
            .I3(n38813), .O(n14489[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_17 (.CI(n38813), .I0(n15136[14]), .I1(GND_net), 
            .CO(n38814));
    SB_LUT4 add_5002_16_lut (.I0(GND_net), .I1(n15136[13]), .I2(n1111), 
            .I3(n38812), .O(n14489[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_16 (.CI(n38812), .I0(n15136[13]), .I1(n1111), .CO(n38813));
    SB_LUT4 add_5002_15_lut (.I0(GND_net), .I1(n15136[12]), .I2(n1038), 
            .I3(n38811), .O(n14489[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_15 (.CI(n38811), .I0(n15136[12]), .I1(n1038), .CO(n38812));
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5002_14_lut (.I0(GND_net), .I1(n15136[11]), .I2(n965), 
            .I3(n38810), .O(n14489[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5002_14 (.CI(n38810), .I0(n15136[11]), .I1(n965), .CO(n38811));
    SB_LUT4 add_5002_13_lut (.I0(GND_net), .I1(n15136[10]), .I2(n892), 
            .I3(n38809), .O(n14489[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_13 (.CI(n38809), .I0(n15136[10]), .I1(n892), .CO(n38810));
    SB_LUT4 add_5002_12_lut (.I0(GND_net), .I1(n15136[9]), .I2(n819), 
            .I3(n38808), .O(n14489[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_12 (.CI(n38808), .I0(n15136[9]), .I1(n819), .CO(n38809));
    SB_LUT4 i19999_2_lut (.I0(n28[17]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19999_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5002_11_lut (.I0(GND_net), .I1(n15136[8]), .I2(n746), 
            .I3(n38807), .O(n14489[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32570_4_lut (.I0(n47329), .I1(n47700), .I2(n45), .I3(n47025), 
            .O(n47702));   // verilog/motorControl.v(31[38:63])
    defparam i32570_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5002_11 (.CI(n38807), .I0(n15136[8]), .I1(n746), .CO(n38808));
    SB_LUT4 add_5002_10_lut (.I0(GND_net), .I1(n15136[7]), .I2(n673), 
            .I3(n38806), .O(n14489[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3772[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_10 (.CI(n38806), .I0(n15136[7]), .I1(n673), .CO(n38807));
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5002_9_lut (.I0(GND_net), .I1(n15136[6]), .I2(n600), .I3(n38805), 
            .O(n14489[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n37722), .I0(GND_net), .I1(n1[19]), 
            .CO(n37723));
    SB_CARRY add_5002_9 (.CI(n38805), .I0(n15136[6]), .I1(n600), .CO(n38806));
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5002_8_lut (.I0(GND_net), .I1(n15136[5]), .I2(n527), .I3(n38804), 
            .O(n14489[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_8 (.CI(n38804), .I0(n15136[5]), .I1(n527), .CO(n38805));
    SB_LUT4 add_5002_7_lut (.I0(GND_net), .I1(n15136[4]), .I2(n454), .I3(n38803), 
            .O(n14489[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_7 (.CI(n38803), .I0(n15136[4]), .I1(n454), .CO(n38804));
    SB_LUT4 add_5002_6_lut (.I0(GND_net), .I1(n15136[3]), .I2(n381), .I3(n38802), 
            .O(n14489[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_6 (.CI(n38802), .I0(n15136[3]), .I1(n381), .CO(n38803));
    SB_LUT4 add_5002_5_lut (.I0(GND_net), .I1(n15136[2]), .I2(n308), .I3(n38801), 
            .O(n14489[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_5 (.CI(n38801), .I0(n15136[2]), .I1(n308), .CO(n38802));
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5002_4_lut (.I0(GND_net), .I1(n15136[1]), .I2(n235), .I3(n38800), 
            .O(n14489[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_4 (.CI(n38800), .I0(n15136[1]), .I1(n235), .CO(n38801));
    SB_LUT4 add_5002_3_lut (.I0(GND_net), .I1(n15136[0]), .I2(n162), .I3(n38799), 
            .O(n14489[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_3 (.CI(n38799), .I0(n15136[0]), .I1(n162), .CO(n38800));
    SB_LUT4 add_5002_2_lut (.I0(GND_net), .I1(n20_adj_4712), .I2(n89), 
            .I3(GND_net), .O(n14489[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5002_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5002_2 (.CI(GND_net), .I0(n20_adj_4712), .I1(n89), .CO(n38799));
    SB_LUT4 add_5036_18_lut (.I0(GND_net), .I1(n15713[15]), .I2(GND_net), 
            .I3(n38798), .O(n15136[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5036_17_lut (.I0(GND_net), .I1(n15713[14]), .I2(GND_net), 
            .I3(n38797), .O(n15136[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_17 (.CI(n38797), .I0(n15713[14]), .I1(GND_net), 
            .CO(n38798));
    SB_LUT4 add_5036_16_lut (.I0(GND_net), .I1(n15713[13]), .I2(n1114), 
            .I3(n38796), .O(n15136[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_16 (.CI(n38796), .I0(n15713[13]), .I1(n1114), .CO(n38797));
    SB_LUT4 add_5036_15_lut (.I0(GND_net), .I1(n15713[12]), .I2(n1041), 
            .I3(n38795), .O(n15136[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_15 (.CI(n38795), .I0(n15713[12]), .I1(n1041), .CO(n38796));
    SB_LUT4 add_5036_14_lut (.I0(GND_net), .I1(n15713[11]), .I2(n968), 
            .I3(n38794), .O(n15136[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_14 (.CI(n38794), .I0(n15713[11]), .I1(n968), .CO(n38795));
    SB_LUT4 add_5036_13_lut (.I0(GND_net), .I1(n15713[10]), .I2(n895), 
            .I3(n38793), .O(n15136[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_13 (.CI(n38793), .I0(n15713[10]), .I1(n895), .CO(n38794));
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4908));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_5036_12_lut (.I0(GND_net), .I1(n15713[9]), .I2(n822), 
            .I3(n38792), .O(n15136[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_12 (.CI(n38792), .I0(n15713[9]), .I1(n822), .CO(n38793));
    SB_LUT4 add_5036_11_lut (.I0(GND_net), .I1(n15713[8]), .I2(n749_adj_4711), 
            .I3(n38791), .O(n15136[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_11 (.CI(n38791), .I0(n15713[8]), .I1(n749_adj_4711), 
            .CO(n38792));
    SB_LUT4 add_5036_10_lut (.I0(GND_net), .I1(n15713[7]), .I2(n676_adj_4710), 
            .I3(n38790), .O(n15136[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4909));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5036_10 (.CI(n38790), .I0(n15713[7]), .I1(n676_adj_4710), 
            .CO(n38791));
    SB_LUT4 add_5036_9_lut (.I0(GND_net), .I1(n15713[6]), .I2(n603), .I3(n38789), 
            .O(n15136[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_9 (.CI(n38789), .I0(n15713[6]), .I1(n603), .CO(n38790));
    SB_LUT4 add_5036_8_lut (.I0(GND_net), .I1(n15713[5]), .I2(n530), .I3(n38788), 
            .O(n15136[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_8 (.CI(n38788), .I0(n15713[5]), .I1(n530), .CO(n38789));
    SB_LUT4 add_5036_7_lut (.I0(GND_net), .I1(n15713[4]), .I2(n457), .I3(n38787), 
            .O(n15136[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_7 (.CI(n38787), .I0(n15713[4]), .I1(n457), .CO(n38788));
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5112_5 (.CI(n38493), .I0(n16869[2]), .I1(n320), .CO(n38494));
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5036_6_lut (.I0(GND_net), .I1(n15713[3]), .I2(n384), .I3(n38786), 
            .O(n15136[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_6 (.CI(n38786), .I0(n15713[3]), .I1(n384), .CO(n38787));
    SB_LUT4 add_5036_5_lut (.I0(GND_net), .I1(n15713[2]), .I2(n311), .I3(n38785), 
            .O(n15136[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5112_4_lut (.I0(GND_net), .I1(n16869[1]), .I2(n247), .I3(n38492), 
            .O(n16449[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23683_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n37160), .I3(n18673[0]), .O(n4_adj_4911));   // verilog/motorControl.v(34[25:36])
    defparam i23683_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(n18673[0]), .I3(n37160), .O(n18649[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i23670_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n18649[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23670_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_CARRY add_5036_5 (.CI(n38785), .I0(n15713[2]), .I1(n311), .CO(n38786));
    SB_LUT4 i23672_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [20]), .I3(\Ki[1] ), 
            .O(n37160));   // verilog/motorControl.v(34[25:36])
    defparam i23672_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n37721), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23767_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n4_adj_4912), .I3(n18609[1]), .O(n6_adj_4913));   // verilog/motorControl.v(34[25:36])
    defparam i23767_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_5036_4_lut (.I0(GND_net), .I1(n15713[1]), .I2(n238), .I3(n38784), 
            .O(n15136[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5036_4 (.CI(n38784), .I0(n15713[1]), .I1(n238), .CO(n38785));
    SB_LUT4 add_5036_3_lut (.I0(GND_net), .I1(n15713[0]), .I2(n165), .I3(n38783), 
            .O(n15136[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1544 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n18609[1]), .I3(n4_adj_4912), .O(n18549[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1544.LUT_INIT = 16'h8778;
    SB_CARRY add_5036_3 (.CI(n38783), .I0(n15713[0]), .I1(n165), .CO(n38784));
    SB_LUT4 add_5036_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n15136[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5036_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4730));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5036_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n38783));
    SB_LUT4 i2_3_lut_4_lut_adj_1545 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n18609[0]), .I3(n37242), .O(n18549[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1545.LUT_INIT = 16'h8778;
    SB_LUT4 i23759_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(n37242), .I3(n18609[0]), .O(n4_adj_4912));   // verilog/motorControl.v(34[25:36])
    defparam i23759_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i23746_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n18549[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23746_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_5244_9_lut (.I0(GND_net), .I1(n18353[6]), .I2(n630), .I3(n38782), 
            .O(n18209[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5112_4 (.CI(n38492), .I0(n16869[1]), .I1(n247), .CO(n38493));
    SB_LUT4 i23748_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), .I3(\Ki[1] ), 
            .O(n37242));   // verilog/motorControl.v(34[25:36])
    defparam i23748_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4727));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5244_8_lut (.I0(GND_net), .I1(n18353[5]), .I2(n557), .I3(n38781), 
            .O(n18209[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5244_8 (.CI(n38781), .I0(n18353[5]), .I1(n557), .CO(n38782));
    SB_LUT4 add_5244_7_lut (.I0(GND_net), .I1(n18353[4]), .I2(n484), .I3(n38780), 
            .O(n18209[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4726));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n37566));
    SB_CARRY add_5244_7 (.CI(n38780), .I0(n18353[4]), .I1(n484), .CO(n38781));
    SB_LUT4 add_5244_6_lut (.I0(GND_net), .I1(n18353[3]), .I2(n411), .I3(n38779), 
            .O(n18209[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5112_3_lut (.I0(GND_net), .I1(n16869[0]), .I2(n174), .I3(n38491), 
            .O(n16449[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i32432_3_lut (.I0(n4_adj_4908), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n47564));   // verilog/motorControl.v(31[10:34])
    defparam i32432_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5112_3 (.CI(n38491), .I0(n16869[0]), .I1(n174), .CO(n38492));
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5244_6 (.CI(n38779), .I0(n18353[3]), .I1(n411), .CO(n38780));
    SB_LUT4 add_5112_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n16449[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5112_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5244_5_lut (.I0(GND_net), .I1(n18353[2]), .I2(n338), .I3(n38778), 
            .O(n18209[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5244_5 (.CI(n38778), .I0(n18353[2]), .I1(n338), .CO(n38779));
    SB_LUT4 add_5244_4_lut (.I0(GND_net), .I1(n18353[1]), .I2(n265), .I3(n38777), 
            .O(n18209[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5244_4 (.CI(n38777), .I0(n18353[1]), .I1(n265), .CO(n38778));
    SB_LUT4 i32433_3_lut (.I0(n47564), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n47565));   // verilog/motorControl.v(31[10:34])
    defparam i32433_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4790));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4914));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4915));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31980_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n48891), 
            .I2(IntegralLimit[16]), .I3(n47374), .O(n47111));
    defparam i31980_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4724));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1546 (.I0(n62), .I1(n131), .I2(n18649[0]), 
            .I3(n204), .O(n18609[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1546.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4789));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5244_3_lut (.I0(GND_net), .I1(n18353[0]), .I2(n192), .I3(n38776), 
            .O(n18209[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5244_3 (.CI(n38776), .I0(n18353[0]), .I1(n192), .CO(n38777));
    SB_LUT4 add_5244_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n18209[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5244_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23721_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n18649[0]), 
            .O(n4_adj_4916));   // verilog/motorControl.v(34[25:36])
    defparam i23721_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i20015_2_lut (.I0(n28[1]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20015_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32536_4_lut (.I0(n30), .I1(n10_adj_4798), .I2(n48914), .I3(n47109), 
            .O(n47668));   // verilog/motorControl.v(31[10:34])
    defparam i32536_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5244_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n38776));
    SB_LUT4 i32181_3_lut (.I0(n47565), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n47313));   // verilog/motorControl.v(31[10:34])
    defparam i32181_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5068_17_lut (.I0(GND_net), .I1(n16224[14]), .I2(GND_net), 
            .I3(n38775), .O(n15713[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4787));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5068_16_lut (.I0(GND_net), .I1(n16224[13]), .I2(n1117_adj_4709), 
            .I3(n38774), .O(n15713[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_16 (.CI(n38774), .I0(n16224[13]), .I1(n1117_adj_4709), 
            .CO(n38775));
    SB_LUT4 add_5068_15_lut (.I0(GND_net), .I1(n16224[12]), .I2(n1044), 
            .I3(n38773), .O(n15713[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_15 (.CI(n38773), .I0(n16224[12]), .I1(n1044), .CO(n38774));
    SB_LUT4 add_5068_14_lut (.I0(GND_net), .I1(n16224[11]), .I2(n971), 
            .I3(n38772), .O(n15713[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_14 (.CI(n38772), .I0(n16224[11]), .I1(n971), .CO(n38773));
    SB_LUT4 add_5068_13_lut (.I0(GND_net), .I1(n16224[10]), .I2(n898), 
            .I3(n38771), .O(n15713[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_13 (.CI(n38771), .I0(n16224[10]), .I1(n898), .CO(n38772));
    SB_LUT4 add_5068_12_lut (.I0(GND_net), .I1(n16224[9]), .I2(n825), 
            .I3(n38770), .O(n15713[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4783));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n37721), .I0(GND_net), .I1(n1[18]), 
            .CO(n37722));
    SB_CARRY add_5068_12 (.CI(n38770), .I0(n16224[9]), .I1(n825), .CO(n38771));
    SB_LUT4 add_5068_11_lut (.I0(GND_net), .I1(n16224[8]), .I2(n752), 
            .I3(n38769), .O(n15713[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5112_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n38491));
    SB_LUT4 i23889_3_lut_4_lut (.I0(\Kp[3] ), .I1(n28[18]), .I2(n4_adj_4917), 
            .I3(n18633[1]), .O(n6_adj_4918));   // verilog/motorControl.v(34[16:22])
    defparam i23889_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_5068_11 (.CI(n38769), .I0(n16224[8]), .I1(n752), .CO(n38770));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n37720), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5068_10_lut (.I0(GND_net), .I1(n16224[7]), .I2(n679), 
            .I3(n38768), .O(n15713[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_10 (.CI(n38768), .I0(n16224[7]), .I1(n679), .CO(n38769));
    SB_CARRY unary_minus_16_add_3_19 (.CI(n37720), .I0(GND_net), .I1(n1[17]), 
            .CO(n37721));
    SB_LUT4 add_5068_9_lut (.I0(GND_net), .I1(n16224[6]), .I2(n606), .I3(n38767), 
            .O(n15713[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_9 (.CI(n38767), .I0(n16224[6]), .I1(n606), .CO(n38768));
    SB_LUT4 add_5266_8_lut (.I0(GND_net), .I1(n18513[5]), .I2(n560), .I3(n38490), 
            .O(n18416[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5266_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5068_8_lut (.I0(GND_net), .I1(n16224[5]), .I2(n533), .I3(n38766), 
            .O(n15713[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_8 (.CI(n38766), .I0(n16224[5]), .I1(n533), .CO(n38767));
    SB_LUT4 add_5068_7_lut (.I0(GND_net), .I1(n16224[4]), .I2(n460), .I3(n38765), 
            .O(n15713[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_7 (.CI(n38765), .I0(n16224[4]), .I1(n460), .CO(n38766));
    SB_LUT4 add_5068_6_lut (.I0(GND_net), .I1(n16224[3]), .I2(n387), .I3(n38764), 
            .O(n15713[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n37719), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_6 (.CI(n38764), .I0(n16224[3]), .I1(n387), .CO(n38765));
    SB_CARRY unary_minus_16_add_3_18 (.CI(n37719), .I0(GND_net), .I1(n1[16]), 
            .CO(n37720));
    SB_LUT4 add_5068_5_lut (.I0(GND_net), .I1(n16224[2]), .I2(n314), .I3(n38763), 
            .O(n15713[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_5 (.CI(n38763), .I0(n16224[2]), .I1(n314), .CO(n38764));
    SB_LUT4 i2_3_lut_4_lut_adj_1547 (.I0(\Kp[3] ), .I1(n28[18]), .I2(n18633[1]), 
            .I3(n4_adj_4917), .O(n18584[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1547.LUT_INIT = 16'h8778;
    SB_LUT4 add_5068_4_lut (.I0(GND_net), .I1(n16224[1]), .I2(n241), .I3(n38762), 
            .O(n15713[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_4 (.CI(n38762), .I0(n16224[1]), .I1(n241), .CO(n38763));
    SB_LUT4 add_5068_3_lut (.I0(GND_net), .I1(n16224[0]), .I2(n168), .I3(n38761), 
            .O(n15713[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_3 (.CI(n38761), .I0(n16224[0]), .I1(n168), .CO(n38762));
    SB_LUT4 add_5068_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n15713[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5068_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n37718), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5068_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n38761));
    SB_LUT4 add_5266_7_lut (.I0(GND_net), .I1(n18513[4]), .I2(n487), .I3(n38489), 
            .O(n18416[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5266_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n37718), .I0(GND_net), .I1(n1[15]), 
            .CO(n37719));
    SB_CARRY add_5266_7 (.CI(n38489), .I0(n18513[4]), .I1(n487), .CO(n38490));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n37717), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n37717), .I0(GND_net), .I1(n1[14]), 
            .CO(n37718));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n37716), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n37716), .I0(GND_net), .I1(n1[13]), 
            .CO(n37717));
    SB_LUT4 add_5098_16_lut (.I0(GND_net), .I1(n16673[13]), .I2(n1120_adj_4920), 
            .I3(n38760), .O(n16224[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n37715), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5266_6_lut (.I0(GND_net), .I1(n18513[3]), .I2(n414), .I3(n38488), 
            .O(n18416[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5266_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n37715), .I0(GND_net), .I1(n1[12]), 
            .CO(n37716));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n37714), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5266_6 (.CI(n38488), .I0(n18513[3]), .I1(n414), .CO(n38489));
    SB_LUT4 add_5098_15_lut (.I0(GND_net), .I1(n16673[12]), .I2(n1047_adj_4923), 
            .I3(n38759), .O(n16224[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_15 (.CI(n38759), .I0(n16673[12]), .I1(n1047_adj_4923), 
            .CO(n38760));
    SB_LUT4 add_5266_5_lut (.I0(GND_net), .I1(n18513[2]), .I2(n341), .I3(n38487), 
            .O(n18416[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5266_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1548 (.I0(\Kp[2] ), .I1(n28[18]), .I2(n18633[0]), 
            .I3(n37374), .O(n18584[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1548.LUT_INIT = 16'h8778;
    SB_LUT4 i23881_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[18]), .I2(n37374), 
            .I3(n18633[0]), .O(n4_adj_4917));   // verilog/motorControl.v(34[16:22])
    defparam i23881_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i23868_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n18584[0]));   // verilog/motorControl.v(34[16:22])
    defparam i23868_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i23870_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n37374));   // verilog/motorControl.v(34[16:22])
    defparam i23870_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_5098_14_lut (.I0(GND_net), .I1(n16673[11]), .I2(n974_adj_4924), 
            .I3(n38758), .O(n16224[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5266_5 (.CI(n38487), .I0(n18513[2]), .I1(n341), .CO(n38488));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n37714), .I0(GND_net), .I1(n1[11]), 
            .CO(n37715));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n37713), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_14 (.CI(n38758), .I0(n16673[11]), .I1(n974_adj_4924), 
            .CO(n38759));
    SB_LUT4 add_5098_13_lut (.I0(GND_net), .I1(n16673[10]), .I2(n901_adj_4926), 
            .I3(n38757), .O(n16224[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4782));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5098_13 (.CI(n38757), .I0(n16673[10]), .I1(n901_adj_4926), 
            .CO(n38758));
    SB_LUT4 add_5098_12_lut (.I0(GND_net), .I1(n16673[9]), .I2(n828_adj_4927), 
            .I3(n38756), .O(n16224[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_12 (.CI(n38756), .I0(n16673[9]), .I1(n828_adj_4927), 
            .CO(n38757));
    SB_LUT4 add_5098_11_lut (.I0(GND_net), .I1(n16673[8]), .I2(n755_adj_4928), 
            .I3(n38755), .O(n16224[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_11 (.CI(n38755), .I0(n16673[8]), .I1(n755_adj_4928), 
            .CO(n38756));
    SB_LUT4 add_5098_10_lut (.I0(GND_net), .I1(n16673[7]), .I2(n682_adj_4929), 
            .I3(n38754), .O(n16224[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_10 (.CI(n38754), .I0(n16673[7]), .I1(n682_adj_4929), 
            .CO(n38755));
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4781));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5266_4_lut (.I0(GND_net), .I1(n18513[1]), .I2(n268_adj_4930), 
            .I3(n38486), .O(n18416[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5266_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4931));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4932));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23805_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[20]), .I2(n37292), 
            .I3(n18681[0]), .O(n4_adj_4934));   // verilog/motorControl.v(34[16:22])
    defparam i23805_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1549 (.I0(\Kp[2] ), .I1(n28[20]), .I2(n18681[0]), 
            .I3(n37292), .O(n18664[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1549.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4778));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5098_9_lut (.I0(GND_net), .I1(n16673[6]), .I2(n609_adj_4935), 
            .I3(n38753), .O(n16224[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n37713), .I0(GND_net), .I1(n1[10]), 
            .CO(n37714));
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5098_9 (.CI(n38753), .I0(n16673[6]), .I1(n609_adj_4935), 
            .CO(n38754));
    SB_LUT4 add_5098_8_lut (.I0(GND_net), .I1(n16673[5]), .I2(n536_adj_4936), 
            .I3(n38752), .O(n16224[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_8 (.CI(n38752), .I0(n16673[5]), .I1(n536_adj_4936), 
            .CO(n38753));
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4937));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5098_7_lut (.I0(GND_net), .I1(n16673[4]), .I2(n463_adj_4938), 
            .I3(n38751), .O(n16224[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_7 (.CI(n38751), .I0(n16673[4]), .I1(n463_adj_4938), 
            .CO(n38752));
    SB_LUT4 add_5098_6_lut (.I0(GND_net), .I1(n16673[3]), .I2(n390_adj_4939), 
            .I3(n38750), .O(n16224[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut_adj_1550 (.I0(n62_adj_4940), .I1(n131_adj_4941), 
            .I2(n18664[0]), .I3(n204_adj_4942), .O(n18633[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1550.LUT_INIT = 16'h8778;
    SB_CARRY add_5098_6 (.CI(n38750), .I0(n16673[3]), .I1(n390_adj_4939), 
            .CO(n38751));
    SB_LUT4 add_5098_5_lut (.I0(GND_net), .I1(n16673[2]), .I2(n317_adj_4943), 
            .I3(n38749), .O(n16224[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_5 (.CI(n38749), .I0(n16673[2]), .I1(n317_adj_4943), 
            .CO(n38750));
    SB_LUT4 add_5098_4_lut (.I0(GND_net), .I1(n16673[1]), .I2(n244_adj_4944), 
            .I3(n38748), .O(n16224[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_4 (.CI(n38748), .I0(n16673[1]), .I1(n244_adj_4944), 
            .CO(n38749));
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5098_3_lut (.I0(GND_net), .I1(n16673[0]), .I2(n171_adj_4946), 
            .I3(n38747), .O(n16224[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5098_3 (.CI(n38747), .I0(n16673[0]), .I1(n171_adj_4946), 
            .CO(n38748));
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4947));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5098_2_lut (.I0(GND_net), .I1(n29_adj_4948), .I2(n98_adj_4949), 
            .I3(GND_net), .O(n16224[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5098_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4951));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5098_2 (.CI(GND_net), .I0(n29_adj_4948), .I1(n98_adj_4949), 
            .CO(n38747));
    SB_CARRY add_5266_4 (.CI(n38486), .I0(n18513[1]), .I1(n268_adj_4930), 
            .CO(n38487));
    SB_LUT4 add_5259_8_lut (.I0(GND_net), .I1(n18465[5]), .I2(n560_adj_4952), 
            .I3(n38746), .O(n18353[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4954));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5266_3_lut (.I0(GND_net), .I1(n18513[0]), .I2(n195_adj_4955), 
            .I3(n38485), .O(n18416[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5266_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5259_7_lut (.I0(GND_net), .I1(n18465[4]), .I2(n487_adj_4956), 
            .I3(n38745), .O(n18353[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_7 (.CI(n38745), .I0(n18465[4]), .I1(n487_adj_4956), 
            .CO(n38746));
    SB_LUT4 add_5259_6_lut (.I0(GND_net), .I1(n18465[3]), .I2(n414_adj_4957), 
            .I3(n38744), .O(n18353[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_6 (.CI(n38744), .I0(n18465[3]), .I1(n414_adj_4957), 
            .CO(n38745));
    SB_CARRY add_5266_3 (.CI(n38485), .I0(n18513[0]), .I1(n195_adj_4955), 
            .CO(n38486));
    SB_LUT4 add_5259_5_lut (.I0(GND_net), .I1(n18465[2]), .I2(n341_adj_4958), 
            .I3(n38743), .O(n18353[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5266_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n18416[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5266_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_5 (.CI(n38743), .I0(n18465[2]), .I1(n341_adj_4958), 
            .CO(n38744));
    SB_CARRY add_5266_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n38485));
    SB_LUT4 add_5259_4_lut (.I0(GND_net), .I1(n18465[1]), .I2(n268_adj_4959), 
            .I3(n38742), .O(n18353[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_4 (.CI(n38742), .I0(n18465[1]), .I1(n268_adj_4959), 
            .CO(n38743));
    SB_LUT4 add_5139_14_lut (.I0(GND_net), .I1(n17233[11]), .I2(n980), 
            .I3(n38484), .O(n16869[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5259_3_lut (.I0(GND_net), .I1(n18465[0]), .I2(n195_adj_4960), 
            .I3(n38741), .O(n18353[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_13_lut (.I0(GND_net), .I1(n17233[10]), .I2(n907), 
            .I3(n38483), .O(n16869[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5259_3 (.CI(n38741), .I0(n18465[0]), .I1(n195_adj_4960), 
            .CO(n38742));
    SB_LUT4 add_5259_2_lut (.I0(GND_net), .I1(n53_adj_4961), .I2(n122_adj_4962), 
            .I3(GND_net), .O(n18353[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5259_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_13 (.CI(n38483), .I0(n17233[10]), .I1(n907), .CO(n38484));
    SB_CARRY add_5259_2 (.CI(GND_net), .I0(n53_adj_4961), .I1(n122_adj_4962), 
            .CO(n38741));
    SB_LUT4 add_5126_15_lut (.I0(GND_net), .I1(n17064[12]), .I2(n1050_adj_4963), 
            .I3(n38740), .O(n16673[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5126_14_lut (.I0(GND_net), .I1(n17064[11]), .I2(n977_adj_4964), 
            .I3(n38739), .O(n16673[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_14 (.CI(n38739), .I0(n17064[11]), .I1(n977_adj_4964), 
            .CO(n38740));
    SB_LUT4 add_5126_13_lut (.I0(GND_net), .I1(n17064[10]), .I2(n904_adj_4965), 
            .I3(n38738), .O(n16673[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_13 (.CI(n38738), .I0(n17064[10]), .I1(n904_adj_4965), 
            .CO(n38739));
    SB_LUT4 add_5126_12_lut (.I0(GND_net), .I1(n17064[9]), .I2(n831_adj_4966), 
            .I3(n38737), .O(n16673[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_12 (.CI(n38737), .I0(n17064[9]), .I1(n831_adj_4966), 
            .CO(n38738));
    SB_LUT4 add_5126_11_lut (.I0(GND_net), .I1(n17064[8]), .I2(n758_adj_4967), 
            .I3(n38736), .O(n16673[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5126_11 (.CI(n38736), .I0(n17064[8]), .I1(n758_adj_4967), 
            .CO(n38737));
    SB_LUT4 add_5126_10_lut (.I0(GND_net), .I1(n17064[7]), .I2(n685_adj_4969), 
            .I3(n38735), .O(n16673[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_10 (.CI(n38735), .I0(n17064[7]), .I1(n685_adj_4969), 
            .CO(n38736));
    SB_LUT4 add_5126_9_lut (.I0(GND_net), .I1(n17064[6]), .I2(n612_adj_4970), 
            .I3(n38734), .O(n16673[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_9 (.CI(n38734), .I0(n17064[6]), .I1(n612_adj_4970), 
            .CO(n38735));
    SB_LUT4 add_5126_8_lut (.I0(GND_net), .I1(n17064[5]), .I2(n539_adj_4971), 
            .I3(n38733), .O(n16673[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_8 (.CI(n38733), .I0(n17064[5]), .I1(n539_adj_4971), 
            .CO(n38734));
    SB_LUT4 add_5126_7_lut (.I0(GND_net), .I1(n17064[4]), .I2(n466_adj_4972), 
            .I3(n38732), .O(n16673[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_7 (.CI(n38732), .I0(n17064[4]), .I1(n466_adj_4972), 
            .CO(n38733));
    SB_LUT4 add_5126_6_lut (.I0(GND_net), .I1(n17064[3]), .I2(n393_adj_4973), 
            .I3(n38731), .O(n16673[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_6 (.CI(n38731), .I0(n17064[3]), .I1(n393_adj_4973), 
            .CO(n38732));
    SB_LUT4 add_5126_5_lut (.I0(GND_net), .I1(n17064[2]), .I2(n320_adj_4974), 
            .I3(n38730), .O(n16673[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_5 (.CI(n38730), .I0(n17064[2]), .I1(n320_adj_4974), 
            .CO(n38731));
    SB_LUT4 add_5126_4_lut (.I0(GND_net), .I1(n17064[1]), .I2(n247_adj_4975), 
            .I3(n38729), .O(n16673[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_4 (.CI(n38729), .I0(n17064[1]), .I1(n247_adj_4975), 
            .CO(n38730));
    SB_LUT4 add_5126_3_lut (.I0(GND_net), .I1(n17064[0]), .I2(n174_adj_4976), 
            .I3(n38728), .O(n16673[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_3 (.CI(n38728), .I0(n17064[0]), .I1(n174_adj_4976), 
            .CO(n38729));
    SB_LUT4 add_5126_2_lut (.I0(GND_net), .I1(n32_adj_4977), .I2(n101_adj_4978), 
            .I3(GND_net), .O(n16673[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5126_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5126_2 (.CI(GND_net), .I0(n32_adj_4977), .I1(n101_adj_4978), 
            .CO(n38728));
    SB_LUT4 add_5152_14_lut (.I0(GND_net), .I1(n17401[11]), .I2(n980_adj_4979), 
            .I3(n38727), .O(n17064[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_12_lut (.I0(GND_net), .I1(n17233[9]), .I2(n834), 
            .I3(n38482), .O(n16869[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_13_lut (.I0(GND_net), .I1(n17401[10]), .I2(n907_adj_4980), 
            .I3(n38726), .O(n17064[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_13 (.CI(n38726), .I0(n17401[10]), .I1(n907_adj_4980), 
            .CO(n38727));
    SB_LUT4 add_5152_12_lut (.I0(GND_net), .I1(n17401[9]), .I2(n834_adj_4981), 
            .I3(n38725), .O(n17064[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_12 (.CI(n38725), .I0(n17401[9]), .I1(n834_adj_4981), 
            .CO(n38726));
    SB_CARRY add_5139_12 (.CI(n38482), .I0(n17233[9]), .I1(n834), .CO(n38483));
    SB_LUT4 add_5152_11_lut (.I0(GND_net), .I1(n17401[8]), .I2(n761), 
            .I3(n38724), .O(n17064[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n37712), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_11_lut (.I0(GND_net), .I1(n17233[8]), .I2(n761_adj_4983), 
            .I3(n38481), .O(n16869[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_11 (.CI(n38481), .I0(n17233[8]), .I1(n761_adj_4983), 
            .CO(n38482));
    SB_CARRY unary_minus_16_add_3_11 (.CI(n37712), .I0(GND_net), .I1(n1[9]), 
            .CO(n37713));
    SB_CARRY add_5152_11 (.CI(n38724), .I0(n17401[8]), .I1(n761), .CO(n38725));
    SB_LUT4 add_5139_10_lut (.I0(GND_net), .I1(n17233[7]), .I2(n688), 
            .I3(n38480), .O(n16869[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_10 (.CI(n38480), .I0(n17233[7]), .I1(n688), .CO(n38481));
    SB_LUT4 add_5139_9_lut (.I0(GND_net), .I1(n17233[6]), .I2(n615), .I3(n38479), 
            .O(n16869[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5152_10_lut (.I0(GND_net), .I1(n17401[7]), .I2(n688_adj_4985), 
            .I3(n38723), .O(n17064[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_10 (.CI(n38723), .I0(n17401[7]), .I1(n688_adj_4985), 
            .CO(n38724));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n37711), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_9_lut (.I0(GND_net), .I1(n17401[6]), .I2(n615_adj_4987), 
            .I3(n38722), .O(n17064[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_9 (.CI(n38479), .I0(n17233[6]), .I1(n615), .CO(n38480));
    SB_LUT4 i32634_4_lut (.I0(n47313), .I1(n47668), .I2(n48914), .I3(n47111), 
            .O(n47766));   // verilog/motorControl.v(31[10:34])
    defparam i32634_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5152_9 (.CI(n38722), .I0(n17401[6]), .I1(n615_adj_4987), 
            .CO(n38723));
    SB_LUT4 i23835_3_lut_4_lut (.I0(n62_adj_4940), .I1(n131_adj_4941), .I2(n204_adj_4942), 
            .I3(n18664[0]), .O(n4_adj_4988));   // verilog/motorControl.v(34[16:22])
    defparam i23835_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4989));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n37711), .I0(GND_net), .I1(n1[8]), 
            .CO(n37712));
    SB_LUT4 add_5139_8_lut (.I0(GND_net), .I1(n17233[5]), .I2(n542), .I3(n38478), 
            .O(n16869[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_8 (.CI(n38478), .I0(n17233[5]), .I1(n542), .CO(n38479));
    SB_LUT4 add_5139_7_lut (.I0(GND_net), .I1(n17233[4]), .I2(n469), .I3(n38477), 
            .O(n16869[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_7 (.CI(n38477), .I0(n17233[4]), .I1(n469), .CO(n38478));
    SB_LUT4 add_5139_6_lut (.I0(GND_net), .I1(n17233[3]), .I2(n396), .I3(n38476), 
            .O(n16869[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n37710), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_6 (.CI(n38476), .I0(n17233[3]), .I1(n396), .CO(n38477));
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4991));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5152_8_lut (.I0(GND_net), .I1(n17401[5]), .I2(n542_adj_4992), 
            .I3(n38721), .O(n17064[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_8 (.CI(n38721), .I0(n17401[5]), .I1(n542_adj_4992), 
            .CO(n38722));
    SB_LUT4 add_5152_7_lut (.I0(GND_net), .I1(n17401[4]), .I2(n469_adj_4993), 
            .I3(n38720), .O(n17064[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_5_lut (.I0(GND_net), .I1(n17233[2]), .I2(n323), .I3(n38475), 
            .O(n16869[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_7 (.CI(n38720), .I0(n17401[4]), .I1(n469_adj_4993), 
            .CO(n38721));
    SB_LUT4 add_5152_6_lut (.I0(GND_net), .I1(n17401[3]), .I2(n396_adj_4994), 
            .I3(n38719), .O(n17064[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_5 (.CI(n38475), .I0(n17233[2]), .I1(n323), .CO(n38476));
    SB_CARRY add_5152_6 (.CI(n38719), .I0(n17401[3]), .I1(n396_adj_4994), 
            .CO(n38720));
    SB_LUT4 add_5152_5_lut (.I0(GND_net), .I1(n17401[2]), .I2(n323_adj_4995), 
            .I3(n38718), .O(n17064[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_5 (.CI(n38718), .I0(n17401[2]), .I1(n323_adj_4995), 
            .CO(n38719));
    SB_LUT4 add_5139_4_lut (.I0(GND_net), .I1(n17233[1]), .I2(n250), .I3(n38474), 
            .O(n16869[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_4 (.CI(n38474), .I0(n17233[1]), .I1(n250), .CO(n38475));
    SB_LUT4 add_5152_4_lut (.I0(GND_net), .I1(n17401[1]), .I2(n250_adj_4996), 
            .I3(n38717), .O(n17064[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5139_3_lut (.I0(GND_net), .I1(n17233[0]), .I2(n177), .I3(n38473), 
            .O(n16869[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5139_3 (.CI(n38473), .I0(n17233[0]), .I1(n177), .CO(n38474));
    SB_LUT4 add_5139_2_lut (.I0(GND_net), .I1(n35_adj_4997), .I2(n104), 
            .I3(GND_net), .O(n16869[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5139_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19998_2_lut (.I0(n28[18]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19998_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5152_4 (.CI(n38717), .I0(n17401[1]), .I1(n250_adj_4996), 
            .CO(n38718));
    SB_CARRY add_5139_2 (.CI(GND_net), .I0(n35_adj_4997), .I1(n104), .CO(n38473));
    SB_LUT4 i23792_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n18664[0]));   // verilog/motorControl.v(34[16:22])
    defparam i23792_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_5152_3_lut (.I0(GND_net), .I1(n17401[0]), .I2(n177_adj_4999), 
            .I3(n38716), .O(n17064[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_3 (.CI(n38716), .I0(n17401[0]), .I1(n177_adj_4999), 
            .CO(n38717));
    SB_LUT4 add_5152_2_lut (.I0(GND_net), .I1(n35_adj_5000), .I2(n104_adj_5001), 
            .I3(GND_net), .O(n17064[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5164_13_lut (.I0(GND_net), .I1(n17545[10]), .I2(n910), 
            .I3(n38472), .O(n17233[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_2 (.CI(GND_net), .I0(n35_adj_5000), .I1(n104_adj_5001), 
            .CO(n38716));
    SB_LUT4 add_5272_7_lut (.I0(GND_net), .I1(n43796), .I2(n490), .I3(n38715), 
            .O(n18465[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5164_12_lut (.I0(GND_net), .I1(n17545[9]), .I2(n837), 
            .I3(n38471), .O(n17233[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5272_6_lut (.I0(GND_net), .I1(n18549[3]), .I2(n417), .I3(n38714), 
            .O(n18465[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_6 (.CI(n38714), .I0(n18549[3]), .I1(n417), .CO(n38715));
    SB_LUT4 add_5272_5_lut (.I0(GND_net), .I1(n18549[2]), .I2(n344), .I3(n38713), 
            .O(n18465[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_5002));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5272_5 (.CI(n38713), .I0(n18549[2]), .I1(n344), .CO(n38714));
    SB_LUT4 add_5272_4_lut (.I0(GND_net), .I1(n18549[1]), .I2(n271_adj_5003), 
            .I3(n38712), .O(n18465[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_4 (.CI(n38712), .I0(n18549[1]), .I1(n271_adj_5003), 
            .CO(n38713));
    SB_CARRY add_5164_12 (.CI(n38471), .I0(n17545[9]), .I1(n837), .CO(n38472));
    SB_LUT4 add_5272_3_lut (.I0(GND_net), .I1(n18549[0]), .I2(n198_adj_5004), 
            .I3(n38711), .O(n18465[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5164_11_lut (.I0(GND_net), .I1(n17545[8]), .I2(n764), 
            .I3(n38470), .O(n17233[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n37710), .I0(GND_net), .I1(n1[7]), 
            .CO(n37711));
    SB_CARRY add_5164_11 (.CI(n38470), .I0(n17545[8]), .I1(n764), .CO(n38471));
    SB_LUT4 add_5164_10_lut (.I0(GND_net), .I1(n17545[7]), .I2(n691), 
            .I3(n38469), .O(n17233[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_10 (.CI(n38469), .I0(n17545[7]), .I1(n691), .CO(n38470));
    SB_CARRY add_5272_3 (.CI(n38711), .I0(n18549[0]), .I1(n198_adj_5004), 
            .CO(n38712));
    SB_LUT4 add_5164_9_lut (.I0(GND_net), .I1(n17545[6]), .I2(n618), .I3(n38468), 
            .O(n17233[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n37709), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n37709), .I0(GND_net), .I1(n1[6]), 
            .CO(n37710));
    SB_CARRY add_5164_9 (.CI(n38468), .I0(n17545[6]), .I1(n618), .CO(n38469));
    SB_LUT4 add_5272_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n18465[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5272_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5164_8_lut (.I0(GND_net), .I1(n17545[5]), .I2(n545), .I3(n38467), 
            .O(n17233[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5272_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n38711));
    SB_LUT4 add_5176_13_lut (.I0(GND_net), .I1(n17688[10]), .I2(n910_adj_5006), 
            .I3(n38710), .O(n17401[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5176_12_lut (.I0(GND_net), .I1(n17688[9]), .I2(n837_adj_5007), 
            .I3(n38709), .O(n17401[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_8 (.CI(n38467), .I0(n17545[5]), .I1(n545), .CO(n38468));
    SB_CARRY add_5176_12 (.CI(n38709), .I0(n17688[9]), .I1(n837_adj_5007), 
            .CO(n38710));
    SB_LUT4 add_5164_7_lut (.I0(GND_net), .I1(n17545[4]), .I2(n472), .I3(n38466), 
            .O(n17233[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_7 (.CI(n38466), .I0(n17545[4]), .I1(n472), .CO(n38467));
    SB_LUT4 add_5164_6_lut (.I0(GND_net), .I1(n17545[3]), .I2(n399), .I3(n38465), 
            .O(n17233[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n37708), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_6 (.CI(n38465), .I0(n17545[3]), .I1(n399), .CO(n38466));
    SB_LUT4 add_5164_5_lut (.I0(GND_net), .I1(n17545[2]), .I2(n326), .I3(n38464), 
            .O(n17233[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n37708), .I0(GND_net), .I1(n1[5]), 
            .CO(n37709));
    SB_CARRY add_5164_5 (.CI(n38464), .I0(n17545[2]), .I1(n326), .CO(n38465));
    SB_LUT4 add_5164_4_lut (.I0(GND_net), .I1(n17545[1]), .I2(n253), .I3(n38463), 
            .O(n17233[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_4 (.CI(n38463), .I0(n17545[1]), .I1(n253), .CO(n38464));
    SB_LUT4 add_5164_3_lut (.I0(GND_net), .I1(n17545[0]), .I2(n180), .I3(n38462), 
            .O(n17233[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_3 (.CI(n38462), .I0(n17545[0]), .I1(n180), .CO(n38463));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n37707), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5164_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n17233[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5176_11_lut (.I0(GND_net), .I1(n17688[8]), .I2(n764_adj_5010), 
            .I3(n38708), .O(n17401[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_11 (.CI(n38708), .I0(n17688[8]), .I1(n764_adj_5010), 
            .CO(n38709));
    SB_LUT4 add_5176_10_lut (.I0(GND_net), .I1(n17688[7]), .I2(n691_adj_5011), 
            .I3(n38707), .O(n17401[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n38462));
    SB_CARRY add_5176_10 (.CI(n38707), .I0(n17688[7]), .I1(n691_adj_5011), 
            .CO(n38708));
    SB_LUT4 add_5278_7_lut (.I0(GND_net), .I1(n44030), .I2(n490_adj_5012), 
            .I3(n38461), .O(n18513[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5176_9_lut (.I0(GND_net), .I1(n17688[6]), .I2(n618_adj_5013), 
            .I3(n38706), .O(n17401[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5278_6_lut (.I0(GND_net), .I1(n18584[3]), .I2(n417_adj_5014), 
            .I3(n38460), .O(n18513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_9 (.CI(n38706), .I0(n17688[6]), .I1(n618_adj_5013), 
            .CO(n38707));
    SB_LUT4 add_5176_8_lut (.I0(GND_net), .I1(n17688[5]), .I2(n545_adj_5015), 
            .I3(n38705), .O(n17401[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_8 (.CI(n38705), .I0(n17688[5]), .I1(n545_adj_5015), 
            .CO(n38706));
    SB_LUT4 add_5176_7_lut (.I0(GND_net), .I1(n17688[4]), .I2(n472_adj_5016), 
            .I3(n38704), .O(n17401[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_7 (.CI(n38704), .I0(n17688[4]), .I1(n472_adj_5016), 
            .CO(n38705));
    SB_LUT4 add_5176_6_lut (.I0(GND_net), .I1(n17688[3]), .I2(n399_adj_5017), 
            .I3(n38703), .O(n17401[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_6 (.CI(n38703), .I0(n17688[3]), .I1(n399_adj_5017), 
            .CO(n38704));
    SB_LUT4 add_5176_5_lut (.I0(GND_net), .I1(n17688[2]), .I2(n326_adj_5018), 
            .I3(n38702), .O(n17401[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_5 (.CI(n38702), .I0(n17688[2]), .I1(n326_adj_5018), 
            .CO(n38703));
    SB_LUT4 add_5176_4_lut (.I0(GND_net), .I1(n17688[1]), .I2(n253_adj_5019), 
            .I3(n38701), .O(n17401[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_4 (.CI(n38701), .I0(n17688[1]), .I1(n253_adj_5019), 
            .CO(n38702));
    SB_LUT4 add_5176_3_lut (.I0(GND_net), .I1(n17688[0]), .I2(n180_adj_5020), 
            .I3(n38700), .O(n17401[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5176_3 (.CI(n38700), .I0(n17688[0]), .I1(n180_adj_5020), 
            .CO(n38701));
    SB_LUT4 add_5176_2_lut (.I0(GND_net), .I1(n38_adj_5021), .I2(n107_adj_5022), 
            .I3(GND_net), .O(n17401[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5176_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23794_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n37292));   // verilog/motorControl.v(34[16:22])
    defparam i23794_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n37707), .I0(GND_net), .I1(n1[4]), 
            .CO(n37708));
    SB_CARRY add_5176_2 (.CI(GND_net), .I0(n38_adj_5021), .I1(n107_adj_5022), 
            .CO(n38700));
    SB_LUT4 add_5198_12_lut (.I0(GND_net), .I1(n17929[9]), .I2(n840_adj_5023), 
            .I3(n38699), .O(n17688[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n37706), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_6 (.CI(n38460), .I0(n18584[3]), .I1(n417_adj_5014), 
            .CO(n38461));
    SB_CARRY unary_minus_16_add_3_5 (.CI(n37706), .I0(GND_net), .I1(n1[3]), 
            .CO(n37707));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n37705), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5198_11_lut (.I0(GND_net), .I1(n17929[8]), .I2(n767_adj_5026), 
            .I3(n38698), .O(n17688[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5278_5_lut (.I0(GND_net), .I1(n18584[2]), .I2(n344_adj_5027), 
            .I3(n38459), .O(n18513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_5028));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5198_11 (.CI(n38698), .I0(n17929[8]), .I1(n767_adj_5026), 
            .CO(n38699));
    SB_CARRY unary_minus_16_add_3_4 (.CI(n37705), .I0(GND_net), .I1(n1[2]), 
            .CO(n37706));
    SB_LUT4 add_5198_10_lut (.I0(GND_net), .I1(n17929[7]), .I2(n694_adj_5029), 
            .I3(n38697), .O(n17688[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n37704), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_10 (.CI(n38697), .I0(n17929[7]), .I1(n694_adj_5029), 
            .CO(n38698));
    SB_LUT4 add_5198_9_lut (.I0(GND_net), .I1(n17929[6]), .I2(n621_adj_5031), 
            .I3(n38696), .O(n17688[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n37704), .I0(GND_net), .I1(n1[1]), 
            .CO(n37705));
    SB_CARRY add_5198_9 (.CI(n38696), .I0(n17929[6]), .I1(n621_adj_5031), 
            .CO(n38697));
    SB_LUT4 add_5198_8_lut (.I0(GND_net), .I1(n17929[5]), .I2(n548_adj_5032), 
            .I3(n38695), .O(n17688[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_8 (.CI(n38695), .I0(n17929[5]), .I1(n548_adj_5032), 
            .CO(n38696));
    SB_LUT4 add_5198_7_lut (.I0(GND_net), .I1(n17929[4]), .I2(n475_adj_5033), 
            .I3(n38694), .O(n17688[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_7 (.CI(n38694), .I0(n17929[4]), .I1(n475_adj_5033), 
            .CO(n38695));
    SB_LUT4 add_5198_6_lut (.I0(GND_net), .I1(n17929[3]), .I2(n402_adj_5034), 
            .I3(n38693), .O(n17688[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_6 (.CI(n38693), .I0(n17929[3]), .I1(n402_adj_5034), 
            .CO(n38694));
    SB_LUT4 add_5198_5_lut (.I0(GND_net), .I1(n17929[2]), .I2(n329_adj_5035), 
            .I3(n38692), .O(n17688[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_5 (.CI(n38459), .I0(n18584[2]), .I1(n344_adj_5027), 
            .CO(n38460));
    SB_CARRY add_5198_5 (.CI(n38692), .I0(n17929[2]), .I1(n329_adj_5035), 
            .CO(n38693));
    SB_LUT4 add_5198_4_lut (.I0(GND_net), .I1(n17929[1]), .I2(n256_adj_5036), 
            .I3(n38691), .O(n17688[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_4 (.CI(n38691), .I0(n17929[1]), .I1(n256_adj_5036), 
            .CO(n38692));
    SB_LUT4 add_5198_3_lut (.I0(GND_net), .I1(n17929[0]), .I2(n183_adj_5037), 
            .I3(n38690), .O(n17688[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_3 (.CI(n38690), .I0(n17929[0]), .I1(n183_adj_5037), 
            .CO(n38691));
    SB_LUT4 add_5198_2_lut (.I0(GND_net), .I1(n41_adj_5038), .I2(n110_adj_5039), 
            .I3(GND_net), .O(n17688[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5198_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5198_2 (.CI(GND_net), .I0(n41_adj_5038), .I1(n110_adj_5039), 
            .CO(n38690));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I1(n10590[21]), .I2(GND_net), .I3(n38689), .O(n10083[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n10590[20]), .I2(GND_net), 
            .I3(n38688), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n38688), .I0(n10590[20]), .I1(GND_net), 
            .CO(n38689));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n10590[19]), .I2(GND_net), 
            .I3(n38687), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n37704));
    SB_CARRY mult_11_add_1225_22 (.CI(n38687), .I0(n10590[19]), .I1(GND_net), 
            .CO(n38688));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n10590[18]), .I2(GND_net), 
            .I3(n38686), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5132[23]), 
            .I3(n37703), .O(\PID_CONTROLLER.integral_23__N_3723 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_5132[22]), .I3(n37702), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n37702), .I0(GND_net), .I1(n1_adj_5132[22]), 
            .CO(n37703));
    SB_CARRY mult_11_add_1225_21 (.CI(n38686), .I0(n10590[18]), .I1(GND_net), 
            .CO(n38687));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n10590[17]), .I2(GND_net), 
            .I3(n38685), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n38685), .I0(n10590[17]), .I1(GND_net), 
            .CO(n38686));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n10590[16]), .I2(GND_net), 
            .I3(n38684), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n38684), .I0(n10590[16]), .I1(GND_net), 
            .CO(n38685));
    SB_LUT4 add_5278_4_lut (.I0(GND_net), .I1(n18584[1]), .I2(n271_adj_5043), 
            .I3(n38458), .O(n18513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n10590[15]), .I2(GND_net), 
            .I3(n38683), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_4 (.CI(n38458), .I0(n18584[1]), .I1(n271_adj_5043), 
            .CO(n38459));
    SB_CARRY mult_11_add_1225_18 (.CI(n38683), .I0(n10590[15]), .I1(GND_net), 
            .CO(n38684));
    SB_LUT4 add_5278_3_lut (.I0(GND_net), .I1(n18584[0]), .I2(n198_adj_5044), 
            .I3(n38457), .O(n18513[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n10590[14]), .I2(GND_net), 
            .I3(n38682), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_3 (.CI(n38457), .I0(n18584[0]), .I1(n198_adj_5044), 
            .CO(n38458));
    SB_CARRY mult_11_add_1225_17 (.CI(n38682), .I0(n10590[14]), .I1(GND_net), 
            .CO(n38683));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n10590[13]), .I2(n1096_adj_5045), 
            .I3(n38681), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n38681), .I0(n10590[13]), .I1(n1096_adj_5045), 
            .CO(n38682));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n10590[12]), .I2(n1023_adj_5046), 
            .I3(n38680), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n38680), .I0(n10590[12]), .I1(n1023_adj_5046), 
            .CO(n38681));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n10590[11]), .I2(n950_adj_5047), 
            .I3(n38679), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5278_2_lut (.I0(GND_net), .I1(n56_adj_5048), .I2(n125_adj_5049), 
            .I3(GND_net), .O(n18513[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5278_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n38679), .I0(n10590[11]), .I1(n950_adj_5047), 
            .CO(n38680));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n10590[10]), .I2(n877_adj_5050), 
            .I3(n38678), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n38678), .I0(n10590[10]), .I1(n877_adj_5050), 
            .CO(n38679));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n10590[9]), .I2(n804_adj_5051), 
            .I3(n38677), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n38677), .I0(n10590[9]), .I1(n804_adj_5051), 
            .CO(n38678));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n10590[8]), .I2(n731_adj_5052), 
            .I3(n38676), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n38676), .I0(n10590[8]), .I1(n731_adj_5052), 
            .CO(n38677));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n10590[7]), .I2(n658_adj_5053), 
            .I3(n38675), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n38675), .I0(n10590[7]), .I1(n658_adj_5053), 
            .CO(n38676));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n10590[6]), .I2(n585_adj_5054), 
            .I3(n38674), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n38674), .I0(n10590[6]), .I1(n585_adj_5054), 
            .CO(n38675));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n10590[5]), .I2(n512_adj_5055), 
            .I3(n38673), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n38673), .I0(n10590[5]), .I1(n512_adj_5055), 
            .CO(n38674));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n10590[4]), .I2(n439_adj_5056), 
            .I3(n38672), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n38672), .I0(n10590[4]), .I1(n439_adj_5056), 
            .CO(n38673));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n10590[3]), .I2(n366_adj_5057), 
            .I3(n38671), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n38671), .I0(n10590[3]), .I1(n366_adj_5057), 
            .CO(n38672));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n10590[2]), .I2(n293_adj_5058), 
            .I3(n38670), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n38670), .I0(n10590[2]), .I1(n293_adj_5058), 
            .CO(n38671));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n10590[1]), .I2(n220_adj_5059), 
            .I3(n38669), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n38669), .I0(n10590[1]), .I1(n220_adj_5059), 
            .CO(n38670));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n10590[0]), .I2(n147_adj_5060), 
            .I3(n38668), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n38668), .I0(n10590[0]), .I1(n147_adj_5060), 
            .CO(n38669));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_5061), .I2(n74_adj_5062), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5278_2 (.CI(GND_net), .I0(n56_adj_5048), .I1(n125_adj_5049), 
            .CO(n38457));
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_5061), .I1(n74_adj_5062), 
            .CO(n38668));
    SB_LUT4 add_4823_23_lut (.I0(GND_net), .I1(n11605[20]), .I2(GND_net), 
            .I3(n38667), .O(n10590[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4823_22_lut (.I0(GND_net), .I1(n11605[19]), .I2(GND_net), 
            .I3(n38666), .O(n10590[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_22 (.CI(n38666), .I0(n11605[19]), .I1(GND_net), 
            .CO(n38667));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_5132[21]), .I3(n37701), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4823_21_lut (.I0(GND_net), .I1(n11605[18]), .I2(GND_net), 
            .I3(n38665), .O(n10590[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_21 (.CI(n38665), .I0(n11605[18]), .I1(GND_net), 
            .CO(n38666));
    SB_LUT4 add_4823_20_lut (.I0(GND_net), .I1(n11605[17]), .I2(GND_net), 
            .I3(n38664), .O(n10590[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_20 (.CI(n38664), .I0(n11605[17]), .I1(GND_net), 
            .CO(n38665));
    SB_LUT4 add_4823_19_lut (.I0(GND_net), .I1(n11605[16]), .I2(GND_net), 
            .I3(n38663), .O(n10590[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_19 (.CI(n38663), .I0(n11605[16]), .I1(GND_net), 
            .CO(n38664));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n37701), .I0(GND_net), .I1(n1_adj_5132[21]), 
            .CO(n37702));
    SB_LUT4 add_4823_18_lut (.I0(GND_net), .I1(n11605[15]), .I2(GND_net), 
            .I3(n38662), .O(n10590[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_18 (.CI(n38662), .I0(n11605[15]), .I1(GND_net), 
            .CO(n38663));
    SB_LUT4 add_4823_17_lut (.I0(GND_net), .I1(n11605[14]), .I2(GND_net), 
            .I3(n38661), .O(n10590[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_17 (.CI(n38661), .I0(n11605[14]), .I1(GND_net), 
            .CO(n38662));
    SB_LUT4 add_4823_16_lut (.I0(GND_net), .I1(n11605[13]), .I2(n1099_adj_5064), 
            .I3(n38660), .O(n10590[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_16 (.CI(n38660), .I0(n11605[13]), .I1(n1099_adj_5064), 
            .CO(n38661));
    SB_LUT4 add_4823_15_lut (.I0(GND_net), .I1(n11605[12]), .I2(n1026_adj_5065), 
            .I3(n38659), .O(n10590[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_15 (.CI(n38659), .I0(n11605[12]), .I1(n1026_adj_5065), 
            .CO(n38660));
    SB_LUT4 add_4823_14_lut (.I0(GND_net), .I1(n11605[11]), .I2(n953_adj_5066), 
            .I3(n38658), .O(n10590[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_14 (.CI(n38658), .I0(n11605[11]), .I1(n953_adj_5066), 
            .CO(n38659));
    SB_LUT4 add_4823_13_lut (.I0(GND_net), .I1(n11605[10]), .I2(n880_adj_5067), 
            .I3(n38657), .O(n10590[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_13 (.CI(n38657), .I0(n11605[10]), .I1(n880_adj_5067), 
            .CO(n38658));
    SB_LUT4 add_4823_12_lut (.I0(GND_net), .I1(n11605[9]), .I2(n807_adj_5068), 
            .I3(n38656), .O(n10590[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_12 (.CI(n38656), .I0(n11605[9]), .I1(n807_adj_5068), 
            .CO(n38657));
    SB_LUT4 add_4823_11_lut (.I0(GND_net), .I1(n11605[8]), .I2(n734_adj_5069), 
            .I3(n38655), .O(n10590[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_11 (.CI(n38655), .I0(n11605[8]), .I1(n734_adj_5069), 
            .CO(n38656));
    SB_LUT4 add_4823_10_lut (.I0(GND_net), .I1(n11605[7]), .I2(n661_adj_5070), 
            .I3(n38654), .O(n10590[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_10 (.CI(n38654), .I0(n11605[7]), .I1(n661_adj_5070), 
            .CO(n38655));
    SB_LUT4 add_4823_9_lut (.I0(GND_net), .I1(n11605[6]), .I2(n588_adj_5071), 
            .I3(n38653), .O(n10590[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_9 (.CI(n38653), .I0(n11605[6]), .I1(n588_adj_5071), 
            .CO(n38654));
    SB_LUT4 add_4823_8_lut (.I0(GND_net), .I1(n11605[5]), .I2(n515_adj_5072), 
            .I3(n38652), .O(n10590[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_8 (.CI(n38652), .I0(n11605[5]), .I1(n515_adj_5072), 
            .CO(n38653));
    SB_LUT4 add_4823_7_lut (.I0(GND_net), .I1(n11605[4]), .I2(n442_adj_5073), 
            .I3(n38651), .O(n10590[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_7 (.CI(n38651), .I0(n11605[4]), .I1(n442_adj_5073), 
            .CO(n38652));
    SB_LUT4 add_4823_6_lut (.I0(GND_net), .I1(n11605[3]), .I2(n369_adj_5074), 
            .I3(n38650), .O(n10590[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_6 (.CI(n38650), .I0(n11605[3]), .I1(n369_adj_5074), 
            .CO(n38651));
    SB_LUT4 add_4823_5_lut (.I0(GND_net), .I1(n11605[2]), .I2(n296_adj_5075), 
            .I3(n38649), .O(n10590[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_5 (.CI(n38649), .I0(n11605[2]), .I1(n296_adj_5075), 
            .CO(n38650));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_5132[20]), .I3(n37700), .O(n41_adj_4905)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4823_4_lut (.I0(GND_net), .I1(n11605[1]), .I2(n223_adj_5077), 
            .I3(n38648), .O(n10590[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_4 (.CI(n38648), .I0(n11605[1]), .I1(n223_adj_5077), 
            .CO(n38649));
    SB_LUT4 add_4823_3_lut (.I0(GND_net), .I1(n11605[0]), .I2(n150_adj_5078), 
            .I3(n38647), .O(n10590[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_3 (.CI(n38647), .I0(n11605[0]), .I1(n150_adj_5078), 
            .CO(n38648));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n37700), .I0(GND_net), .I1(n1_adj_5132[20]), 
            .CO(n37701));
    SB_LUT4 add_4823_2_lut (.I0(GND_net), .I1(n8_adj_5079), .I2(n77_adj_5080), 
            .I3(GND_net), .O(n10590[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4823_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4823_2 (.CI(GND_net), .I0(n8_adj_5079), .I1(n77_adj_5080), 
            .CO(n38647));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_5132[19]), .I3(n37699), .O(n39_adj_4903)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4867_22_lut (.I0(GND_net), .I1(n12529[19]), .I2(GND_net), 
            .I3(n38646), .O(n11605[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4867_21_lut (.I0(GND_net), .I1(n12529[18]), .I2(GND_net), 
            .I3(n38645), .O(n11605[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_21 (.CI(n38645), .I0(n12529[18]), .I1(GND_net), 
            .CO(n38646));
    SB_CARRY unary_minus_5_add_3_21 (.CI(n37699), .I0(GND_net), .I1(n1_adj_5132[19]), 
            .CO(n37700));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_5132[18]), .I3(n37698), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n37698), .I0(GND_net), .I1(n1_adj_5132[18]), 
            .CO(n37699));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_5132[17]), .I3(n37697), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n37697), .I0(GND_net), .I1(n1_adj_5132[17]), 
            .CO(n37698));
    SB_LUT4 add_4867_20_lut (.I0(GND_net), .I1(n12529[17]), .I2(GND_net), 
            .I3(n38644), .O(n11605[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_20 (.CI(n38644), .I0(n12529[17]), .I1(GND_net), 
            .CO(n38645));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_5132[16]), .I3(n37696), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4867_19_lut (.I0(GND_net), .I1(n12529[16]), .I2(GND_net), 
            .I3(n38643), .O(n11605[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_19 (.CI(n38643), .I0(n12529[16]), .I1(GND_net), 
            .CO(n38644));
    SB_LUT4 add_4867_18_lut (.I0(GND_net), .I1(n12529[15]), .I2(GND_net), 
            .I3(n38642), .O(n11605[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_18 (.CI(n38642), .I0(n12529[15]), .I1(GND_net), 
            .CO(n38643));
    SB_LUT4 add_4867_17_lut (.I0(GND_net), .I1(n12529[14]), .I2(GND_net), 
            .I3(n38641), .O(n11605[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_17 (.CI(n38641), .I0(n12529[14]), .I1(GND_net), 
            .CO(n38642));
    SB_CARRY unary_minus_5_add_3_18 (.CI(n37696), .I0(GND_net), .I1(n1_adj_5132[16]), 
            .CO(n37697));
    SB_LUT4 add_4867_16_lut (.I0(GND_net), .I1(n12529[13]), .I2(n1102_adj_5085), 
            .I3(n38640), .O(n11605[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_5132[15]), .I3(n37695), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4867_16 (.CI(n38640), .I0(n12529[13]), .I1(n1102_adj_5085), 
            .CO(n38641));
    SB_LUT4 add_4867_15_lut (.I0(GND_net), .I1(n12529[12]), .I2(n1029_adj_5087), 
            .I3(n38639), .O(n11605[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_15 (.CI(n38639), .I0(n12529[12]), .I1(n1029_adj_5087), 
            .CO(n38640));
    SB_LUT4 add_4867_14_lut (.I0(GND_net), .I1(n12529[11]), .I2(n956_adj_5088), 
            .I3(n38638), .O(n11605[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_14 (.CI(n38638), .I0(n12529[11]), .I1(n956_adj_5088), 
            .CO(n38639));
    SB_LUT4 add_4867_13_lut (.I0(GND_net), .I1(n12529[10]), .I2(n883_adj_5089), 
            .I3(n38637), .O(n11605[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_13 (.CI(n38637), .I0(n12529[10]), .I1(n883_adj_5089), 
            .CO(n38638));
    SB_LUT4 add_4867_12_lut (.I0(GND_net), .I1(n12529[9]), .I2(n810_adj_5090), 
            .I3(n38636), .O(n11605[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_12 (.CI(n38636), .I0(n12529[9]), .I1(n810_adj_5090), 
            .CO(n38637));
    SB_LUT4 add_4867_11_lut (.I0(GND_net), .I1(n12529[8]), .I2(n737_adj_5091), 
            .I3(n38635), .O(n11605[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_11 (.CI(n38635), .I0(n12529[8]), .I1(n737_adj_5091), 
            .CO(n38636));
    SB_CARRY unary_minus_5_add_3_17 (.CI(n37695), .I0(GND_net), .I1(n1_adj_5132[15]), 
            .CO(n37696));
    SB_LUT4 add_4867_10_lut (.I0(GND_net), .I1(n12529[7]), .I2(n664_adj_5092), 
            .I3(n38634), .O(n11605[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_10 (.CI(n38634), .I0(n12529[7]), .I1(n664_adj_5092), 
            .CO(n38635));
    SB_LUT4 add_4867_9_lut (.I0(GND_net), .I1(n12529[6]), .I2(n591_adj_5093), 
            .I3(n38633), .O(n11605[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_9 (.CI(n38633), .I0(n12529[6]), .I1(n591_adj_5093), 
            .CO(n38634));
    SB_LUT4 add_4867_8_lut (.I0(GND_net), .I1(n12529[5]), .I2(n518_adj_5094), 
            .I3(n38632), .O(n11605[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_8 (.CI(n38632), .I0(n12529[5]), .I1(n518_adj_5094), 
            .CO(n38633));
    SB_LUT4 add_4867_7_lut (.I0(GND_net), .I1(n12529[4]), .I2(n445_adj_5095), 
            .I3(n38631), .O(n11605[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_7 (.CI(n38631), .I0(n12529[4]), .I1(n445_adj_5095), 
            .CO(n38632));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_5132[14]), .I3(n37694), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4867_6_lut (.I0(GND_net), .I1(n12529[3]), .I2(n372_adj_5097), 
            .I3(n38630), .O(n11605[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_6 (.CI(n38630), .I0(n12529[3]), .I1(n372_adj_5097), 
            .CO(n38631));
    SB_LUT4 add_958_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n4236[23]), .I3(n37611), .O(\PID_CONTROLLER.integral_23__N_3672 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n37694), .I0(GND_net), .I1(n1_adj_5132[14]), 
            .CO(n37695));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_5132[13]), .I3(n37693), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_958_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n4236[22]), .I3(n37610), .O(\PID_CONTROLLER.integral_23__N_3672 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n37693), .I0(GND_net), .I1(n1_adj_5132[13]), 
            .CO(n37694));
    SB_CARRY add_958_24 (.CI(n37610), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n4236[22]), .CO(n37611));
    SB_LUT4 add_4867_5_lut (.I0(GND_net), .I1(n12529[2]), .I2(n299_adj_5099), 
            .I3(n38629), .O(n11605[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_5 (.CI(n38629), .I0(n12529[2]), .I1(n299_adj_5099), 
            .CO(n38630));
    SB_LUT4 add_4867_4_lut (.I0(GND_net), .I1(n12529[1]), .I2(n226_adj_5100), 
            .I3(n38628), .O(n11605[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_4 (.CI(n38628), .I0(n12529[1]), .I1(n226_adj_5100), 
            .CO(n38629));
    SB_LUT4 add_4867_3_lut (.I0(GND_net), .I1(n12529[0]), .I2(n153_adj_5101), 
            .I3(n38627), .O(n11605[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_3 (.CI(n38627), .I0(n12529[0]), .I1(n153_adj_5101), 
            .CO(n38628));
    SB_LUT4 add_4867_2_lut (.I0(GND_net), .I1(n11_adj_5102), .I2(n80_adj_5103), 
            .I3(GND_net), .O(n11605[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4867_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4867_2 (.CI(GND_net), .I0(n11_adj_5102), .I1(n80_adj_5103), 
            .CO(n38627));
    SB_LUT4 add_4908_21_lut (.I0(GND_net), .I1(n13369[18]), .I2(GND_net), 
            .I3(n38626), .O(n12529[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4908_20_lut (.I0(GND_net), .I1(n13369[17]), .I2(GND_net), 
            .I3(n38625), .O(n12529[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_20 (.CI(n38625), .I0(n13369[17]), .I1(GND_net), 
            .CO(n38626));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_5132[12]), .I3(n37692), .O(n25_adj_4794)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_958_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n4236[21]), .I3(n37609), .O(\PID_CONTROLLER.integral_23__N_3672 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n37692), .I0(GND_net), .I1(n1_adj_5132[12]), 
            .CO(n37693));
    SB_CARRY add_958_23 (.CI(n37609), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n4236[21]), .CO(n37610));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_5132[11]), .I3(n37691), .O(n23_adj_4795)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_958_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n4236[20]), .I3(n37608), .O(\PID_CONTROLLER.integral_23__N_3672 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n37691), .I0(GND_net), .I1(n1_adj_5132[11]), 
            .CO(n37692));
    SB_LUT4 add_4908_19_lut (.I0(GND_net), .I1(n13369[16]), .I2(GND_net), 
            .I3(n38624), .O(n12529[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_19 (.CI(n38624), .I0(n13369[16]), .I1(GND_net), 
            .CO(n38625));
    SB_LUT4 add_4908_18_lut (.I0(GND_net), .I1(n13369[15]), .I2(GND_net), 
            .I3(n38623), .O(n12529[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_18 (.CI(n38623), .I0(n13369[15]), .I1(GND_net), 
            .CO(n38624));
    SB_LUT4 add_4908_17_lut (.I0(GND_net), .I1(n13369[14]), .I2(GND_net), 
            .I3(n38622), .O(n12529[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_17 (.CI(n38622), .I0(n13369[14]), .I1(GND_net), 
            .CO(n38623));
    SB_LUT4 add_4908_16_lut (.I0(GND_net), .I1(n13369[13]), .I2(n1105_adj_5106), 
            .I3(n38621), .O(n12529[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_16 (.CI(n38621), .I0(n13369[13]), .I1(n1105_adj_5106), 
            .CO(n38622));
    SB_LUT4 add_4908_15_lut (.I0(GND_net), .I1(n13369[12]), .I2(n1032_adj_5107), 
            .I3(n38620), .O(n12529[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_15 (.CI(n38620), .I0(n13369[12]), .I1(n1032_adj_5107), 
            .CO(n38621));
    SB_CARRY add_958_22 (.CI(n37608), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n4236[20]), .CO(n37609));
    SB_LUT4 add_4908_14_lut (.I0(GND_net), .I1(n13369[11]), .I2(n959_adj_5108), 
            .I3(n38619), .O(n12529[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_14 (.CI(n38619), .I0(n13369[11]), .I1(n959_adj_5108), 
            .CO(n38620));
    SB_LUT4 add_4908_13_lut (.I0(GND_net), .I1(n13369[10]), .I2(n886_adj_5109), 
            .I3(n38618), .O(n12529[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_13 (.CI(n38618), .I0(n13369[10]), .I1(n886_adj_5109), 
            .CO(n38619));
    SB_LUT4 add_4908_12_lut (.I0(GND_net), .I1(n13369[9]), .I2(n813_adj_5110), 
            .I3(n38617), .O(n12529[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_12 (.CI(n38617), .I0(n13369[9]), .I1(n813_adj_5110), 
            .CO(n38618));
    SB_LUT4 add_4908_11_lut (.I0(GND_net), .I1(n13369[8]), .I2(n740_adj_5111), 
            .I3(n38616), .O(n12529[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_11 (.CI(n38616), .I0(n13369[8]), .I1(n740_adj_5111), 
            .CO(n38617));
    SB_LUT4 add_4908_10_lut (.I0(GND_net), .I1(n13369[7]), .I2(n667_adj_5112), 
            .I3(n38615), .O(n12529[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n4236[19]), .I3(n37607), .O(\PID_CONTROLLER.integral_23__N_3672 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_10 (.CI(n38615), .I0(n13369[7]), .I1(n667_adj_5112), 
            .CO(n38616));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_5132[10]), .I3(n37690), .O(n21_adj_4772)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_958_21 (.CI(n37607), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n4236[19]), .CO(n37608));
    SB_LUT4 add_4908_9_lut (.I0(GND_net), .I1(n13369[6]), .I2(n594_adj_5114), 
            .I3(n38614), .O(n12529[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_9 (.CI(n38614), .I0(n13369[6]), .I1(n594_adj_5114), 
            .CO(n38615));
    SB_LUT4 add_4908_8_lut (.I0(GND_net), .I1(n13369[5]), .I2(n521_adj_5115), 
            .I3(n38613), .O(n12529[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_8 (.CI(n38613), .I0(n13369[5]), .I1(n521_adj_5115), 
            .CO(n38614));
    SB_LUT4 add_4908_7_lut (.I0(GND_net), .I1(n13369[4]), .I2(n448_adj_5116), 
            .I3(n38612), .O(n12529[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_7 (.CI(n38612), .I0(n13369[4]), .I1(n448_adj_5116), 
            .CO(n38613));
    SB_LUT4 add_4908_6_lut (.I0(GND_net), .I1(n13369[3]), .I2(n375_adj_5117), 
            .I3(n38611), .O(n12529[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_6 (.CI(n38611), .I0(n13369[3]), .I1(n375_adj_5117), 
            .CO(n38612));
    SB_LUT4 add_4908_5_lut (.I0(GND_net), .I1(n13369[2]), .I2(n302_adj_5118), 
            .I3(n38610), .O(n12529[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_5 (.CI(n38610), .I0(n13369[2]), .I1(n302_adj_5118), 
            .CO(n38611));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n37690), .I0(GND_net), .I1(n1_adj_5132[10]), 
            .CO(n37691));
    SB_LUT4 add_4908_4_lut (.I0(GND_net), .I1(n13369[1]), .I2(n229_adj_5028), 
            .I3(n38609), .O(n12529[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_4 (.CI(n38609), .I0(n13369[1]), .I1(n229_adj_5028), 
            .CO(n38610));
    SB_LUT4 add_4908_3_lut (.I0(GND_net), .I1(n13369[0]), .I2(n156_adj_5002), 
            .I3(n38608), .O(n12529[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4236[18]), .I3(n37606), .O(\PID_CONTROLLER.integral_23__N_3672 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4908_3 (.CI(n38608), .I0(n13369[0]), .I1(n156_adj_5002), 
            .CO(n38609));
    SB_LUT4 add_4908_2_lut (.I0(GND_net), .I1(n14_adj_4991), .I2(n83_adj_4989), 
            .I3(GND_net), .O(n12529[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4908_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_5132[9]), .I3(n37689), .O(n19_adj_4773)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4908_2 (.CI(GND_net), .I0(n14_adj_4991), .I1(n83_adj_4989), 
            .CO(n38608));
    SB_LUT4 add_5218_11_lut (.I0(GND_net), .I1(n18128[8]), .I2(n770_adj_4968), 
            .I3(n38607), .O(n17929[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n37689), .I0(GND_net), .I1(n1_adj_5132[9]), 
            .CO(n37690));
    SB_LUT4 add_5218_10_lut (.I0(GND_net), .I1(n18128[7]), .I2(n697_adj_4954), 
            .I3(n38606), .O(n17929[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_5118));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5218_10 (.CI(n38606), .I0(n18128[7]), .I1(n697_adj_4954), 
            .CO(n38607));
    SB_LUT4 add_5218_9_lut (.I0(GND_net), .I1(n18128[6]), .I2(n624_adj_4953), 
            .I3(n38605), .O(n17929[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_20 (.CI(n37606), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n4236[18]), .CO(n37607));
    SB_CARRY add_5218_9 (.CI(n38605), .I0(n18128[6]), .I1(n624_adj_4953), 
            .CO(n38606));
    SB_LUT4 add_5218_8_lut (.I0(GND_net), .I1(n18128[5]), .I2(n551_adj_4951), 
            .I3(n38604), .O(n17929[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_8 (.CI(n38604), .I0(n18128[5]), .I1(n551_adj_4951), 
            .CO(n38605));
    SB_LUT4 add_5218_7_lut (.I0(GND_net), .I1(n18128[4]), .I2(n478_adj_4950), 
            .I3(n38603), .O(n17929[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_7 (.CI(n38603), .I0(n18128[4]), .I1(n478_adj_4950), 
            .CO(n38604));
    SB_LUT4 add_5218_6_lut (.I0(GND_net), .I1(n18128[3]), .I2(n405_adj_4947), 
            .I3(n38602), .O(n17929[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_6 (.CI(n38602), .I0(n18128[3]), .I1(n405_adj_4947), 
            .CO(n38603));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_5132[8]), .I3(n37688), .O(n17_adj_4774)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5218_5_lut (.I0(GND_net), .I1(n18128[2]), .I2(n332_adj_4937), 
            .I3(n38601), .O(n17929[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_5 (.CI(n38601), .I0(n18128[2]), .I1(n332_adj_4937), 
            .CO(n38602));
    SB_LUT4 add_5218_4_lut (.I0(GND_net), .I1(n18128[1]), .I2(n259_adj_4932), 
            .I3(n38600), .O(n17929[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_4 (.CI(n38600), .I0(n18128[1]), .I1(n259_adj_4932), 
            .CO(n38601));
    SB_LUT4 add_5218_3_lut (.I0(GND_net), .I1(n18128[0]), .I2(n186_adj_4931), 
            .I3(n38599), .O(n17929[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n37688), .I0(GND_net), .I1(n1_adj_5132[8]), 
            .CO(n37689));
    SB_CARRY add_5218_3 (.CI(n38599), .I0(n18128[0]), .I1(n186_adj_4931), 
            .CO(n38600));
    SB_LUT4 add_5218_2_lut (.I0(GND_net), .I1(n44_adj_4915), .I2(n113_adj_4914), 
            .I3(GND_net), .O(n17929[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_2 (.CI(GND_net), .I0(n44_adj_4915), .I1(n113_adj_4914), 
            .CO(n38599));
    SB_LUT4 add_4947_20_lut (.I0(GND_net), .I1(n14129[17]), .I2(GND_net), 
            .I3(n38598), .O(n13369[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4947_19_lut (.I0(GND_net), .I1(n14129[16]), .I2(GND_net), 
            .I3(n38597), .O(n13369[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_19 (.CI(n38597), .I0(n14129[16]), .I1(GND_net), 
            .CO(n38598));
    SB_LUT4 add_4947_18_lut (.I0(GND_net), .I1(n14129[15]), .I2(GND_net), 
            .I3(n38596), .O(n13369[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_18 (.CI(n38596), .I0(n14129[15]), .I1(GND_net), 
            .CO(n38597));
    SB_LUT4 add_4947_17_lut (.I0(GND_net), .I1(n14129[14]), .I2(GND_net), 
            .I3(n38595), .O(n13369[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_17 (.CI(n38595), .I0(n14129[14]), .I1(GND_net), 
            .CO(n38596));
    SB_LUT4 add_4947_16_lut (.I0(GND_net), .I1(n14129[13]), .I2(n1108_adj_4910), 
            .I3(n38594), .O(n13369[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_16 (.CI(n38594), .I0(n14129[13]), .I1(n1108_adj_4910), 
            .CO(n38595));
    SB_LUT4 add_4947_15_lut (.I0(GND_net), .I1(n14129[12]), .I2(n1035_adj_4909), 
            .I3(n38593), .O(n13369[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_15 (.CI(n38593), .I0(n14129[12]), .I1(n1035_adj_4909), 
            .CO(n38594));
    SB_LUT4 add_4947_14_lut (.I0(GND_net), .I1(n14129[11]), .I2(n962_adj_4907), 
            .I3(n38592), .O(n13369[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_14 (.CI(n38592), .I0(n14129[11]), .I1(n962_adj_4907), 
            .CO(n38593));
    SB_LUT4 add_958_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n4236[17]), .I3(n37605), .O(\PID_CONTROLLER.integral_23__N_3672 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_19 (.CI(n37605), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n4236[17]), .CO(n37606));
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_5132[7]), .I3(n37687), .O(n15_adj_4756)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_958_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n4236[16]), .I3(n37604), .O(\PID_CONTROLLER.integral_23__N_3672 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_18 (.CI(n37604), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n4236[16]), .CO(n37605));
    SB_LUT4 add_958_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n4236[15]), .I3(n37603), .O(\PID_CONTROLLER.integral_23__N_3672 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4947_13_lut (.I0(GND_net), .I1(n14129[10]), .I2(n889_adj_4902), 
            .I3(n38591), .O(n13369[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_13 (.CI(n38591), .I0(n14129[10]), .I1(n889_adj_4902), 
            .CO(n38592));
    SB_LUT4 add_4947_12_lut (.I0(GND_net), .I1(n14129[9]), .I2(n816_adj_4901), 
            .I3(n38590), .O(n13369[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_12 (.CI(n38590), .I0(n14129[9]), .I1(n816_adj_4901), 
            .CO(n38591));
    SB_LUT4 add_4947_11_lut (.I0(GND_net), .I1(n14129[8]), .I2(n743_adj_4899), 
            .I3(n38589), .O(n13369[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_11 (.CI(n38589), .I0(n14129[8]), .I1(n743_adj_4899), 
            .CO(n38590));
    SB_LUT4 add_4947_10_lut (.I0(GND_net), .I1(n14129[7]), .I2(n670_adj_4898), 
            .I3(n38588), .O(n13369[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_10 (.CI(n38588), .I0(n14129[7]), .I1(n670_adj_4898), 
            .CO(n38589));
    SB_LUT4 add_4947_9_lut (.I0(GND_net), .I1(n14129[6]), .I2(n597_adj_4897), 
            .I3(n38587), .O(n13369[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_9 (.CI(n38587), .I0(n14129[6]), .I1(n597_adj_4897), 
            .CO(n38588));
    SB_LUT4 add_4947_8_lut (.I0(GND_net), .I1(n14129[5]), .I2(n524_adj_4896), 
            .I3(n38586), .O(n13369[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_8 (.CI(n38586), .I0(n14129[5]), .I1(n524_adj_4896), 
            .CO(n38587));
    SB_LUT4 add_4947_7_lut (.I0(GND_net), .I1(n14129[4]), .I2(n451_adj_4895), 
            .I3(n38585), .O(n13369[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_7 (.CI(n38585), .I0(n14129[4]), .I1(n451_adj_4895), 
            .CO(n38586));
    SB_LUT4 add_4947_6_lut (.I0(GND_net), .I1(n14129[3]), .I2(n378_adj_4894), 
            .I3(n38584), .O(n13369[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_6 (.CI(n38584), .I0(n14129[3]), .I1(n378_adj_4894), 
            .CO(n38585));
    SB_LUT4 add_4947_5_lut (.I0(GND_net), .I1(n14129[2]), .I2(n305_adj_4893), 
            .I3(n38583), .O(n13369[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_5 (.CI(n38583), .I0(n14129[2]), .I1(n305_adj_4893), 
            .CO(n38584));
    SB_LUT4 add_4947_4_lut (.I0(GND_net), .I1(n14129[1]), .I2(n232_adj_4891), 
            .I3(n38582), .O(n13369[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_4 (.CI(n38582), .I0(n14129[1]), .I1(n232_adj_4891), 
            .CO(n38583));
    SB_LUT4 add_4947_3_lut (.I0(GND_net), .I1(n14129[0]), .I2(n159_adj_4890), 
            .I3(n38581), .O(n13369[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_3 (.CI(n38581), .I0(n14129[0]), .I1(n159_adj_4890), 
            .CO(n38582));
    SB_LUT4 add_4947_2_lut (.I0(GND_net), .I1(n17_adj_4887), .I2(n86_adj_4886), 
            .I3(GND_net), .O(n13369[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4947_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4947_2 (.CI(GND_net), .I0(n17_adj_4887), .I1(n86_adj_4886), 
            .CO(n38581));
    SB_LUT4 add_4984_19_lut (.I0(GND_net), .I1(n14813[16]), .I2(GND_net), 
            .I3(n38580), .O(n14129[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4984_18_lut (.I0(GND_net), .I1(n14813[15]), .I2(GND_net), 
            .I3(n38579), .O(n14129[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_18 (.CI(n38579), .I0(n14813[15]), .I1(GND_net), 
            .CO(n38580));
    SB_LUT4 add_4984_17_lut (.I0(GND_net), .I1(n14813[14]), .I2(GND_net), 
            .I3(n38578), .O(n14129[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_17 (.CI(n38578), .I0(n14813[14]), .I1(GND_net), 
            .CO(n38579));
    SB_LUT4 add_4984_16_lut (.I0(GND_net), .I1(n14813[13]), .I2(n1111_adj_4883), 
            .I3(n38577), .O(n14129[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_5117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32635_3_lut (.I0(n47766), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n47767));   // verilog/motorControl.v(31[10:34])
    defparam i32635_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_5116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_5115));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_5114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19997_2_lut (.I0(n28[19]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19997_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4984_16 (.CI(n38577), .I0(n14813[13]), .I1(n1111_adj_4883), 
            .CO(n38578));
    SB_LUT4 add_4984_15_lut (.I0(GND_net), .I1(n14813[12]), .I2(n1038_adj_4863), 
            .I3(n38576), .O(n14129[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_15 (.CI(n38576), .I0(n14813[12]), .I1(n1038_adj_4863), 
            .CO(n38577));
    SB_LUT4 add_4984_14_lut (.I0(GND_net), .I1(n14813[11]), .I2(n965_adj_4862), 
            .I3(n38575), .O(n14129[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_5112));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4984_14 (.CI(n38575), .I0(n14813[11]), .I1(n965_adj_4862), 
            .CO(n38576));
    SB_LUT4 add_4984_13_lut (.I0(GND_net), .I1(n14813[10]), .I2(n892_adj_4861), 
            .I3(n38574), .O(n14129[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_13 (.CI(n38574), .I0(n14813[10]), .I1(n892_adj_4861), 
            .CO(n38575));
    SB_LUT4 add_4984_12_lut (.I0(GND_net), .I1(n14813[9]), .I2(n819_adj_4860), 
            .I3(n38573), .O(n14129[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_12 (.CI(n38573), .I0(n14813[9]), .I1(n819_adj_4860), 
            .CO(n38574));
    SB_LUT4 add_4984_11_lut (.I0(GND_net), .I1(n14813[8]), .I2(n746_adj_4855), 
            .I3(n38572), .O(n14129[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_11 (.CI(n38572), .I0(n14813[8]), .I1(n746_adj_4855), 
            .CO(n38573));
    SB_LUT4 add_4984_10_lut (.I0(GND_net), .I1(n14813[7]), .I2(n673_adj_4853), 
            .I3(n38571), .O(n14129[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_10 (.CI(n38571), .I0(n14813[7]), .I1(n673_adj_4853), 
            .CO(n38572));
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_5111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4984_9_lut (.I0(GND_net), .I1(n14813[6]), .I2(n600_adj_4852), 
            .I3(n38570), .O(n14129[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_9 (.CI(n38570), .I0(n14813[6]), .I1(n600_adj_4852), 
            .CO(n38571));
    SB_LUT4 add_4984_8_lut (.I0(GND_net), .I1(n14813[5]), .I2(n527_adj_4849), 
            .I3(n38569), .O(n14129[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_8 (.CI(n38569), .I0(n14813[5]), .I1(n527_adj_4849), 
            .CO(n38570));
    SB_LUT4 add_4984_7_lut (.I0(GND_net), .I1(n14813[4]), .I2(n454_adj_4846), 
            .I3(n38568), .O(n14129[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_7 (.CI(n38568), .I0(n14813[4]), .I1(n454_adj_4846), 
            .CO(n38569));
    SB_LUT4 add_4984_6_lut (.I0(GND_net), .I1(n14813[3]), .I2(n381_adj_4843), 
            .I3(n38567), .O(n14129[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_6 (.CI(n38567), .I0(n14813[3]), .I1(n381_adj_4843), 
            .CO(n38568));
    SB_LUT4 add_4984_5_lut (.I0(GND_net), .I1(n14813[2]), .I2(n308_adj_4842), 
            .I3(n38566), .O(n14129[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_5 (.CI(n38566), .I0(n14813[2]), .I1(n308_adj_4842), 
            .CO(n38567));
    SB_LUT4 add_4984_4_lut (.I0(GND_net), .I1(n14813[1]), .I2(n235_adj_4840), 
            .I3(n38565), .O(n14129[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_4 (.CI(n38565), .I0(n14813[1]), .I1(n235_adj_4840), 
            .CO(n38566));
    SB_LUT4 add_4984_3_lut (.I0(GND_net), .I1(n14813[0]), .I2(n162_adj_4839), 
            .I3(n38564), .O(n14129[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_3 (.CI(n38564), .I0(n14813[0]), .I1(n162_adj_4839), 
            .CO(n38565));
    SB_LUT4 add_4984_2_lut (.I0(GND_net), .I1(n20_adj_4838), .I2(n89_adj_4836), 
            .I3(GND_net), .O(n14129[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4984_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n37687), .I0(GND_net), .I1(n1_adj_5132[7]), 
            .CO(n37688));
    SB_CARRY add_958_17 (.CI(n37603), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n4236[15]), .CO(n37604));
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_5110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_958_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n4236[14]), .I3(n37602), .O(\PID_CONTROLLER.integral_23__N_3672 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4984_2 (.CI(GND_net), .I0(n20_adj_4838), .I1(n89_adj_4836), 
            .CO(n38564));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_5132[6]), .I3(n37686), .O(n13_adj_4757)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5236_10_lut (.I0(GND_net), .I1(n18289[7]), .I2(n700_adj_4834), 
            .I3(n38563), .O(n18128[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_5109));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_5108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_5107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_958_16 (.CI(n37602), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n4236[14]), .CO(n37603));
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_5106));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19996_2_lut (.I0(n28[20]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19996_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19995_2_lut (.I0(n28[21]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19995_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n37686), .I0(GND_net), .I1(n1_adj_5132[6]), 
            .CO(n37687));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_5132[5]), .I3(n37685), .O(n11_adj_4758)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n37685), .I0(GND_net), .I1(n1_adj_5132[5]), 
            .CO(n37686));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_5132[4]), .I3(n37684), .O(n9_adj_4775)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5236_9_lut (.I0(GND_net), .I1(n18289[6]), .I2(n627_adj_4819), 
            .I3(n38562), .O(n18128[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n37684), .I0(GND_net), .I1(n1_adj_5132[4]), 
            .CO(n37685));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_5132[3]), .I3(n37683), .O(n7_adj_4792)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_958_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n4236[13]), .I3(n37601), .O(\PID_CONTROLLER.integral_23__N_3672 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_15 (.CI(n37601), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n4236[13]), .CO(n37602));
    SB_CARRY add_5236_9 (.CI(n38562), .I0(n18289[6]), .I1(n627_adj_4819), 
            .CO(n38563));
    SB_LUT4 add_958_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n4236[12]), .I3(n37600), .O(\PID_CONTROLLER.integral_23__N_3672 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_14 (.CI(n37600), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n4236[12]), .CO(n37601));
    SB_CARRY unary_minus_5_add_3_5 (.CI(n37683), .I0(GND_net), .I1(n1_adj_5132[3]), 
            .CO(n37684));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_5132[2]), .I3(n37682), .O(n5_adj_4793)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_958_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n4236[11]), .I3(n37599), .O(\PID_CONTROLLER.integral_23__N_3672 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n37682), .I0(GND_net), .I1(n1_adj_5132[2]), 
            .CO(n37683));
    SB_CARRY add_958_13 (.CI(n37599), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n4236[11]), .CO(n37600));
    SB_LUT4 add_958_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n4236[10]), .I3(n37598), .O(\PID_CONTROLLER.integral_23__N_3672 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5236_8_lut (.I0(GND_net), .I1(n18289[5]), .I2(n554_adj_4784), 
            .I3(n38561), .O(n18128[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_12 (.CI(n37598), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n4236[10]), .CO(n37599));
    SB_LUT4 add_958_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n4236[9]), .I3(n37597), .O(\PID_CONTROLLER.integral_23__N_3672 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_5132[1]), .I3(n37681), .O(n3_adj_4850)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_958_11 (.CI(n37597), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n4236[9]), .CO(n37598));
    SB_CARRY unary_minus_5_add_3_3 (.CI(n37681), .I0(GND_net), .I1(n1_adj_5132[1]), 
            .CO(n37682));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_5132[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3723 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_958_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n4236[8]), .I3(n37596), .O(\PID_CONTROLLER.integral_23__N_3672 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_10 (.CI(n37596), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n4236[8]), .CO(n37597));
    SB_LUT4 i23708_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .O(n18609[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23708_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_958_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n4236[7]), .I3(n37595), .O(\PID_CONTROLLER.integral_23__N_3672 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_958_9 (.CI(n37595), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n4236[7]), .CO(n37596));
    SB_LUT4 add_958_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n4236[6]), .I3(n37594), .O(\PID_CONTROLLER.integral_23__N_3672 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_8 (.CI(n38561), .I0(n18289[5]), .I1(n554_adj_4784), 
            .CO(n38562));
    SB_LUT4 add_5236_7_lut (.I0(GND_net), .I1(n18289[4]), .I2(n481_adj_4769), 
            .I3(n38560), .O(n18128[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_7 (.CI(n38560), .I0(n18289[4]), .I1(n481_adj_4769), 
            .CO(n38561));
    SB_LUT4 add_5236_6_lut (.I0(GND_net), .I1(n18289[3]), .I2(n408_adj_4768), 
            .I3(n38559), .O(n18128[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_6 (.CI(n38559), .I0(n18289[3]), .I1(n408_adj_4768), 
            .CO(n38560));
    SB_CARRY add_958_8 (.CI(n37594), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n4236[6]), .CO(n37595));
    SB_LUT4 add_5236_5_lut (.I0(GND_net), .I1(n18289[2]), .I2(n335_adj_4767), 
            .I3(n38558), .O(n18128[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_5 (.CI(n38558), .I0(n18289[2]), .I1(n335_adj_4767), 
            .CO(n38559));
    SB_LUT4 add_5236_4_lut (.I0(GND_net), .I1(n18289[1]), .I2(n262_adj_4766), 
            .I3(n38557), .O(n18128[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_4 (.CI(n38557), .I0(n18289[1]), .I1(n262_adj_4766), 
            .CO(n38558));
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_5132[0]), 
            .CO(n37681));
    SB_LUT4 add_5236_3_lut (.I0(GND_net), .I1(n18289[0]), .I2(n189_adj_4765), 
            .I3(n38556), .O(n18128[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_3 (.CI(n38556), .I0(n18289[0]), .I1(n189_adj_4765), 
            .CO(n38557));
    SB_LUT4 add_958_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n4236[5]), .I3(n37593), .O(\PID_CONTROLLER.integral_23__N_3672 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5236_2_lut (.I0(GND_net), .I1(n47_adj_4759), .I2(n116_adj_4755), 
            .I3(GND_net), .O(n18128[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_2 (.CI(GND_net), .I0(n47_adj_4759), .I1(n116_adj_4755), 
            .CO(n38556));
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n37680), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_18_lut (.I0(GND_net), .I1(n15425[15]), .I2(GND_net), 
            .I3(n38555), .O(n14813[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5019_17_lut (.I0(GND_net), .I1(n15425[14]), .I2(GND_net), 
            .I3(n38554), .O(n14813[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n37679), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n37679), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n37680));
    SB_CARRY add_5019_17 (.CI(n38554), .I0(n15425[14]), .I1(GND_net), 
            .CO(n38555));
    SB_LUT4 add_5019_16_lut (.I0(GND_net), .I1(n15425[13]), .I2(n1114_adj_4750), 
            .I3(n38553), .O(n14813[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n37678), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_5103));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_958_7 (.CI(n37593), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n4236[5]), .CO(n37594));
    SB_LUT4 add_958_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n4236[4]), .I3(n37592), .O(\PID_CONTROLLER.integral_23__N_3672 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_958_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_16 (.CI(n38553), .I0(n15425[13]), .I1(n1114_adj_4750), 
            .CO(n38554));
    SB_CARRY add_958_6 (.CI(n37592), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n4236[4]), .CO(n37593));
    SB_CARRY sub_3_add_2_23 (.CI(n37678), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n37679));
    SB_LUT4 add_5019_15_lut (.I0(GND_net), .I1(n15425[12]), .I2(n1041_adj_4748), 
            .I3(n38552), .O(n14813[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n37677), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5019_15 (.CI(n38552), .I0(n15425[12]), .I1(n1041_adj_4748), 
            .CO(n38553));
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_5102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5019_14_lut (.I0(GND_net), .I1(n15425[11]), .I2(n968_adj_4746), 
            .I3(n38551), .O(n14813[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_22 (.CI(n37677), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n37678));
    SB_CARRY add_5019_14 (.CI(n38551), .I0(n15425[11]), .I1(n968_adj_4746), 
            .CO(n38552));
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_5101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_5100));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5019_13_lut (.I0(GND_net), .I1(n15425[10]), .I2(n895_adj_4745), 
            .I3(n38550), .O(n14813[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_5099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_13 (.CI(n38550), .I0(n15425[10]), .I1(n895_adj_4745), 
            .CO(n38551));
    SB_LUT4 add_5019_12_lut (.I0(GND_net), .I1(n15425[9]), .I2(n822_adj_4744), 
            .I3(n38549), .O(n14813[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19994_2_lut (.I0(n28[22]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19994_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19993_2_lut (.I0(n28[23]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19993_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5019_12 (.CI(n38549), .I0(n15425[9]), .I1(n822_adj_4744), 
            .CO(n38550));
    SB_LUT4 add_5019_11_lut (.I0(GND_net), .I1(n15425[8]), .I2(n749), 
            .I3(n38548), .O(n14813[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5019_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4771));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4722));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_5097));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23822_2_lut_4_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(\Kp[1] ), 
            .I3(n28[19]), .O(n18633[0]));   // verilog/motorControl.v(34[16:22])
    defparam i23822_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_5095));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_5094));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_5093));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_5092));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_5091));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_5090));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_5089));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_5088));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_5087));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_5085));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_5080));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_5079));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_5078));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_5077));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_5075));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_5074));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_5073));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_5072));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_5071));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_5070));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_5069));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_5068));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_5067));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_5066));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_5065));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_5064));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_5062));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_5061));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_5060));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_5059));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_5058));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_5057));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_5056));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_5055));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_5054));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_5053));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_5052));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_5051));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_5050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_5049));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n28[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_5048));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_5047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_5046));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_5045));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_5044));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_5043));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_5132[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_5039));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_5037));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4763));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_5036));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_5035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_5034));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_5033));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31789_2_lut_4_lut (.I0(duty_23__N_3772[21]), .I1(n257[21]), 
            .I2(duty_23__N_3772[9]), .I3(n257[9]), .O(n46920));
    defparam i31789_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_5032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_5031));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4762));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_5029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4760));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31804_2_lut_4_lut (.I0(duty_23__N_3772[16]), .I1(n257[16]), 
            .I2(duty_23__N_3772[7]), .I3(n257[7]), .O(n46935));
    defparam i31804_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_5027));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_5026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4754));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_5023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4753));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_5022));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_5021));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_5020));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_5019));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326_adj_5018));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399_adj_5017));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_5016));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_5015));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_5014));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4918), .I1(\Kp[4] ), .I2(n18633[2]), 
            .I3(n28[18]), .O(n18584[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_5013));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4841));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(n28[19]), .I2(GND_net), 
            .I3(GND_net), .O(n204_adj_4942));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31831_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3772[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3772[9]), .O(n46962));
    defparam i31831_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i31844_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3772[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3772[7]), .O(n46975));
    defparam i31844_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i23693_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n18681[0]));   // verilog/motorControl.v(34[16:22])
    defparam i23693_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(n28[19]), .I2(GND_net), 
            .I3(GND_net), .O(n131_adj_4941));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(GND_net), 
            .I3(GND_net), .O(n62_adj_4940));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20014_2_lut (.I0(n28[2]), .I1(\PID_CONTROLLER.integral_23__N_3720 ), 
            .I2(GND_net), .I3(GND_net), .O(n4236[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20014_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32627_3_lut (.I0(n47767), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n47759));   // verilog/motorControl.v(31[10:34])
    defparam i32627_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i2_4_lut_adj_1551 (.I0(n4_adj_4988), .I1(\Kp[3] ), .I2(n18664[1]), 
            .I3(n28[19]), .O(n18633[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1551.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_5012));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1552 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n28[23]), 
            .I3(n28[20]), .O(n12_adj_5120));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1552.LUT_INIT = 16'h9c50;
    SB_LUT4 i23897_4_lut (.I0(n18633[2]), .I1(\Kp[4] ), .I2(n6_adj_4918), 
            .I3(n28[18]), .O(n8_adj_5121));   // verilog/motorControl.v(34[16:22])
    defparam i23897_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n28[19]), .I3(n28[21]), 
            .O(n11_adj_5122));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23843_4_lut (.I0(n18664[1]), .I1(\Kp[3] ), .I2(n4_adj_4988), 
            .I3(n28[19]), .O(n6_adj_5123));   // verilog/motorControl.v(34[16:22])
    defparam i23843_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i23695_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n37185));   // verilog/motorControl.v(34[16:22])
    defparam i23695_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_5123), .I1(n11_adj_5122), .I2(n8_adj_5121), 
            .I3(n12_adj_5120), .O(n18_adj_5124));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n28[18]), .I3(n28[22]), 
            .O(n13_adj_5125));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_5125), .I1(n18_adj_5124), .I2(n37185), 
            .I3(n4_adj_4934), .O(n44030));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_5011));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_5010));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_5007));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_5006));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_5004));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_5003));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1553 (.I0(n6_adj_4913), .I1(\Ki[4] ), .I2(n18609[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), .O(n18549[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1553.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1554 (.I0(n4_adj_4916), .I1(\Ki[3] ), .I2(n18649[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), .O(n18609[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1554.LUT_INIT = 16'h965a;
    SB_LUT4 i23853_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n18673[0]));   // verilog/motorControl.v(34[25:36])
    defparam i23853_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1555 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [20]), .O(n12_adj_5126));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1555.LUT_INIT = 16'h9c50;
    SB_LUT4 i23775_4_lut (.I0(n18609[2]), .I1(\Ki[4] ), .I2(n6_adj_4913), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [18]), .O(n8_adj_5127));   // verilog/motorControl.v(34[25:36])
    defparam i23775_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1556 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n11_adj_5128));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut_adj_1556.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23729_4_lut (.I0(n18649[1]), .I1(\Ki[3] ), .I2(n4_adj_4916), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [19]), .O(n6_adj_5129));   // verilog/motorControl.v(34[25:36])
    defparam i23729_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i23855_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [21]), .O(n37358));   // verilog/motorControl.v(34[25:36])
    defparam i23855_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1557 (.I0(n6_adj_5129), .I1(n11_adj_5128), .I2(n8_adj_5127), 
            .I3(n12_adj_5126), .O(n18_adj_5130));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut_adj_1557.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1558 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3672 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3672 [22]), .O(n13_adj_5131));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut_adj_1558.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1559 (.I0(n13_adj_5131), .I1(n18_adj_5130), .I2(n37358), 
            .I3(n4_adj_4911), .O(n43796));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut_adj_1559.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_5001));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5000));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4999));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4997));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4996));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4995));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4994));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4993));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4992));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4987));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4985));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4983));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4981));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4979));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4978));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4976));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4975));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4974));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4973));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4972));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4970));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685_adj_4969));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758_adj_4967));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831_adj_4966));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904_adj_4965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4964));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4963));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31972_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n48882), 
            .I2(IntegralLimit[21]), .I3(n47780), .O(n47103));
    defparam i31972_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4961));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4960));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4959));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4751));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4958));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4957));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4955));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4952));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4949));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4948));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4946));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4944));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4943));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4939));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4938));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4936));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4935));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4930));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4929));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i31829_3_lut_4_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3772[2]), .O(n46960));   // verilog/motorControl.v(38[19:35])
    defparam i31829_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4928));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4927));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4926));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3772[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4885));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4747));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4924));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3672 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4923));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4920));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module \grp_debouncer(3,1000) 
//

module \grp_debouncer(3,1000)  (reg_B, CLK_c, GND_net, VCC_net, data_i, 
            n28167, data_o, n44732, n28614, n28613);
    output [2:0]reg_B;
    input CLK_c;
    input GND_net;
    input VCC_net;
    input [2:0]data_i;
    input n28167;
    output [2:0]data_o;
    output n44732;
    input n28614;
    input n28613;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [9:0]n45;
    wire [9:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n38309, n38308, n38307, n38306, n38305, n38304, n38303, 
        n38302, n38301, cnt_next_9__N_812, n16, n17, n6;
    
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(CLK_c), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_2191_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[9]), 
            .I3(n38309), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_2191_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[8]), 
            .I3(n38308), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_10 (.CI(n38308), .I0(GND_net), .I1(cnt_reg[8]), 
            .CO(n38309));
    SB_LUT4 cnt_reg_2191_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[7]), 
            .I3(n38307), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_9 (.CI(n38307), .I0(GND_net), .I1(cnt_reg[7]), 
            .CO(n38308));
    SB_LUT4 cnt_reg_2191_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n38306), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_8 (.CI(n38306), .I0(GND_net), .I1(cnt_reg[6]), 
            .CO(n38307));
    SB_LUT4 cnt_reg_2191_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n38305), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_7 (.CI(n38305), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n38306));
    SB_LUT4 cnt_reg_2191_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n38304), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_6 (.CI(n38304), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n38305));
    SB_LUT4 cnt_reg_2191_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n38303), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_5 (.CI(n38303), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n38304));
    SB_LUT4 cnt_reg_2191_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n38302), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_4 (.CI(n38302), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n38303));
    SB_LUT4 cnt_reg_2191_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n38301), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_3 (.CI(n38301), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n38302));
    SB_LUT4 cnt_reg_2191_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_2191_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_2191_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n38301));
    SB_DFFSR cnt_reg_2191__i9 (.Q(cnt_reg[9]), .C(CLK_c), .D(n45[9]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i8 (.Q(cnt_reg[8]), .C(CLK_c), .D(n45[8]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i7 (.Q(cnt_reg[7]), .C(CLK_c), .D(n45[7]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i6 (.Q(cnt_reg[6]), .C(CLK_c), .D(n45[6]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i5 (.Q(cnt_reg[5]), .C(CLK_c), .D(n45[5]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i4 (.Q(cnt_reg[4]), .C(CLK_c), .D(n45[4]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i3 (.Q(cnt_reg[3]), .C(CLK_c), .D(n45[3]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i2 (.Q(cnt_reg[2]), .C(CLK_c), .D(n45[2]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_2191__i1 (.Q(cnt_reg[1]), .C(CLK_c), .D(n45[1]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i2 (.Q(reg_B[2]), .C(CLK_c), .D(reg_A[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(CLK_c), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(CLK_c), .D(data_i[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(CLK_c), .D(data_i[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_2191__i0 (.Q(cnt_reg[0]), .C(CLK_c), .D(n45[0]), 
            .R(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(CLK_c), .D(n28167));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 i6_4_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[7]), 
            .I3(cnt_reg[2]), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut (.I0(cnt_reg[4]), .I1(cnt_reg[3]), .I2(cnt_reg[8]), 
            .I3(cnt_reg[9]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(cnt_reg[6]), .I2(n16), .I3(cnt_reg[5]), 
            .O(n44732));
    defparam i9_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(reg_B[1]), .I2(reg_A[0]), .I3(reg_A[1]), 
            .O(n6));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut (.I0(n44732), .I1(n6), .I2(reg_B[2]), .I3(reg_A[2]), 
            .O(cnt_next_9__N_812));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i3_4_lut.LUT_INIT = 16'hdffd;
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(CLK_c), .D(n28614));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i2 (.Q(data_o[2]), .C(CLK_c), .D(n28613));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i2 (.Q(reg_A[2]), .C(CLK_c), .D(data_i[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (a_new, ENCODER1_B_N_keep, n1668, 
            ENCODER1_A_N_keep, encoder1_position, GND_net, VCC_net, 
            direction_N_3907, b_prev, n28480, n1673) /* synthesis lattice_noprune=1 */ ;
    output [1:0]a_new;
    input ENCODER1_B_N_keep;
    input n1668;
    input ENCODER1_A_N_keep;
    output [31:0]encoder1_position;
    input GND_net;
    input VCC_net;
    output direction_N_3907;
    output b_prev;
    input n28480;
    output n1673;
    
    
    wire debounce_cnt, a_prev_N_3913, a_prev, n28388;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [31:0]n133;
    
    wire direction_N_3906, n38347, n38346, n38345, n38344, n38343, 
        n38342, n38341, n38340, n38339, n38338, n38337, n38336, 
        n38335, n38334, n38333, n38332, n38331, n38330, n38329, 
        n38328, n38327, n38326, n38325, n38324, n38323, n38322, 
        n38321, n38320, n38319, n38318, n38317, direction_N_3910, 
        n28481;
    
    SB_LUT4 i14874_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(a_new[1]), 
            .I3(a_prev), .O(n28388));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14874_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1668), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1668), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2193_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[31]), .I3(n38347), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2193_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[30]), .I3(n38346), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_32 (.CI(n38346), .I0(direction_N_3906), 
            .I1(encoder1_position[30]), .CO(n38347));
    SB_LUT4 position_2193_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[29]), .I3(n38345), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_31 (.CI(n38345), .I0(direction_N_3906), 
            .I1(encoder1_position[29]), .CO(n38346));
    SB_LUT4 position_2193_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[28]), .I3(n38344), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_30 (.CI(n38344), .I0(direction_N_3906), 
            .I1(encoder1_position[28]), .CO(n38345));
    SB_LUT4 position_2193_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[27]), .I3(n38343), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1668), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_CARRY position_2193_add_4_29 (.CI(n38343), .I0(direction_N_3906), 
            .I1(encoder1_position[27]), .CO(n38344));
    SB_LUT4 position_2193_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[26]), .I3(n38342), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_28 (.CI(n38342), .I0(direction_N_3906), 
            .I1(encoder1_position[26]), .CO(n38343));
    SB_LUT4 position_2193_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[25]), .I3(n38341), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_27 (.CI(n38341), .I0(direction_N_3906), 
            .I1(encoder1_position[25]), .CO(n38342));
    SB_LUT4 position_2193_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[24]), .I3(n38340), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_26 (.CI(n38340), .I0(direction_N_3906), 
            .I1(encoder1_position[24]), .CO(n38341));
    SB_LUT4 position_2193_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[23]), .I3(n38339), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_25 (.CI(n38339), .I0(direction_N_3906), 
            .I1(encoder1_position[23]), .CO(n38340));
    SB_LUT4 position_2193_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[22]), .I3(n38338), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_24 (.CI(n38338), .I0(direction_N_3906), 
            .I1(encoder1_position[22]), .CO(n38339));
    SB_LUT4 position_2193_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[21]), .I3(n38337), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_23 (.CI(n38337), .I0(direction_N_3906), 
            .I1(encoder1_position[21]), .CO(n38338));
    SB_LUT4 position_2193_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[20]), .I3(n38336), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_22 (.CI(n38336), .I0(direction_N_3906), 
            .I1(encoder1_position[20]), .CO(n38337));
    SB_LUT4 position_2193_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[19]), .I3(n38335), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_21 (.CI(n38335), .I0(direction_N_3906), 
            .I1(encoder1_position[19]), .CO(n38336));
    SB_LUT4 position_2193_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[18]), .I3(n38334), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_20 (.CI(n38334), .I0(direction_N_3906), 
            .I1(encoder1_position[18]), .CO(n38335));
    SB_LUT4 position_2193_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[17]), .I3(n38333), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_19 (.CI(n38333), .I0(direction_N_3906), 
            .I1(encoder1_position[17]), .CO(n38334));
    SB_LUT4 position_2193_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[16]), .I3(n38332), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_18 (.CI(n38332), .I0(direction_N_3906), 
            .I1(encoder1_position[16]), .CO(n38333));
    SB_LUT4 position_2193_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[15]), .I3(n38331), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_17 (.CI(n38331), .I0(direction_N_3906), 
            .I1(encoder1_position[15]), .CO(n38332));
    SB_LUT4 position_2193_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[14]), .I3(n38330), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_16 (.CI(n38330), .I0(direction_N_3906), 
            .I1(encoder1_position[14]), .CO(n38331));
    SB_LUT4 position_2193_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[13]), .I3(n38329), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_15 (.CI(n38329), .I0(direction_N_3906), 
            .I1(encoder1_position[13]), .CO(n38330));
    SB_LUT4 position_2193_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[12]), .I3(n38328), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_14 (.CI(n38328), .I0(direction_N_3906), 
            .I1(encoder1_position[12]), .CO(n38329));
    SB_LUT4 position_2193_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[11]), .I3(n38327), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_13 (.CI(n38327), .I0(direction_N_3906), 
            .I1(encoder1_position[11]), .CO(n38328));
    SB_LUT4 position_2193_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[10]), .I3(n38326), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_12 (.CI(n38326), .I0(direction_N_3906), 
            .I1(encoder1_position[10]), .CO(n38327));
    SB_LUT4 position_2193_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[9]), .I3(n38325), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_11 (.CI(n38325), .I0(direction_N_3906), 
            .I1(encoder1_position[9]), .CO(n38326));
    SB_LUT4 position_2193_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[8]), .I3(n38324), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_10 (.CI(n38324), .I0(direction_N_3906), 
            .I1(encoder1_position[8]), .CO(n38325));
    SB_LUT4 position_2193_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[7]), .I3(n38323), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_9 (.CI(n38323), .I0(direction_N_3906), 
            .I1(encoder1_position[7]), .CO(n38324));
    SB_LUT4 position_2193_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[6]), .I3(n38322), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_8 (.CI(n38322), .I0(direction_N_3906), 
            .I1(encoder1_position[6]), .CO(n38323));
    SB_LUT4 position_2193_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[5]), .I3(n38321), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_7 (.CI(n38321), .I0(direction_N_3906), 
            .I1(encoder1_position[5]), .CO(n38322));
    SB_LUT4 position_2193_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[4]), .I3(n38320), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_6 (.CI(n38320), .I0(direction_N_3906), 
            .I1(encoder1_position[4]), .CO(n38321));
    SB_LUT4 position_2193_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[3]), .I3(n38319), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_5 (.CI(n38319), .I0(direction_N_3906), 
            .I1(encoder1_position[3]), .CO(n38320));
    SB_LUT4 position_2193_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[2]), .I3(n38318), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_4 (.CI(n38318), .I0(direction_N_3906), 
            .I1(encoder1_position[2]), .CO(n38319));
    SB_LUT4 position_2193_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder1_position[1]), .I3(n38317), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_3 (.CI(n38317), .I0(direction_N_3906), 
            .I1(encoder1_position[1]), .CO(n38318));
    SB_LUT4 position_2193_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2193_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2193_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n38317));
    SB_DFFE position_2193__i31 (.Q(encoder1_position[31]), .C(n1668), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i30 (.Q(encoder1_position[30]), .C(n1668), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i29 (.Q(encoder1_position[29]), .C(n1668), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i28 (.Q(encoder1_position[28]), .C(n1668), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i27 (.Q(encoder1_position[27]), .C(n1668), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i26 (.Q(encoder1_position[26]), .C(n1668), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i25 (.Q(encoder1_position[25]), .C(n1668), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i24 (.Q(encoder1_position[24]), .C(n1668), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i23 (.Q(encoder1_position[23]), .C(n1668), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i22 (.Q(encoder1_position[22]), .C(n1668), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i21 (.Q(encoder1_position[21]), .C(n1668), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i20 (.Q(encoder1_position[20]), .C(n1668), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i19 (.Q(encoder1_position[19]), .C(n1668), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i18 (.Q(encoder1_position[18]), .C(n1668), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i17 (.Q(encoder1_position[17]), .C(n1668), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i16 (.Q(encoder1_position[16]), .C(n1668), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i15 (.Q(encoder1_position[15]), .C(n1668), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i14 (.Q(encoder1_position[14]), .C(n1668), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i13 (.Q(encoder1_position[13]), .C(n1668), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i12 (.Q(encoder1_position[12]), .C(n1668), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i11 (.Q(encoder1_position[11]), .C(n1668), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i10 (.Q(encoder1_position[10]), .C(n1668), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i9 (.Q(encoder1_position[9]), .C(n1668), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i8 (.Q(encoder1_position[8]), .C(n1668), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i7 (.Q(encoder1_position[7]), .C(n1668), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i6 (.Q(encoder1_position[6]), .C(n1668), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i5 (.Q(encoder1_position[5]), .C(n1668), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i4 (.Q(encoder1_position[4]), .C(n1668), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i3 (.Q(encoder1_position[3]), .C(n1668), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i2 (.Q(encoder1_position[2]), .C(n1668), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i1 (.Q(encoder1_position[1]), .C(n1668), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2193__i0 (.Q(encoder1_position[0]), .C(n1668), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1668), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1668), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(a_new[1]), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1668), .D(n28481));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1673), .C(n1668), .D(n28480));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1668), .D(n28388));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i32748_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i32748_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i14967_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n28481));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14967_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (CLK_c, read, \state[0] , enable_slow_N_4190, n5614, 
            \state[1] , n41883, n41869, n28229, rw, n41973, data_ready, 
            \state[3] , n6, GND_net, \state[2] , n7, n33881, n43114, 
            n42289, scl_enable, scl, \state_7__N_4103[3] , \state[0]_adj_13 , 
            n33185, n6692, \saved_addr[0] , VCC_net, n4, n4_adj_14, 
            n33292, sda_enable, \state_7__N_4087[0] , n28193, data, 
            n28192, n28191, n28190, n28189, n28188, n28187, n10, 
            n8, n28330, n28315, n7233, n26424, n26409, sda_out, 
            n46890) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    input read;
    output \state[0] ;
    output enable_slow_N_4190;
    output [0:0]n5614;
    output \state[1] ;
    input n41883;
    input n41869;
    input n28229;
    output rw;
    input n41973;
    output data_ready;
    output \state[3] ;
    output n6;
    input GND_net;
    output \state[2] ;
    output n7;
    output n33881;
    input n43114;
    output n42289;
    output scl_enable;
    output scl;
    input \state_7__N_4103[3] ;
    output \state[0]_adj_13 ;
    output n33185;
    output n6692;
    output \saved_addr[0] ;
    input VCC_net;
    output n4;
    output n4_adj_14;
    output n33292;
    output sda_enable;
    output \state_7__N_4087[0] ;
    input n28193;
    output [7:0]data;
    input n28192;
    input n28191;
    input n28190;
    input n28189;
    input n28188;
    input n28187;
    output n10;
    input n8;
    input n28330;
    input n28315;
    input n7233;
    output n26424;
    output n26409;
    output sda_out;
    output n46890;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3989;
    
    wire n27777;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n28001, n28, n26, n27, n25, n26287, enable;
    wire [15:0]n4272;
    
    wire n37626, n37625, n37624, n37623, n37622, n37621, n37620, 
        n37619, n37618, n37617, n37616, n37615, n37614, n37613, 
        n37612;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[1]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[2]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[3]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[4]), .S(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[5]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[6]), .S(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[7]), .S(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[8]), .S(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[9]), .S(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[10]), .S(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[11]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[12]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n26287));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_1410_Mux_0_i1_4_lut (.I0(read), .I1(n26287), .I2(\state[0] ), 
            .I3(enable_slow_N_4190), .O(n5614[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_1410_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[13]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n5614[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[14]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[15]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n27777), 
            .D(delay_counter_15__N_3989[0]), .R(n28001));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n41883));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n41869));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n28229));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n41973));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i2_2_lut (.I0(n26287), .I1(\state[3] ), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14500_2_lut (.I0(n27777), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28001));   // verilog/eeprom.v(26[8] 58[4])
    defparam i14500_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n27777));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 add_962_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n4272[15]), 
            .I3(n37626), .O(delay_counter_15__N_3989[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_962_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n4272[15]), 
            .I3(n37625), .O(delay_counter_15__N_3989[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_16 (.CI(n37625), .I0(delay_counter[14]), .I1(n4272[15]), 
            .CO(n37626));
    SB_LUT4 add_962_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n4272[15]), 
            .I3(n37624), .O(delay_counter_15__N_3989[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_15 (.CI(n37624), .I0(delay_counter[13]), .I1(n4272[15]), 
            .CO(n37625));
    SB_LUT4 add_962_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n4272[15]), 
            .I3(n37623), .O(delay_counter_15__N_3989[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_14 (.CI(n37623), .I0(delay_counter[12]), .I1(n4272[15]), 
            .CO(n37624));
    SB_LUT4 add_962_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n4272[15]), 
            .I3(n37622), .O(delay_counter_15__N_3989[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_13 (.CI(n37622), .I0(delay_counter[11]), .I1(n4272[15]), 
            .CO(n37623));
    SB_LUT4 add_962_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n4272[15]), 
            .I3(n37621), .O(delay_counter_15__N_3989[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_12 (.CI(n37621), .I0(delay_counter[10]), .I1(n4272[15]), 
            .CO(n37622));
    SB_LUT4 add_962_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n4272[15]), 
            .I3(n37620), .O(delay_counter_15__N_3989[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_11 (.CI(n37620), .I0(delay_counter[9]), .I1(n4272[15]), 
            .CO(n37621));
    SB_LUT4 add_962_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n4272[15]), 
            .I3(n37619), .O(delay_counter_15__N_3989[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_10 (.CI(n37619), .I0(delay_counter[8]), .I1(n4272[15]), 
            .CO(n37620));
    SB_LUT4 add_962_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n4272[15]), 
            .I3(n37618), .O(delay_counter_15__N_3989[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_9 (.CI(n37618), .I0(delay_counter[7]), .I1(n4272[15]), 
            .CO(n37619));
    SB_LUT4 add_962_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n4272[15]), 
            .I3(n37617), .O(delay_counter_15__N_3989[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_8 (.CI(n37617), .I0(delay_counter[6]), .I1(n4272[15]), 
            .CO(n37618));
    SB_LUT4 add_962_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n4272[15]), 
            .I3(n37616), .O(delay_counter_15__N_3989[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_7 (.CI(n37616), .I0(delay_counter[5]), .I1(n4272[15]), 
            .CO(n37617));
    SB_LUT4 add_962_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n4272[15]), 
            .I3(n37615), .O(delay_counter_15__N_3989[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_6 (.CI(n37615), .I0(delay_counter[4]), .I1(n4272[15]), 
            .CO(n37616));
    SB_LUT4 add_962_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n4272[15]), 
            .I3(n37614), .O(delay_counter_15__N_3989[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_5 (.CI(n37614), .I0(delay_counter[3]), .I1(n4272[15]), 
            .CO(n37615));
    SB_LUT4 add_962_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n4272[15]), 
            .I3(n37613), .O(delay_counter_15__N_3989[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_4 (.CI(n37613), .I0(delay_counter[2]), .I1(n4272[15]), 
            .CO(n37614));
    SB_LUT4 add_962_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n4272[15]), 
            .I3(n37612), .O(delay_counter_15__N_3989[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_3 (.CI(n37612), .I0(delay_counter[1]), .I1(n4272[15]), 
            .CO(n37613));
    SB_LUT4 add_962_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n4272[15]), 
            .I3(GND_net), .O(delay_counter_15__N_3989[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_962_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_962_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n4272[15]), 
            .CO(n37612));
    SB_LUT4 i2_2_lut_adj_1543 (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut_adj_1543.LUT_INIT = 16'heeee;
    SB_LUT4 i20376_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4190), 
            .I3(GND_net), .O(n33881));   // verilog/eeprom.v(51[5:9])
    defparam i20376_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4190), 
            .I3(n43114), .O(n42289));   // verilog/eeprom.v(51[5:9])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 i32793_2_lut (.I0(n26287), .I1(enable_slow_N_4190), .I2(GND_net), 
            .I3(GND_net), .O(n4272[15]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i32793_2_lut.LUT_INIT = 16'h2222;
    i2c_controller i2c (.scl_enable(scl_enable), .scl(scl), .GND_net(GND_net), 
            .\state_7__N_4103[3] (\state_7__N_4103[3] ), .\state[0] (\state[0]_adj_13 ), 
            .\state[1] (state[1]), .\state[2] (\state[2] ), .\state[3] (\state[3] ), 
            .n33185(n33185), .n6692(n6692), .\saved_addr[0] (\saved_addr[0] ), 
            .CLK_c(CLK_c), .VCC_net(VCC_net), .n4(n4), .n4_adj_12(n4_adj_14), 
            .n33292(n33292), .sda_enable(sda_enable), .\state_7__N_4087[0] (\state_7__N_4087[0] ), 
            .n28193(n28193), .data({data}), .n28192(n28192), .n28191(n28191), 
            .n28190(n28190), .n28189(n28189), .n28188(n28188), .n28187(n28187), 
            .n10(n10), .enable(enable), .enable_slow_N_4190(enable_slow_N_4190), 
            .n8(n8), .n28330(n28330), .n28315(n28315), .n7233(n7233), 
            .n26424(n26424), .n26409(n26409), .sda_out(sda_out), .n46890(n46890)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (scl_enable, scl, GND_net, \state_7__N_4103[3] , 
            \state[0] , \state[1] , \state[2] , \state[3] , n33185, 
            n6692, \saved_addr[0] , CLK_c, VCC_net, n4, n4_adj_12, 
            n33292, sda_enable, \state_7__N_4087[0] , n28193, data, 
            n28192, n28191, n28190, n28189, n28188, n28187, n10, 
            enable, enable_slow_N_4190, n8, n28330, n28315, n7233, 
            n26424, n26409, sda_out, n46890) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output scl_enable;
    output scl;
    input GND_net;
    input \state_7__N_4103[3] ;
    output \state[0] ;
    output \state[1] ;
    output \state[2] ;
    output \state[3] ;
    output n33185;
    output n6692;
    output \saved_addr[0] ;
    input CLK_c;
    input VCC_net;
    output n4;
    output n4_adj_12;
    output n33292;
    output sda_enable;
    output \state_7__N_4087[0] ;
    input n28193;
    output [7:0]data;
    input n28192;
    input n28191;
    input n28190;
    input n28189;
    input n28188;
    input n28187;
    output n10;
    input enable;
    output enable_slow_N_4190;
    input n8;
    input n28330;
    input n28315;
    input n7233;
    output n26424;
    output n26409;
    output sda_out;
    output n46890;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n11, n33476, n9, n10_c, state_7__N_4086, n6685, n11_adj_4695, 
        n11_adj_4696, n5;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n46843, n46827, n6502;
    wire [0:0]n6538;
    
    wire n28015, i2c_clk_N_4176, n7, n33, n37, n27999, n34, n39, 
        n7136, n19183;
    wire [7:0]n119;
    
    wire n27820, n28070;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n38415, n38414, n38413, n38412, n38411, scl_enable_N_4177, 
        n41911, sda_out_adj_4700, n33966, n33485, n42053, n44346, 
        enable_slow_N_4189, n27745, n37765, n37764, n37763, n37762, 
        n37761, n37760, n37759, n10_adj_4701, n12, n10_adj_4703, 
        n11_adj_4704, n15, n43122, n46897;
    
    SB_LUT4 i19777_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i19777_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i33082_2_lut (.I0(\state_7__N_4103[3] ), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n33476));
    defparam i33082_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_c));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i32700_4_lut (.I0(state_7__N_4086), .I1(n6685), .I2(n11_adj_4695), 
            .I3(n33185), .O(n6692));
    defparam i32700_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_4_lut (.I0(n11_adj_4696), .I1(n11), .I2(\state_7__N_4103[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'h5755;
    SB_LUT4 i31850_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n46843));   // verilog/i2c_controller.v(198[28:35])
    defparam i31850_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31802_4_lut (.I0(n46843), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n46827));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i31802_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 mux_1621_i1_4_lut (.I0(n46827), .I1(\state[0] ), .I2(n6502), 
            .I3(\state[2] ), .O(n6538[0]));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam mux_1621_i1_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i1_2_lut (.I0(i2c_clk), .I1(n28015), .I2(GND_net), .I3(GND_net), 
            .O(i2c_clk_N_4176));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1537 (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1537.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n27999));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_1538 (.I0(n34), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i1_2_lut_adj_1538.LUT_INIT = 16'heeee;
    SB_LUT4 i32800_4_lut (.I0(n6502), .I1(n39), .I2(\state[2] ), .I3(\state[1] ), 
            .O(n7136));
    defparam i32800_4_lut.LUT_INIT = 16'hc8cc;
    SB_LUT4 i32795_2_lut (.I0(\state[0] ), .I1(n6502), .I2(GND_net), .I3(GND_net), 
            .O(n19183));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i32795_2_lut.LUT_INIT = 16'h4444;
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27820), .D(n119[1]), 
            .S(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27820), .D(n119[2]), 
            .S(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27820), .D(n119[3]), 
            .R(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27820), .D(n119[4]), 
            .R(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27820), .D(n119[5]), 
            .R(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27820), .D(n119[6]), 
            .R(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27820), .D(n119[7]), 
            .R(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_2203_2204__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n28015));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 counter2_2203_2204_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n38415), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_2203_2204_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n38414), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_6 (.CI(n38414), .I0(GND_net), .I1(counter2[4]), 
            .CO(n38415));
    SB_LUT4 counter2_2203_2204_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n38413), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_5 (.CI(n38413), .I0(GND_net), .I1(counter2[3]), 
            .CO(n38414));
    SB_LUT4 counter2_2203_2204_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n38412), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_4 (.CI(n38412), .I0(GND_net), .I1(counter2[2]), 
            .CO(n38413));
    SB_LUT4 counter2_2203_2204_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n38411), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_3 (.CI(n38411), .I0(GND_net), .I1(counter2[1]), 
            .CO(n38412));
    SB_LUT4 counter2_2203_2204_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_2203_2204_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_2203_2204_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n38411));
    SB_LUT4 equal_340_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_340_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_339_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_12));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_339_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i19795_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33292));
    defparam i19795_2_lut.LUT_INIT = 16'h8888;
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n7136), 
            .D(n19183), .S(n27999));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4176));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4177));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4700), .C(i2c_clk), .E(n41911), 
            .D(n6538[0]));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27820), .D(n119[0]), 
            .S(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n6692), .D(n5), 
            .S(n33966));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n6692), .D(n33476), 
            .S(n33485));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n6692), .D(n42053), 
            .S(n44346));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE enable_slow_120 (.Q(\state_7__N_4087[0] ), .C(CLK_c), .E(n27745), 
            .D(enable_slow_N_4189));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n37765), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n37764), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n37764), .I0(counter[6]), .I1(VCC_net), 
            .CO(n37765));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n37763), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n37763), .I0(counter[5]), .I1(VCC_net), 
            .CO(n37764));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n37762), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n37762), .I0(counter[4]), .I1(VCC_net), 
            .CO(n37763));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n37761), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n37761), .I0(counter[3]), .I1(VCC_net), 
            .CO(n37762));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n37760), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n37760), .I0(counter[2]), .I1(VCC_net), 
            .CO(n37761));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n37759), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_3 (.CI(n37759), .I0(counter[1]), .I1(VCC_net), 
            .CO(n37760));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n37759));
    SB_DFFSR counter2_2203_2204__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n28015));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2203_2204__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n28015));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2203_2204__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n28015));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2203_2204__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n28015));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_2203_2204__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n28015));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n28193));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n28192));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n28191));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n28190));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n28189));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n28188));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n28187));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4701));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4701), .I2(counter2[0]), 
            .I3(GND_net), .O(n28015));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i32798_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n41911));
    defparam i32798_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i33085_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n6692), .O(n44346));
    defparam i33085_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n6685));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_264_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4703));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_264_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut (.I0(enable), .I1(\state_7__N_4087[0] ), .I2(enable_slow_N_4190), 
            .I3(GND_net), .O(n27745));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i33087_3_lut_4_lut (.I0(n9), .I1(n10_c), .I2(n11_adj_4704), 
            .I3(n6692), .O(n33485));   // verilog/i2c_controller.v(151[5:14])
    defparam i33087_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i28099_2_lut (.I0(\state_7__N_4103[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n43122));
    defparam i28099_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n28330));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4704));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n28315));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i17_4_lut (.I0(n6685), .I1(n43122), .I2(n7233), .I3(n37), 
            .O(n27820));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 equal_2182_i19_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4190));   // verilog/i2c_controller.v(77[47:62])
    defparam equal_2182_i19_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i28065_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n43122), .O(n28070));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i28065_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 equal_264_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_264_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4696));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 i1_2_lut_3_lut_adj_1539 (.I0(n9), .I1(n10_c), .I2(counter[0]), 
            .I3(GND_net), .O(n26424));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_1539.LUT_INIT = 16'hefef;
    SB_LUT4 i20340_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4177));   // verilog/i2c_controller.v(77[47:62])
    defparam i20340_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i3_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(\state[2] ), .O(n6502));   // verilog/i2c_controller.v(77[47:62])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h001a;
    SB_LUT4 i1_2_lut_3_lut_adj_1540 (.I0(n9), .I1(n10_c), .I2(counter[0]), 
            .I3(GND_net), .O(n26409));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_1540.LUT_INIT = 16'hfefe;
    SB_LUT4 i2604_2_lut (.I0(sda_out_adj_4700), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i2604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i32687_2_lut (.I0(\state_7__N_4087[0] ), .I1(enable_slow_N_4190), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4189));   // verilog/i2c_controller.v(62[6:32])
    defparam i32687_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut_4_lut_adj_1541 (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut_adj_1541.LUT_INIT = 16'h0510;
    SB_LUT4 i31820_3_lut_4_lut (.I0(n11_adj_4695), .I1(n11_adj_4704), .I2(enable_slow_N_4190), 
            .I3(\state_7__N_4087[0] ), .O(n46890));
    defparam i31820_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i33089_3_lut_4_lut (.I0(n11_adj_4695), .I1(n11_adj_4704), .I2(n15), 
            .I3(n6692), .O(n33966));
    defparam i33089_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i31999_4_lut (.I0(n10_adj_4703), .I1(n10_c), .I2(\state_7__N_4103[3] ), 
            .I3(enable), .O(n46897));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i31999_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut_adj_1542 (.I0(\state[1] ), .I1(n7), .I2(n46897), 
            .I3(\state[0] ), .O(n42053));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_1542.LUT_INIT = 16'ha088;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4695));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i19817_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33185));
    defparam i19817_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i20360_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_4086));
    defparam i20360_3_lut_4_lut.LUT_INIT = 16'hf800;
    
endmodule
//
// Verilog Description of module TLI4970
//

module TLI4970 (GND_net, CS_c, CS_CLK_c, n5, n5_adj_11, n33328, 
            CLK_c, VCC_net, \data[15] , n43722, n28227, current, 
            n28692, n28691, n28690, n28689, n28688, n28687, n28686, 
            n28685, n28684, n28683, n28682, n28681, n28185, n28184, 
            \data[12] , n28183, \data[11] , n28182, \data[10] , n28181, 
            \data[9] , n28180, \data[8] , n28179, \data[7] , n28178, 
            \data[6] , n28177, \data[5] , n28176, \data[4] , n28175, 
            \data[3] , n28174, \data[2] , n28173, \data[1] , state_7__N_4293, 
            n28458, \data[0] , n9, n11, n26432, n26440, n26445, 
            n26435) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    output CS_c;
    output CS_CLK_c;
    output n5;
    output n5_adj_11;
    output n33328;
    input CLK_c;
    input VCC_net;
    output \data[15] ;
    output n43722;
    input n28227;
    output [12:0]current;
    input n28692;
    input n28691;
    input n28690;
    input n28689;
    input n28688;
    input n28687;
    input n28686;
    input n28685;
    input n28684;
    input n28683;
    input n28682;
    input n28681;
    input n28185;
    input n28184;
    output \data[12] ;
    input n28183;
    output \data[11] ;
    input n28182;
    output \data[10] ;
    input n28181;
    output \data[9] ;
    input n28180;
    output \data[8] ;
    input n28179;
    output \data[7] ;
    input n28178;
    output \data[6] ;
    input n28177;
    output \data[5] ;
    input n28176;
    output \data[4] ;
    input n28175;
    output \data[3] ;
    input n28174;
    output \data[2] ;
    input n28173;
    output \data[1] ;
    output state_7__N_4293;
    input n28458;
    output \data[0] ;
    output n9;
    output n11;
    output n26432;
    output n26440;
    output n26445;
    output n26435;
    
    wire clk_slow /* synthesis is_clock=1, SET_AS_NETWORK=\tli/clk_slow */ ;   // verilog/tli4970.v(11[7:15])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n10078, n27869;
    wire [7:0]state;   // verilog/tli4970.v(29[13:18])
    
    wire n27983;
    wire [7:0]n37;
    
    wire n27779;
    wire [7:0]bit_counter;   // verilog/tli4970.v(26[13:24])
    
    wire n28035;
    wire [7:0]counter;   // verilog/tli4970.v(12[13:20])
    
    wire n6, clk_slow_N_4207, clk_slow_N_4206, clk_out;
    wire [4:0]n25;
    
    wire n38364, n38363, n38362, n38361;
    wire [13:0]n61;
    wire [15:0]delay_counter;   // verilog/tli4970.v(28[14:27])
    
    wire n38360, n38359, n38358, n38357, n38356, n38355, n38354, 
        n38353, n38352, n38351, n38350, n38349, n38348, n46880, 
        n23333, n38316, n38315, n38314, n38313, n46832, n38312, 
        n1, n46831, n38311, n46830, n38310, n33707, delay_counter_15__N_4288, 
        n23302, n23304, n23306, n9_c, n28230, n15, n6_adj_4693, 
        n6_adj_4694, n43806, n43723, n44313;
    
    SB_DFFNESR state_i1 (.Q(state[1]), .C(clk_slow), .E(n27869), .D(n10078), 
            .R(n27983));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNESR bit_counter_2192__i4 (.Q(bit_counter[4]), .C(clk_slow), .E(n27779), 
            .D(n37[4]), .R(n28035));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2192__i5 (.Q(bit_counter[5]), .C(clk_slow), .E(n27779), 
            .D(n37[5]), .R(n28035));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2192__i6 (.Q(bit_counter[6]), .C(clk_slow), .E(n27779), 
            .D(n37[6]), .R(n28035));   // verilog/tli4970.v(53[24:39])
    SB_DFFNESR bit_counter_2192__i7 (.Q(bit_counter[7]), .C(clk_slow), .E(n27779), 
            .D(n37[7]), .R(n28035));   // verilog/tli4970.v(53[24:39])
    SB_LUT4 i2_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2298_4_lut (.I0(counter[0]), .I1(counter[4]), .I2(n6), .I3(counter[3]), 
            .O(clk_slow_N_4207));
    defparam i2298_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 clk_slow_I_0_71_2_lut (.I0(clk_slow), .I1(clk_slow_N_4207), 
            .I2(GND_net), .I3(GND_net), .O(clk_slow_N_4206));   // verilog/tli4970.v(15[5] 18[8])
    defparam clk_slow_I_0_71_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 spi_clk_I_0_i1_3_lut (.I0(clk_slow), .I1(clk_out), .I2(CS_c), 
            .I3(GND_net), .O(CS_CLK_c));   // verilog/tli4970.v(23[20:53])
    defparam spi_clk_I_0_i1_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 equal_314_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/tli4970.v(52[9:26])
    defparam equal_314_i5_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_313_i5_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_11));   // verilog/tli4970.v(52[9:26])
    defparam equal_313_i5_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i19830_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n33328));
    defparam i19830_2_lut.LUT_INIT = 16'h8888;
    SB_DFF clk_slow_62 (.Q(clk_slow), .C(CLK_c), .D(clk_slow_N_4206));   // verilog/tli4970.v(13[10] 19[6])
    SB_LUT4 counter_2196_2197_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(counter[4]), 
            .I3(n38364), .O(n25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter_2196_2197_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(counter[3]), 
            .I3(n38363), .O(n25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_5 (.CI(n38363), .I0(GND_net), .I1(counter[3]), 
            .CO(n38364));
    SB_LUT4 counter_2196_2197_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(counter[2]), 
            .I3(n38362), .O(n25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_4 (.CI(n38362), .I0(GND_net), .I1(counter[2]), 
            .CO(n38363));
    SB_LUT4 counter_2196_2197_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(counter[1]), 
            .I3(n38361), .O(n25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_3 (.CI(n38361), .I0(GND_net), .I1(counter[1]), 
            .CO(n38362));
    SB_LUT4 counter_2196_2197_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(counter[0]), 
            .I3(VCC_net), .O(n25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter_2196_2197_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter_2196_2197_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter[0]), 
            .CO(n38361));
    SB_LUT4 delay_counter_2194_2195_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[13]), .I3(n38360), .O(n61[13])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_2194_2195_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[12]), .I3(n38359), .O(n61[12])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_14 (.CI(n38359), .I0(GND_net), 
            .I1(delay_counter[12]), .CO(n38360));
    SB_LUT4 delay_counter_2194_2195_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n38358), .O(n61[11])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_13 (.CI(n38358), .I0(GND_net), 
            .I1(delay_counter[11]), .CO(n38359));
    SB_LUT4 delay_counter_2194_2195_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n38357), .O(n61[10])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_12 (.CI(n38357), .I0(GND_net), 
            .I1(delay_counter[10]), .CO(n38358));
    SB_LUT4 delay_counter_2194_2195_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n38356), .O(n61[9])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_11 (.CI(n38356), .I0(GND_net), 
            .I1(delay_counter[9]), .CO(n38357));
    SB_LUT4 delay_counter_2194_2195_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n38355), .O(n61[8])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_10 (.CI(n38355), .I0(GND_net), 
            .I1(delay_counter[8]), .CO(n38356));
    SB_LUT4 delay_counter_2194_2195_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n38354), .O(n61[7])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_9 (.CI(n38354), .I0(GND_net), 
            .I1(delay_counter[7]), .CO(n38355));
    SB_LUT4 delay_counter_2194_2195_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n38353), .O(n61[6])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_8 (.CI(n38353), .I0(GND_net), 
            .I1(delay_counter[6]), .CO(n38354));
    SB_LUT4 delay_counter_2194_2195_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n38352), .O(n61[5])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_7 (.CI(n38352), .I0(GND_net), 
            .I1(delay_counter[5]), .CO(n38353));
    SB_LUT4 delay_counter_2194_2195_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n38351), .O(n61[4])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_6 (.CI(n38351), .I0(GND_net), 
            .I1(delay_counter[4]), .CO(n38352));
    SB_LUT4 delay_counter_2194_2195_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n38350), .O(n61[3])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_5 (.CI(n38350), .I0(GND_net), 
            .I1(delay_counter[3]), .CO(n38351));
    SB_LUT4 delay_counter_2194_2195_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n38349), .O(n61[2])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_4 (.CI(n38349), .I0(GND_net), 
            .I1(delay_counter[2]), .CO(n38350));
    SB_LUT4 delay_counter_2194_2195_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n38348), .O(n61[1])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_3 (.CI(n38348), .I0(GND_net), 
            .I1(delay_counter[1]), .CO(n38349));
    SB_LUT4 delay_counter_2194_2195_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n61[0])) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_2194_2195_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_2194_2195_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(delay_counter[0]), .CO(n38348));
    SB_LUT4 i9860_3_lut (.I0(state[0]), .I1(n46880), .I2(state[1]), .I3(GND_net), 
            .O(n23333));   // verilog/tli4970.v(53[24:39])
    defparam i9860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 bit_counter_2192_add_4_9_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[7]), 
            .I3(n38316), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 bit_counter_2192_add_4_8_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[6]), 
            .I3(n38315), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2192_add_4_8 (.CI(n38315), .I0(VCC_net), .I1(bit_counter[6]), 
            .CO(n38316));
    SB_LUT4 bit_counter_2192_add_4_7_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[5]), 
            .I3(n38314), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2192_add_4_7 (.CI(n38314), .I0(VCC_net), .I1(bit_counter[5]), 
            .CO(n38315));
    SB_LUT4 bit_counter_2192_add_4_6_lut (.I0(GND_net), .I1(VCC_net), .I2(bit_counter[4]), 
            .I3(n38313), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY bit_counter_2192_add_4_6 (.CI(n38313), .I0(VCC_net), .I1(bit_counter[4]), 
            .CO(n38314));
    SB_LUT4 bit_counter_2192_add_4_5_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[3]), 
            .I3(n38312), .O(n46832)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_5 (.CI(n38312), .I0(VCC_net), .I1(bit_counter[3]), 
            .CO(n38313));
    SB_LUT4 bit_counter_2192_add_4_4_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[2]), 
            .I3(n38311), .O(n46831)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_4 (.CI(n38311), .I0(VCC_net), .I1(bit_counter[2]), 
            .CO(n38312));
    SB_LUT4 bit_counter_2192_add_4_3_lut (.I0(n1), .I1(VCC_net), .I2(bit_counter[1]), 
            .I3(n38310), .O(n46830)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_3 (.CI(n38310), .I0(VCC_net), .I1(bit_counter[1]), 
            .CO(n38311));
    SB_LUT4 bit_counter_2192_add_4_2_lut (.I0(n1), .I1(GND_net), .I2(bit_counter[0]), 
            .I3(VCC_net), .O(n46880)) /* synthesis syn_instantiated=1 */ ;
    defparam bit_counter_2192_add_4_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY bit_counter_2192_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(bit_counter[0]), 
            .CO(n38310));
    SB_DFFNESS state_i0 (.Q(state[0]), .C(clk_slow), .E(n27869), .D(n33707), 
            .S(n27983));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFSR counter_2196_2197__i5 (.Q(counter[4]), .C(CLK_c), .D(n25[4]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2196_2197__i4 (.Q(counter[3]), .C(CLK_c), .D(n25[3]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2196_2197__i3 (.Q(counter[2]), .C(CLK_c), .D(n25[2]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFSR counter_2196_2197__i2 (.Q(counter[1]), .C(CLK_c), .D(n25[1]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFNSR delay_counter_2194_2195__i14 (.Q(delay_counter[13]), .C(clk_slow), 
            .D(n61[13]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i13 (.Q(delay_counter[12]), .C(clk_slow), 
            .D(n61[12]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i12 (.Q(delay_counter[11]), .C(clk_slow), 
            .D(n61[11]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i11 (.Q(delay_counter[10]), .C(clk_slow), 
            .D(n61[10]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i10 (.Q(delay_counter[9]), .C(clk_slow), 
            .D(n61[9]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i9 (.Q(delay_counter[8]), .C(clk_slow), 
            .D(n61[8]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i8 (.Q(delay_counter[7]), .C(clk_slow), 
            .D(n61[7]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i7 (.Q(delay_counter[6]), .C(clk_slow), 
            .D(n61[6]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i6 (.Q(delay_counter[5]), .C(clk_slow), 
            .D(n61[5]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i5 (.Q(delay_counter[4]), .C(clk_slow), 
            .D(n61[4]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i4 (.Q(delay_counter[3]), .C(clk_slow), 
            .D(n61[3]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i3 (.Q(delay_counter[2]), .C(clk_slow), 
            .D(n61[2]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNSR delay_counter_2194_2195__i2 (.Q(delay_counter[1]), .C(clk_slow), 
            .D(n61[1]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFNE bit_counter_2192__i3 (.Q(bit_counter[3]), .C(clk_slow), .E(n27779), 
            .D(n23302));   // verilog/tli4970.v(53[24:39])
    SB_DFFNE bit_counter_2192__i2 (.Q(bit_counter[2]), .C(clk_slow), .E(n27779), 
            .D(n23304));   // verilog/tli4970.v(53[24:39])
    SB_DFFNE bit_counter_2192__i1 (.Q(bit_counter[1]), .C(clk_slow), .E(n27779), 
            .D(n23306));   // verilog/tli4970.v(53[24:39])
    SB_LUT4 i2_3_lut (.I0(\data[15] ), .I1(state[1]), .I2(state[0]), .I3(GND_net), 
            .O(n43722));
    defparam i2_3_lut.LUT_INIT = 16'hbfbf;
    SB_DFFN clk_out_66 (.Q(clk_out), .C(clk_slow), .D(n9_c));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN slave_select_65 (.Q(CS_c), .C(clk_slow), .D(n28230));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i0 (.Q(current[0]), .C(clk_slow), .D(n28227));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i1 (.Q(current[1]), .C(clk_slow), .D(n28692));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i2 (.Q(current[2]), .C(clk_slow), .D(n28691));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i3 (.Q(current[3]), .C(clk_slow), .D(n28690));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i4 (.Q(current[4]), .C(clk_slow), .D(n28689));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i5 (.Q(current[5]), .C(clk_slow), .D(n28688));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNE bit_counter_2192__i0 (.Q(bit_counter[0]), .C(clk_slow), .E(n27779), 
            .D(n23333));   // verilog/tli4970.v(53[24:39])
    SB_DFFN current_i0_i6 (.Q(current[6]), .C(clk_slow), .D(n28687));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i7 (.Q(current[7]), .C(clk_slow), .D(n28686));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFNSR delay_counter_2194_2195__i1 (.Q(delay_counter[0]), .C(clk_slow), 
            .D(n61[0]), .R(delay_counter_15__N_4288));   // verilog/tli4970.v(38[24:39])
    SB_DFFN current_i0_i8 (.Q(current[8]), .C(clk_slow), .D(n28685));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFSR counter_2196_2197__i1 (.Q(counter[0]), .C(CLK_c), .D(n25[0]), 
            .R(clk_slow_N_4207));   // verilog/tli4970.v(14[16:27])
    SB_DFFN current_i0_i9 (.Q(current[9]), .C(clk_slow), .D(n28684));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i10 (.Q(current[10]), .C(clk_slow), .D(n28683));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i11 (.Q(current[11]), .C(clk_slow), .D(n28682));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN current_i0_i12 (.Q(current[12]), .C(clk_slow), .D(n28681));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i15 (.Q(\data[15] ), .C(clk_slow), .D(n28185));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i12 (.Q(\data[12] ), .C(clk_slow), .D(n28184));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i11 (.Q(\data[11] ), .C(clk_slow), .D(n28183));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i10 (.Q(\data[10] ), .C(clk_slow), .D(n28182));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i9 (.Q(\data[9] ), .C(clk_slow), .D(n28181));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i8 (.Q(\data[8] ), .C(clk_slow), .D(n28180));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i7 (.Q(\data[7] ), .C(clk_slow), .D(n28179));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i6 (.Q(\data[6] ), .C(clk_slow), .D(n28178));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i5 (.Q(\data[5] ), .C(clk_slow), .D(n28177));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i4 (.Q(\data[4] ), .C(clk_slow), .D(n28176));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i3 (.Q(\data[3] ), .C(clk_slow), .D(n28175));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i2 (.Q(\data[2] ), .C(clk_slow), .D(n28174));   // verilog/tli4970.v(33[10] 66[6])
    SB_DFFN data_i1 (.Q(\data[1] ), .C(clk_slow), .D(n28173));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 i9833_3_lut (.I0(state[0]), .I1(n46830), .I2(state[1]), .I3(GND_net), 
            .O(n23306));   // verilog/tli4970.v(53[24:39])
    defparam i9833_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9831_3_lut (.I0(state[0]), .I1(n46831), .I2(state[1]), .I3(GND_net), 
            .O(n23304));   // verilog/tli4970.v(53[24:39])
    defparam i9831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9829_3_lut (.I0(state[0]), .I1(n46832), .I2(state[1]), .I3(GND_net), 
            .O(n23302));   // verilog/tli4970.v(53[24:39])
    defparam i9829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32803_2_lut (.I0(n15), .I1(state[0]), .I2(GND_net), .I3(GND_net), 
            .O(n33707));
    defparam i32803_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_76_i9_2_lut (.I0(state[0]), .I1(state[1]), .I2(GND_net), 
            .I3(GND_net), .O(state_7__N_4293));   // verilog/tli4970.v(51[7:17])
    defparam state_7__I_0_76_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i14396_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27779));
    defparam i14396_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i14716_3_lut_3_lut (.I0(state[0]), .I1(state[1]), .I2(CS_c), 
            .I3(GND_net), .O(n28230));   // verilog/tli4970.v(41[5] 65[12])
    defparam i14716_3_lut_3_lut.LUT_INIT = 16'hd1d1;
    SB_LUT4 i33428_4_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(clk_out), 
            .I3(n15), .O(n9_c));   // verilog/tli4970.v(41[5] 65[12])
    defparam i33428_4_lut_4_lut.LUT_INIT = 16'hf2b2;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15), .I1(state[1]), .I2(state[0]), .I3(delay_counter_15__N_4288), 
            .O(n27869));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfff4;
    SB_LUT4 i14469_2_lut_4_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(delay_counter_15__N_4288), .O(n27983));
    defparam i14469_2_lut_4_lut.LUT_INIT = 16'h0b00;
    SB_DFFN data_i0 (.Q(\data[0] ), .C(clk_slow), .D(n28458));   // verilog/tli4970.v(33[10] 66[6])
    SB_LUT4 equal_257_i9_2_lut (.I0(bit_counter[0]), .I1(bit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/tli4970.v(54[12:26])
    defparam equal_257_i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(bit_counter[5]), .I1(bit_counter[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4693));   // verilog/tli4970.v(54[12:26])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut (.I0(bit_counter[6]), .I1(bit_counter[7]), .I2(n11), 
            .I3(n6_adj_4693), .O(n15));   // verilog/tli4970.v(54[12:26])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1532 (.I0(delay_counter[5]), .I1(delay_counter[6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4694));
    defparam i2_2_lut_adj_1532.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(delay_counter[0]), .I1(delay_counter[1]), .I2(delay_counter[3]), 
            .I3(delay_counter[2]), .O(n43806));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1533 (.I0(n43806), .I1(n6_adj_4694), .I2(delay_counter[7]), 
            .I3(delay_counter[4]), .O(n43723));
    defparam i3_4_lut_adj_1533.LUT_INIT = 16'hfefc;
    SB_LUT4 i3_4_lut_adj_1534 (.I0(n43723), .I1(delay_counter[8]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n44313));
    defparam i3_4_lut_adj_1534.LUT_INIT = 16'h8000;
    SB_LUT4 i2303_4_lut (.I0(n44313), .I1(delay_counter[13]), .I2(delay_counter[12]), 
            .I3(delay_counter[11]), .O(delay_counter_15__N_4288));
    defparam i2303_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 mux_2295_i2_3_lut (.I0(n15), .I1(state[1]), .I2(state[0]), 
            .I3(GND_net), .O(n10078));
    defparam mux_2295_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(state[0]), .I1(state[1]), .I2(bit_counter[2]), 
            .I3(bit_counter[3]), .O(n26432));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1535 (.I0(state[0]), .I1(state[1]), 
            .I2(bit_counter[2]), .I3(bit_counter[3]), .O(n26440));   // verilog/tli4970.v(41[5] 65[12])
    defparam i1_2_lut_3_lut_4_lut_adj_1535.LUT_INIT = 16'hffbf;
    SB_LUT4 equal_257_i11_2_lut_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(bit_counter[0]), .I3(bit_counter[1]), .O(n11));   // verilog/tli4970.v(54[12:26])
    defparam equal_257_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1536 (.I0(bit_counter[2]), .I1(bit_counter[3]), 
            .I2(state[0]), .I3(state[1]), .O(n26445));   // verilog/tli4970.v(54[12:26])
    defparam i1_2_lut_3_lut_4_lut_adj_1536.LUT_INIT = 16'hfeff;
    SB_LUT4 i14522_2_lut_2_lut (.I0(state[1]), .I1(state[0]), .I2(GND_net), 
            .I3(GND_net), .O(n28035));   // verilog/tli4970.v(53[24:39])
    defparam i14522_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4796_1_lut (.I0(state[0]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));   // verilog/tli4970.v(41[5] 65[12])
    defparam i4796_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(bit_counter[2]), .I1(bit_counter[3]), .I2(state[0]), 
            .I3(state[1]), .O(n26435));   // verilog/tli4970.v(41[5] 65[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfbff;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (b_prev, a_new, encoder0_position, 
            GND_net, ENCODER0_B_N_keep, n1668, ENCODER0_A_N_keep, VCC_net, 
            direction_N_3907, n28461, n1632) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    output [1:0]a_new;
    output [31:0]encoder0_position;
    input GND_net;
    input ENCODER0_B_N_keep;
    input n1668;
    input ENCODER0_A_N_keep;
    input VCC_net;
    output direction_N_3907;
    input n28461;
    output n1632;
    
    
    wire debounce_cnt, a_prev_N_3913;
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire n28460, a_prev, n28459;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [31:0]n133;
    
    wire direction_N_3906, n38410, n38409, n38408, n38407, n38406, 
        n38405, n38404, n38403, n38402, n38401, n38400, n38399, 
        n38398, n38397, n38396, n38395, n38394, n38393, n38392, 
        n38391, n38390, n38389, n38388, n38387, n38386, n38385, 
        n38384, n38383, n38382, n38381, n38380, direction_N_3910;
    
    SB_LUT4 i14946_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(b_new[1]), 
            .I3(b_prev), .O(n28460));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14946_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14945_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3913), .I2(a_new[1]), 
            .I3(a_prev), .O(n28459));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i14945_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i32714_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(57[8:58])
    defparam i32714_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 position_2202_add_4_33_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[31]), .I3(n38410), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_2202_add_4_32_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[30]), .I3(n38409), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_32 (.CI(n38409), .I0(direction_N_3906), 
            .I1(encoder0_position[30]), .CO(n38410));
    SB_LUT4 position_2202_add_4_31_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[29]), .I3(n38408), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_31 (.CI(n38408), .I0(direction_N_3906), 
            .I1(encoder0_position[29]), .CO(n38409));
    SB_LUT4 position_2202_add_4_30_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[28]), .I3(n38407), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_30 (.CI(n38407), .I0(direction_N_3906), 
            .I1(encoder0_position[28]), .CO(n38408));
    SB_LUT4 position_2202_add_4_29_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[27]), .I3(n38406), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_29 (.CI(n38406), .I0(direction_N_3906), 
            .I1(encoder0_position[27]), .CO(n38407));
    SB_LUT4 position_2202_add_4_28_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[26]), .I3(n38405), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_28 (.CI(n38405), .I0(direction_N_3906), 
            .I1(encoder0_position[26]), .CO(n38406));
    SB_LUT4 position_2202_add_4_27_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[25]), .I3(n38404), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_27 (.CI(n38404), .I0(direction_N_3906), 
            .I1(encoder0_position[25]), .CO(n38405));
    SB_LUT4 position_2202_add_4_26_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[24]), .I3(n38403), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_26 (.CI(n38403), .I0(direction_N_3906), 
            .I1(encoder0_position[24]), .CO(n38404));
    SB_LUT4 position_2202_add_4_25_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[23]), .I3(n38402), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_25 (.CI(n38402), .I0(direction_N_3906), 
            .I1(encoder0_position[23]), .CO(n38403));
    SB_LUT4 position_2202_add_4_24_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[22]), .I3(n38401), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_24 (.CI(n38401), .I0(direction_N_3906), 
            .I1(encoder0_position[22]), .CO(n38402));
    SB_LUT4 position_2202_add_4_23_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[21]), .I3(n38400), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_23 (.CI(n38400), .I0(direction_N_3906), 
            .I1(encoder0_position[21]), .CO(n38401));
    SB_LUT4 position_2202_add_4_22_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[20]), .I3(n38399), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_22 (.CI(n38399), .I0(direction_N_3906), 
            .I1(encoder0_position[20]), .CO(n38400));
    SB_LUT4 position_2202_add_4_21_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[19]), .I3(n38398), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_21 (.CI(n38398), .I0(direction_N_3906), 
            .I1(encoder0_position[19]), .CO(n38399));
    SB_LUT4 position_2202_add_4_20_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[18]), .I3(n38397), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_20 (.CI(n38397), .I0(direction_N_3906), 
            .I1(encoder0_position[18]), .CO(n38398));
    SB_LUT4 position_2202_add_4_19_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[17]), .I3(n38396), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_19 (.CI(n38396), .I0(direction_N_3906), 
            .I1(encoder0_position[17]), .CO(n38397));
    SB_LUT4 position_2202_add_4_18_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[16]), .I3(n38395), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_18 (.CI(n38395), .I0(direction_N_3906), 
            .I1(encoder0_position[16]), .CO(n38396));
    SB_LUT4 position_2202_add_4_17_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[15]), .I3(n38394), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_17 (.CI(n38394), .I0(direction_N_3906), 
            .I1(encoder0_position[15]), .CO(n38395));
    SB_LUT4 position_2202_add_4_16_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[14]), .I3(n38393), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_16 (.CI(n38393), .I0(direction_N_3906), 
            .I1(encoder0_position[14]), .CO(n38394));
    SB_LUT4 position_2202_add_4_15_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[13]), .I3(n38392), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_15 (.CI(n38392), .I0(direction_N_3906), 
            .I1(encoder0_position[13]), .CO(n38393));
    SB_LUT4 position_2202_add_4_14_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[12]), .I3(n38391), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_14 (.CI(n38391), .I0(direction_N_3906), 
            .I1(encoder0_position[12]), .CO(n38392));
    SB_LUT4 position_2202_add_4_13_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[11]), .I3(n38390), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_13 (.CI(n38390), .I0(direction_N_3906), 
            .I1(encoder0_position[11]), .CO(n38391));
    SB_LUT4 position_2202_add_4_12_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[10]), .I3(n38389), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_12 (.CI(n38389), .I0(direction_N_3906), 
            .I1(encoder0_position[10]), .CO(n38390));
    SB_LUT4 position_2202_add_4_11_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[9]), .I3(n38388), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_11 (.CI(n38388), .I0(direction_N_3906), 
            .I1(encoder0_position[9]), .CO(n38389));
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1668), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_2202_add_4_10_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[8]), .I3(n38387), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_10 (.CI(n38387), .I0(direction_N_3906), 
            .I1(encoder0_position[8]), .CO(n38388));
    SB_LUT4 position_2202_add_4_9_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[7]), .I3(n38386), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_9 (.CI(n38386), .I0(direction_N_3906), 
            .I1(encoder0_position[7]), .CO(n38387));
    SB_LUT4 position_2202_add_4_8_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[6]), .I3(n38385), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_8 (.CI(n38385), .I0(direction_N_3906), 
            .I1(encoder0_position[6]), .CO(n38386));
    SB_LUT4 position_2202_add_4_7_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[5]), .I3(n38384), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1668), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_CARRY position_2202_add_4_7 (.CI(n38384), .I0(direction_N_3906), 
            .I1(encoder0_position[5]), .CO(n38385));
    SB_LUT4 position_2202_add_4_6_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[4]), .I3(n38383), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_6 (.CI(n38383), .I0(direction_N_3906), 
            .I1(encoder0_position[4]), .CO(n38384));
    SB_LUT4 position_2202_add_4_5_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[3]), .I3(n38382), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_5 (.CI(n38382), .I0(direction_N_3906), 
            .I1(encoder0_position[3]), .CO(n38383));
    SB_LUT4 position_2202_add_4_4_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[2]), .I3(n38381), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_4 (.CI(n38381), .I0(direction_N_3906), 
            .I1(encoder0_position[2]), .CO(n38382));
    SB_LUT4 position_2202_add_4_3_lut (.I0(GND_net), .I1(direction_N_3906), 
            .I2(encoder0_position[1]), .I3(n38380), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_3 (.CI(n38380), .I0(direction_N_3906), 
            .I1(encoder0_position[1]), .CO(n38381));
    SB_LUT4 position_2202_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_2202_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_2202_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n38380));
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1668), .D(a_prev_N_3913));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_2202__i31 (.Q(encoder0_position[31]), .C(n1668), .E(direction_N_3907), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i30 (.Q(encoder0_position[30]), .C(n1668), .E(direction_N_3907), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i29 (.Q(encoder0_position[29]), .C(n1668), .E(direction_N_3907), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i28 (.Q(encoder0_position[28]), .C(n1668), .E(direction_N_3907), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i27 (.Q(encoder0_position[27]), .C(n1668), .E(direction_N_3907), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i26 (.Q(encoder0_position[26]), .C(n1668), .E(direction_N_3907), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i25 (.Q(encoder0_position[25]), .C(n1668), .E(direction_N_3907), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i24 (.Q(encoder0_position[24]), .C(n1668), .E(direction_N_3907), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i23 (.Q(encoder0_position[23]), .C(n1668), .E(direction_N_3907), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i22 (.Q(encoder0_position[22]), .C(n1668), .E(direction_N_3907), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i21 (.Q(encoder0_position[21]), .C(n1668), .E(direction_N_3907), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i20 (.Q(encoder0_position[20]), .C(n1668), .E(direction_N_3907), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i19 (.Q(encoder0_position[19]), .C(n1668), .E(direction_N_3907), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i18 (.Q(encoder0_position[18]), .C(n1668), .E(direction_N_3907), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i17 (.Q(encoder0_position[17]), .C(n1668), .E(direction_N_3907), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i16 (.Q(encoder0_position[16]), .C(n1668), .E(direction_N_3907), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i15 (.Q(encoder0_position[15]), .C(n1668), .E(direction_N_3907), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i14 (.Q(encoder0_position[14]), .C(n1668), .E(direction_N_3907), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i13 (.Q(encoder0_position[13]), .C(n1668), .E(direction_N_3907), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i12 (.Q(encoder0_position[12]), .C(n1668), .E(direction_N_3907), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i11 (.Q(encoder0_position[11]), .C(n1668), .E(direction_N_3907), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i10 (.Q(encoder0_position[10]), .C(n1668), .E(direction_N_3907), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i9 (.Q(encoder0_position[9]), .C(n1668), .E(direction_N_3907), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i8 (.Q(encoder0_position[8]), .C(n1668), .E(direction_N_3907), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i7 (.Q(encoder0_position[7]), .C(n1668), .E(direction_N_3907), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i6 (.Q(encoder0_position[6]), .C(n1668), .E(direction_N_3907), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i5 (.Q(encoder0_position[5]), .C(n1668), .E(direction_N_3907), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i4 (.Q(encoder0_position[4]), .C(n1668), .E(direction_N_3907), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i3 (.Q(encoder0_position[3]), .C(n1668), .E(direction_N_3907), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i2 (.Q(encoder0_position[2]), .C(n1668), .E(direction_N_3907), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i1 (.Q(encoder0_position[1]), .C(n1668), .E(direction_N_3907), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_2202__i0 (.Q(encoder0_position[0]), .C(n1668), .E(direction_N_3907), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1668), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1668), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3906));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3910));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3910), 
            .I3(a_new[1]), .O(direction_N_3907));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_DFF direction_57 (.Q(n1632), .C(n1668), .D(n28461));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1668), .D(n28460));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1668), .D(n28459));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (pwm_out, clk32MHz, GND_net, VCC_net, pwm_setpoint) /* synthesis syn_module_defined=1 */ ;
    output pwm_out;
    input clk32MHz;
    input GND_net;
    input VCC_net;
    input [23:0]pwm_setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire pwm_out_N_797;
    wire [23:0]n101;
    wire [23:0]pwm_counter;   // verilog/pwm.v(11[19:30])
    
    wire n38300, n38299, n38298, n38297, n38296, n38295, n38294, 
        n38293, n38292, n38291, n38290, n38289, n38288, n38287, 
        n38286, n38285, n38284, n38283, n38282, n38281, n38280, 
        n38279, n38278, pwm_counter_23__N_795, n44075, n18, n21, 
        n20, n24, n19, n47169, n6, n8, n47135, n16, n10, n47146, 
        n12, n41, n39, n45, n37, n43, n29, n31, n23, n25, 
        n35, n33, n11, n13, n15, n27, n9, n17, n19_adj_4688, 
        n21_adj_4689, n47159, n47152, n30, n47420, n47416, n47734, 
        n47580, n47760, n47652, n47653, n24_adj_4690, n47138, n47516, 
        n47291, n4, n47650, n47651, n47148, n47736, n47293, n47786, 
        n47787, n47783, n47140, n47694, n47299, n47748;
    
    SB_DFF pwm_out_12 (.Q(pwm_out), .C(clk32MHz), .D(pwm_out_N_797));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_2190_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n38300), .O(n101[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_2190_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n38299), .O(n101[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_24 (.CI(n38299), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n38300));
    SB_LUT4 pwm_counter_2190_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n38298), .O(n101[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_23 (.CI(n38298), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n38299));
    SB_LUT4 pwm_counter_2190_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n38297), .O(n101[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_22 (.CI(n38297), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n38298));
    SB_LUT4 pwm_counter_2190_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n38296), .O(n101[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_21 (.CI(n38296), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n38297));
    SB_LUT4 pwm_counter_2190_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n38295), .O(n101[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_20 (.CI(n38295), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n38296));
    SB_LUT4 pwm_counter_2190_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n38294), .O(n101[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_19 (.CI(n38294), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n38295));
    SB_LUT4 pwm_counter_2190_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n38293), .O(n101[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_18 (.CI(n38293), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n38294));
    SB_LUT4 pwm_counter_2190_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n38292), .O(n101[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_17 (.CI(n38292), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n38293));
    SB_LUT4 pwm_counter_2190_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n38291), .O(n101[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_16 (.CI(n38291), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n38292));
    SB_LUT4 pwm_counter_2190_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n38290), .O(n101[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_15 (.CI(n38290), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n38291));
    SB_LUT4 pwm_counter_2190_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n38289), .O(n101[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_14 (.CI(n38289), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n38290));
    SB_LUT4 pwm_counter_2190_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n38288), .O(n101[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_13 (.CI(n38288), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n38289));
    SB_LUT4 pwm_counter_2190_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n38287), .O(n101[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_12 (.CI(n38287), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n38288));
    SB_LUT4 pwm_counter_2190_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n38286), .O(n101[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_11 (.CI(n38286), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n38287));
    SB_LUT4 pwm_counter_2190_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n38285), .O(n101[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_10 (.CI(n38285), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n38286));
    SB_LUT4 pwm_counter_2190_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n38284), .O(n101[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_9 (.CI(n38284), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n38285));
    SB_LUT4 pwm_counter_2190_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n38283), .O(n101[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_8 (.CI(n38283), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n38284));
    SB_LUT4 pwm_counter_2190_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n38282), .O(n101[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_7 (.CI(n38282), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n38283));
    SB_LUT4 pwm_counter_2190_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n38281), .O(n101[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_6 (.CI(n38281), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n38282));
    SB_LUT4 pwm_counter_2190_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n38280), .O(n101[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_5 (.CI(n38280), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n38281));
    SB_LUT4 pwm_counter_2190_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n38279), .O(n101[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_4 (.CI(n38279), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n38280));
    SB_LUT4 pwm_counter_2190_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n38278), .O(n101[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_3 (.CI(n38278), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n38279));
    SB_LUT4 pwm_counter_2190_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n101[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_2190_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_2190_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n38278));
    SB_DFFSR pwm_counter_2190__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n101[23]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n101[22]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n101[21]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n101[20]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n101[19]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n101[18]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n101[17]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n101[16]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n101[15]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n101[14]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n101[13]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n101[12]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n101[11]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n101[10]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n101[9]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n101[8]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n101[7]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n101[6]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n101[5]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n101[4]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n101[3]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n101[2]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n101[1]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_2190__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n101[0]), 
            .R(pwm_counter_23__N_795));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n44075));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut (.I0(pwm_counter[19]), .I1(n44075), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n18));
    defparam i5_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i8_4_lut (.I0(pwm_counter[22]), .I1(pwm_counter[14]), .I2(pwm_counter[15]), 
            .I3(pwm_counter[17]), .O(n21));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(pwm_counter[20]), .I1(pwm_counter[21]), .I2(pwm_counter[11]), 
            .I3(GND_net), .O(n20));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n21), .I1(pwm_counter[18]), .I2(n18), .I3(pwm_counter[16]), 
            .O(n24));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(pwm_counter[13]), .I1(pwm_counter[12]), .I2(GND_net), 
            .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33433_4_lut (.I0(pwm_counter[23]), .I1(n19), .I2(n24), .I3(n20), 
            .O(pwm_counter_23__N_795));   // verilog/pwm.v(18[8:40])
    defparam i33433_4_lut.LUT_INIT = 16'h5554;
    SB_LUT4 i32038_3_lut_4_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(pwm_counter[2]), .O(n47169));   // verilog/pwm.v(21[8:24])
    defparam i32038_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(pwm_setpoint[2]), .I3(GND_net), .O(n6));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32004_2_lut_4_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[9]), .I3(pwm_setpoint[9]), .O(n47135));
    defparam i32004_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(pwm_setpoint[9]), .I1(pwm_setpoint[21]), 
            .I2(pwm_counter[21]), .I3(GND_net), .O(n16));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i32015_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n47146));
    defparam i32015_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(pwm_counter[20]), .I1(pwm_setpoint[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(pwm_counter[19]), .I1(pwm_setpoint[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(pwm_counter[22]), .I1(pwm_setpoint[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(pwm_counter[18]), .I1(pwm_setpoint[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(pwm_counter[21]), .I1(pwm_setpoint[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4688));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4689));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i32028_4_lut (.I0(n21_adj_4689), .I1(n19_adj_4688), .I2(n17), 
            .I3(n9), .O(n47159));
    defparam i32028_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32021_4_lut (.I0(n27), .I1(n15), .I2(n13), .I3(n11), .O(n47152));
    defparam i32021_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12), .I1(pwm_setpoint[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32288_4_lut (.I0(n13), .I1(n11), .I2(n9), .I3(n47169), 
            .O(n47420));
    defparam i32288_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32284_4_lut (.I0(n19_adj_4688), .I1(n17), .I2(n15), .I3(n47420), 
            .O(n47416));
    defparam i32284_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i32602_4_lut (.I0(n25), .I1(n23), .I2(n21_adj_4689), .I3(n47416), 
            .O(n47734));
    defparam i32602_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32448_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n47734), 
            .O(n47580));
    defparam i32448_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i32628_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n47580), 
            .O(n47760));
    defparam i32628_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i32520_3_lut (.I0(n6), .I1(pwm_setpoint[10]), .I2(n21_adj_4689), 
            .I3(GND_net), .O(n47652));   // verilog/pwm.v(21[8:24])
    defparam i32520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32521_3_lut (.I0(n47652), .I1(pwm_setpoint[11]), .I2(n23), 
            .I3(GND_net), .O(n47653));   // verilog/pwm.v(21[8:24])
    defparam i32521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16), .I1(pwm_setpoint[22]), .I2(n45), 
            .I3(GND_net), .O(n24_adj_4690));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32007_4_lut (.I0(n43), .I1(n25), .I2(n23), .I3(n47159), 
            .O(n47138));
    defparam i32007_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32384_4_lut (.I0(n24_adj_4690), .I1(n8), .I2(n45), .I3(n47135), 
            .O(n47516));   // verilog/pwm.v(21[8:24])
    defparam i32384_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32159_3_lut (.I0(n47653), .I1(pwm_setpoint[12]), .I2(n25), 
            .I3(GND_net), .O(n47291));   // verilog/pwm.v(21[8:24])
    defparam i32159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4));   // verilog/pwm.v(21[8:24])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i32518_3_lut (.I0(n4), .I1(pwm_setpoint[13]), .I2(n27), .I3(GND_net), 
            .O(n47650));   // verilog/pwm.v(21[8:24])
    defparam i32518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32519_3_lut (.I0(n47650), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n47651));   // verilog/pwm.v(21[8:24])
    defparam i32519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32017_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n47152), 
            .O(n47148));
    defparam i32017_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32604_4_lut (.I0(n30), .I1(n10), .I2(n35), .I3(n47146), 
            .O(n47736));   // verilog/pwm.v(21[8:24])
    defparam i32604_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i32161_3_lut (.I0(n47651), .I1(pwm_setpoint[15]), .I2(n31), 
            .I3(GND_net), .O(n47293));   // verilog/pwm.v(21[8:24])
    defparam i32161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32654_4_lut (.I0(n47293), .I1(n47736), .I2(n35), .I3(n47148), 
            .O(n47786));   // verilog/pwm.v(21[8:24])
    defparam i32654_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32655_3_lut (.I0(n47786), .I1(pwm_setpoint[18]), .I2(n37), 
            .I3(GND_net), .O(n47787));   // verilog/pwm.v(21[8:24])
    defparam i32655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32651_3_lut (.I0(n47787), .I1(pwm_setpoint[19]), .I2(n39), 
            .I3(GND_net), .O(n47783));   // verilog/pwm.v(21[8:24])
    defparam i32651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32009_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n47760), 
            .O(n47140));
    defparam i32009_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i32562_4_lut (.I0(n47291), .I1(n47516), .I2(n45), .I3(n47138), 
            .O(n47694));   // verilog/pwm.v(21[8:24])
    defparam i32562_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32167_3_lut (.I0(n47783), .I1(pwm_setpoint[20]), .I2(n41), 
            .I3(GND_net), .O(n47299));   // verilog/pwm.v(21[8:24])
    defparam i32167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i32616_4_lut (.I0(n47299), .I1(n47694), .I2(n45), .I3(n47140), 
            .O(n47748));   // verilog/pwm.v(21[8:24])
    defparam i32616_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i32617_3_lut (.I0(n47748), .I1(pwm_counter[23]), .I2(pwm_setpoint[23]), 
            .I3(GND_net), .O(pwm_out_N_797));   // verilog/pwm.v(21[8:24])
    defparam i32617_3_lut.LUT_INIT = 16'h8e8e;
    
endmodule
//
// Verilog Description of module coms
//

module coms (n28303, \data_out_frame[18] , CLK_c, \data_out_frame[20] , 
            GND_net, n28302, \data_out_frame[19] , n28301, n28300, 
            n28299, n28298, n28297, n28296, \data_out_frame[25] , 
            \data_out_frame[14] , n27647, \data_out_frame[16] , \data_out_frame[15] , 
            n40583, n28295, n28294, n28293, n28292, \data_out_frame[10] , 
            \data_out_frame[6] , \data_out_frame[5] , \data_out_frame[9] , 
            \data_out_frame[8] , \data_out_frame[11] , \data_out_frame[13] , 
            \data_out_frame[12] , \data_out_frame[4] , \data_out_frame[22] , 
            \data_out_frame[23] , \data_out_frame[24] , \data_out_frame[21][2] , 
            \data_out_frame[7] , \FRAME_MATCHER.state , n28291, \data_out_frame[17] , 
            \data_out_frame[21][1] , n28290, \data_in_frame[14] , \data_in_frame[19] , 
            \data_in_frame[11] , \data_in_frame[15] , \data_in_frame[12] , 
            \data_in_frame[2] , \data_in_frame[9] , \data_in_frame[13] , 
            \data_in_frame[10] , \data_in_frame[3] , \data_in_frame[7] , 
            \data_in_frame[5] , \data_in_frame[6] , \data_in_frame[1] , 
            n28289, \data_in_frame[8] , n27617, rx_data, \data_in_frame[4] , 
            \data_in_frame[21] , \r_SM_Main_2__N_3616[0] , \data_out_frame[21][0] , 
            rx_data_ready, setpoint, \data_out_frame[21][3] , n28288, 
            n28287, n28286, n28285, n28284, n28283, n28282, \data_out_frame[21][4] , 
            n28281, n28280, n28279, n28278, n28277, n28276, n28275, 
            n28274, n28273, \Kp[13] , n42276, n42287, n42266, n28272, 
            n28271, \Ki[11] , DE_c, n28270, \Kp[12] , n28269, \Ki[12] , 
            n28268, \Ki[13] , n28267, \Ki[14] , n28266, n28265, 
            \Kp[11] , n28264, \Ki[15] , n28263, n28262, n28261, 
            n28260, n28259, n28258, n28257, n28256, n28255, n28254, 
            n28253, \data_out_frame[27][0] , n28252, ID, n122, \FRAME_MATCHER.state_31__N_2660[2] , 
            n26494, n4452, n7, n3303, \FRAME_MATCHER.state_31__N_2788[2] , 
            n28251, n28783, neopxl_color, n28782, n28781, n28780, 
            n28779, n28778, n28777, n28776, n28775, n28774, n28773, 
            n28772, n28771, n28770, n28250, n28249, n28248, n28247, 
            n28246, n28245, n28244, n28243, \Kp[14] , n28242, n28241, 
            \data_in[2] , n28240, n28239, n28238, n28237, n28236, 
            n28234, \Kp[10] , n28233, \Kp[9] , n28232, n28226, \Kp[8] , 
            n28225, \Kp[7] , n28224, \Kp[6] , n28223, \Kp[5] , n28222, 
            \Kp[4] , n28221, n41665, n28219, PWMLimit, n28218, \data_in[3] , 
            LED_c, n28217, control_mode, n28215, n28214, \Kp[3] , 
            n28213, \Ki[0] , n28212, \Kp[0] , n28211, \data_in[0] , 
            n28210, \Kp[2] , n28209, \Kp[1] , n28208, n28207, n28206, 
            n28205, n28204, n28202, n28746, n28745, n28744, n28743, 
            n28742, n28741, n28740, n28739, n28730, n28729, n28728, 
            n28727, n28726, n28725, n28724, n28723, n28714, n28713, 
            n28712, n28711, n28710, n28709, n28708, n28707, n28169, 
            n28168, IntegralLimit, n28166, n28164, n28163, n28162, 
            n28161, n28160, n19799, n34010, n23516, n28159, n28158, 
            \data_in[1] , n23622, n42267, n42288, n28669, n28157, 
            n28668, n28667, n28666, n28665, n42244, n43094, n26482, 
            n62, n28664, n28663, n28662, n19, n28652, n28651, 
            n28650, n28618, n28617, n28616, n28615, n28612, n28604, 
            n28603, n28602, n28601, n28600, n28599, n28598, n28597, 
            n28596, n28595, n28594, n28593, n28592, n28591, n28590, 
            n28589, n28588, n28587, n28586, n28585, n28584, n28583, 
            n28582, n28581, n28580, n28579, n28578, n28577, n28576, 
            n28575, n28574, n28573, n28572, n28571, n20, n28546, 
            n28545, n28544, n28543, n28542, n28541, n28540, n28539, 
            n28530, n28529, n28528, n28527, n28526, n28525, n28524, 
            n28523, n28522, n28521, n28520, n28519, n28518, n28517, 
            n28516, n28515, n28514, n28510, n28509, n28508, n28507, 
            n28506, n28505, n28501, n28500, n28499, n28498, n28497, 
            n28496, n28495, n28494, n28493, n28492, n28491, n28490, 
            n28489, n28488, n28487, n28483, n28482, n28479, n28478, 
            n28477, n28476, n28475, n28474, n28473, n28472, n28471, 
            n48873, n28469, n28468, n28467, n28466, n28465, n28464, 
            n28463, n28462, n28457, n28456, n28455, n28454, n28453, 
            n28452, n28451, n28450, n28449, n28448, n28447, n28446, 
            n28445, n28444, n28443, n28442, n28441, n28440, n28439, 
            n28438, n28433, n28432, n28428, n28426, \Ki[1] , n28425, 
            n28424, \Ki[2] , n28423, n28422, n28421, n28420, n28419, 
            n28418, n28417, n28416, n28415, n28414, n28413, n28412, 
            n28411, n28410, n28409, n28408, n28407, n28406, n28405, 
            n28404, n28403, n28402, n28401, n28400, n28399, n28398, 
            n28397, n28396, n28395, n28394, n28393, n28392, n28391, 
            n28390, n28389, n28384, n28383, \Ki[3] , n28382, \Ki[4] , 
            n28381, n28380, n28379, \Ki[5] , n28378, n28377, n28376, 
            n28375, n28374, n28373, n28372, n28371, n28370, n28369, 
            n28368, n28367, n28366, n28365, n28364, n28363, n28362, 
            n28361, n28360, n28359, n28358, n28357, n28356, n28355, 
            n28354, n28353, n28352, n28351, n28350, n28349, n28348, 
            n28347, n28346, n28345, n28344, n28343, n28342, n28341, 
            n28340, n28335, n28331, n28329, n28328, n28327, n28326, 
            n28325, n28324, n28323, n28322, n28321, n28320, n28319, 
            \Ki[6] , n28317, n28316, n28314, \Kp[15] , n28313, n28312, 
            n28311, \Ki[7] , n28310, \Ki[8] , n28309, \Ki[9] , n28308, 
            n28156, n28307, \Ki[10] , n28306, n28305, n28304, n60, 
            n6, tx_active, \state[0] , \state[2] , \state[3] , n7233, 
            n43068, n42251, n42255, n42299, n32652, n42277, n42264, 
            n42285, n44019, \r_Bit_Index[0] , n27840, r_SM_Main, n28123, 
            \r_SM_Main_2__N_3613[1] , tx_o, VCC_net, n28387, n28235, 
            n18934, n4, n48874, tx_enable, \r_Bit_Index[0]_adj_3 , 
            n27844, r_SM_Main_adj_10, n28125, \r_SM_Main_2__N_3542[2] , 
            r_Rx_Data, RX_N_10, n4_adj_7, n4_adj_8, n4_adj_9, n26398, 
            n26390, n33332, n28431, n41875, n28203, n28201, n28200, 
            n28199, n28198, n28197, n28196, n42166, n28437) /* synthesis syn_module_defined=1 */ ;
    input n28303;
    output [7:0]\data_out_frame[18] ;
    input CLK_c;
    output [7:0]\data_out_frame[20] ;
    input GND_net;
    input n28302;
    output [7:0]\data_out_frame[19] ;
    input n28301;
    input n28300;
    input n28299;
    input n28298;
    input n28297;
    input n28296;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[14] ;
    output n27647;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[15] ;
    output n40583;
    input n28295;
    input n28294;
    input n28293;
    input n28292;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[22] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[24] ;
    output \data_out_frame[21][2] ;
    output [7:0]\data_out_frame[7] ;
    output [31:0]\FRAME_MATCHER.state ;
    input n28291;
    output [7:0]\data_out_frame[17] ;
    output \data_out_frame[21][1] ;
    input n28290;
    output [7:0]\data_in_frame[14] ;
    output [7:0]\data_in_frame[19] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[15] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[7] ;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[1] ;
    input n28289;
    output [7:0]\data_in_frame[8] ;
    output n27617;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[21] ;
    output \r_SM_Main_2__N_3616[0] ;
    output \data_out_frame[21][0] ;
    output rx_data_ready;
    output [23:0]setpoint;
    output \data_out_frame[21][3] ;
    input n28288;
    input n28287;
    input n28286;
    input n28285;
    input n28284;
    input n28283;
    input n28282;
    output \data_out_frame[21][4] ;
    input n28281;
    input n28280;
    input n28279;
    input n28278;
    input n28277;
    input n28276;
    input n28275;
    input n28274;
    input n28273;
    output \Kp[13] ;
    output n42276;
    output n42287;
    output n42266;
    input n28272;
    input n28271;
    output \Ki[11] ;
    output DE_c;
    input n28270;
    output \Kp[12] ;
    input n28269;
    output \Ki[12] ;
    input n28268;
    output \Ki[13] ;
    input n28267;
    output \Ki[14] ;
    input n28266;
    input n28265;
    output \Kp[11] ;
    input n28264;
    output \Ki[15] ;
    input n28263;
    input n28262;
    input n28261;
    input n28260;
    input n28259;
    input n28258;
    input n28257;
    input n28256;
    input n28255;
    input n28254;
    input n28253;
    output \data_out_frame[27][0] ;
    input n28252;
    input [7:0]ID;
    output n122;
    output \FRAME_MATCHER.state_31__N_2660[2] ;
    output n26494;
    output n4452;
    output n7;
    output n3303;
    output \FRAME_MATCHER.state_31__N_2788[2] ;
    input n28251;
    input n28783;
    output [23:0]neopxl_color;
    input n28782;
    input n28781;
    input n28780;
    input n28779;
    input n28778;
    input n28777;
    input n28776;
    input n28775;
    input n28774;
    input n28773;
    input n28772;
    input n28771;
    input n28770;
    input n28250;
    input n28249;
    input n28248;
    input n28247;
    input n28246;
    input n28245;
    input n28244;
    input n28243;
    output \Kp[14] ;
    input n28242;
    input n28241;
    output [7:0]\data_in[2] ;
    input n28240;
    input n28239;
    input n28238;
    input n28237;
    input n28236;
    input n28234;
    output \Kp[10] ;
    input n28233;
    output \Kp[9] ;
    input n28232;
    input n28226;
    output \Kp[8] ;
    input n28225;
    output \Kp[7] ;
    input n28224;
    output \Kp[6] ;
    input n28223;
    output \Kp[5] ;
    input n28222;
    output \Kp[4] ;
    input n28221;
    input n41665;
    input n28219;
    output [23:0]PWMLimit;
    input n28218;
    output [7:0]\data_in[3] ;
    output LED_c;
    input n28217;
    output [7:0]control_mode;
    input n28215;
    input n28214;
    output \Kp[3] ;
    input n28213;
    output \Ki[0] ;
    input n28212;
    output \Kp[0] ;
    input n28211;
    output [7:0]\data_in[0] ;
    input n28210;
    output \Kp[2] ;
    input n28209;
    output \Kp[1] ;
    input n28208;
    input n28207;
    input n28206;
    input n28205;
    input n28204;
    input n28202;
    input n28746;
    input n28745;
    input n28744;
    input n28743;
    input n28742;
    input n28741;
    input n28740;
    input n28739;
    input n28730;
    input n28729;
    input n28728;
    input n28727;
    input n28726;
    input n28725;
    input n28724;
    input n28723;
    input n28714;
    input n28713;
    input n28712;
    input n28711;
    input n28710;
    input n28709;
    input n28708;
    input n28707;
    input n28169;
    input n28168;
    output [23:0]IntegralLimit;
    input n28166;
    input n28164;
    input n28163;
    input n28162;
    input n28161;
    input n28160;
    output n19799;
    output n34010;
    output n23516;
    input n28159;
    input n28158;
    output [7:0]\data_in[1] ;
    output n23622;
    output n42267;
    output n42288;
    input n28669;
    input n28157;
    input n28668;
    input n28667;
    input n28666;
    input n28665;
    output n42244;
    input n43094;
    output n26482;
    output n62;
    input n28664;
    input n28663;
    input n28662;
    input n19;
    input n28652;
    input n28651;
    input n28650;
    input n28618;
    input n28617;
    input n28616;
    input n28615;
    input n28612;
    input n28604;
    input n28603;
    input n28602;
    input n28601;
    input n28600;
    input n28599;
    input n28598;
    input n28597;
    input n28596;
    input n28595;
    input n28594;
    input n28593;
    input n28592;
    input n28591;
    input n28590;
    input n28589;
    input n28588;
    input n28587;
    input n28586;
    input n28585;
    input n28584;
    input n28583;
    input n28582;
    input n28581;
    input n28580;
    input n28579;
    input n28578;
    input n28577;
    input n28576;
    input n28575;
    input n28574;
    input n28573;
    input n28572;
    input n28571;
    output n20;
    input n28546;
    input n28545;
    input n28544;
    input n28543;
    input n28542;
    input n28541;
    input n28540;
    input n28539;
    input n28530;
    input n28529;
    input n28528;
    input n28527;
    input n28526;
    input n28525;
    input n28524;
    input n28523;
    input n28522;
    input n28521;
    input n28520;
    input n28519;
    input n28518;
    input n28517;
    input n28516;
    input n28515;
    input n28514;
    input n28510;
    input n28509;
    input n28508;
    input n28507;
    input n28506;
    input n28505;
    input n28501;
    input n28500;
    input n28499;
    input n28498;
    input n28497;
    input n28496;
    input n28495;
    input n28494;
    input n28493;
    input n28492;
    input n28491;
    input n28490;
    input n28489;
    input n28488;
    input n28487;
    input n28483;
    input n28482;
    input n28479;
    input n28478;
    input n28477;
    input n28476;
    input n28475;
    input n28474;
    input n28473;
    input n28472;
    input n28471;
    input n48873;
    input n28469;
    input n28468;
    input n28467;
    input n28466;
    input n28465;
    input n28464;
    input n28463;
    input n28462;
    input n28457;
    input n28456;
    input n28455;
    input n28454;
    input n28453;
    input n28452;
    input n28451;
    input n28450;
    input n28449;
    input n28448;
    input n28447;
    input n28446;
    input n28445;
    input n28444;
    input n28443;
    input n28442;
    input n28441;
    input n28440;
    input n28439;
    input n28438;
    input n28433;
    input n28432;
    input n28428;
    input n28426;
    output \Ki[1] ;
    input n28425;
    input n28424;
    output \Ki[2] ;
    input n28423;
    input n28422;
    input n28421;
    input n28420;
    input n28419;
    input n28418;
    input n28417;
    input n28416;
    input n28415;
    input n28414;
    input n28413;
    input n28412;
    input n28411;
    input n28410;
    input n28409;
    input n28408;
    input n28407;
    input n28406;
    input n28405;
    input n28404;
    input n28403;
    input n28402;
    input n28401;
    input n28400;
    input n28399;
    input n28398;
    input n28397;
    input n28396;
    input n28395;
    input n28394;
    input n28393;
    input n28392;
    input n28391;
    input n28390;
    input n28389;
    input n28384;
    input n28383;
    output \Ki[3] ;
    input n28382;
    output \Ki[4] ;
    input n28381;
    input n28380;
    input n28379;
    output \Ki[5] ;
    input n28378;
    input n28377;
    input n28376;
    input n28375;
    input n28374;
    input n28373;
    input n28372;
    input n28371;
    input n28370;
    input n28369;
    input n28368;
    input n28367;
    input n28366;
    input n28365;
    input n28364;
    input n28363;
    input n28362;
    input n28361;
    input n28360;
    input n28359;
    input n28358;
    input n28357;
    input n28356;
    input n28355;
    input n28354;
    input n28353;
    input n28352;
    input n28351;
    input n28350;
    input n28349;
    input n28348;
    input n28347;
    input n28346;
    input n28345;
    input n28344;
    input n28343;
    input n28342;
    input n28341;
    input n28340;
    input n28335;
    input n28331;
    input n28329;
    input n28328;
    input n28327;
    input n28326;
    input n28325;
    input n28324;
    input n28323;
    input n28322;
    input n28321;
    input n28320;
    input n28319;
    output \Ki[6] ;
    input n28317;
    input n28316;
    input n28314;
    output \Kp[15] ;
    input n28313;
    input n28312;
    input n28311;
    output \Ki[7] ;
    input n28310;
    output \Ki[8] ;
    input n28309;
    output \Ki[9] ;
    input n28308;
    input n28156;
    input n28307;
    output \Ki[10] ;
    input n28306;
    input n28305;
    input n28304;
    output n60;
    output n6;
    output tx_active;
    input \state[0] ;
    input \state[2] ;
    input \state[3] ;
    output n7233;
    input n43068;
    output n42251;
    output n42255;
    output n42299;
    output n32652;
    output n42277;
    output n42264;
    output n42285;
    output n44019;
    output \r_Bit_Index[0] ;
    output n27840;
    output [2:0]r_SM_Main;
    output n28123;
    output \r_SM_Main_2__N_3613[1] ;
    output tx_o;
    input VCC_net;
    input n28387;
    input n28235;
    output n18934;
    output n4;
    input n48874;
    output tx_enable;
    output \r_Bit_Index[0]_adj_3 ;
    output n27844;
    output [2:0]r_SM_Main_adj_10;
    output n28125;
    output \r_SM_Main_2__N_3542[2] ;
    output r_Rx_Data;
    input RX_N_10;
    output n4_adj_7;
    output n4_adj_8;
    output n4_adj_9;
    output n26398;
    output n26390;
    output n33332;
    input n28431;
    input n41875;
    input n28203;
    input n28201;
    input n28200;
    input n28199;
    input n28198;
    input n28197;
    input n28196;
    input n42166;
    input n28437;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n42503, n39859;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3846, n3, n39586, n40632, n42655, n42687, n24648, n44126, 
        n4_c, n3_adj_4405, n44528;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n42923, n40485, n10, n42968, n40535, n42785, n40513, 
        n14, n39685, n27602, n26860, n3_adj_4406, n43493, n27027, 
        n42699, n42944, n14_adj_4407, n44255, n43687, n44708, n43608;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n27558, n26965, n27257, n42769, n9, n40489, n42477, n42702, 
        n42965, n10_adj_4408, n42367, n42788, n26722, n27309, n14_adj_4409, 
        n42838, n42564, n15, n27329, n26511, n27374, n27507, n10_adj_4410, 
        n39567, n26912, n42844, n42403;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n48832, n42905, n6_c, n42760, n42576, n40525, n42741, 
        n39574, n42348, n42313, n10_adj_4411, n26748, n42484, n3_adj_4412, 
        n3_adj_4413, n42529, n12, n26097, n42878, n39506, n42814, 
        n42385, n42452, n12_adj_4414, n1516, n42458, n26989, n3_adj_4415, 
        n3_adj_4416, n6_adj_4417, n27084, n3_adj_4418, n48808, n48811, 
        n3_adj_4419, n48850, n48853, n45861, n45862, n45860, n48583, 
        n48589, n14_adj_4420, n48793, n46849, n48757, n48835, n47458, 
        n45856, n45854, n48751, n48613, n14_adj_4421, n48799, n46834, 
        n42754, n6_adj_4422, n44033;
    wire [31:0]\FRAME_MATCHER.state_c ;   // verilog/coms.v(112[11:16])
    
    wire n23237, n3_adj_4423, n2134, n42417, n6_adj_4424, n43653, 
        n24129, n45899;
    wire [7:0]n8825;
    
    wire n27701, n28149, n45900, n3_adj_4425, n42613, n27282, n42850, 
        n10_adj_4426, n40529, n44014, n3_adj_4427, n45906, n26899, 
        n45905, n3_adj_4428, n3_adj_4429, n42309, n42696, n42413, 
        n42757, n45849, n45850, n3_adj_4430, n45848, n48697, n48649, 
        n14_adj_4431, n42521, n40487, n43490, n3_adj_4432, n42953, 
        n42884, n43563, n42887, n42799, n42956, n10_adj_4433, n3_adj_4434, 
        n3_adj_4435, n42649, n42868, n10_adj_4436;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n40264, n44109, n40531, n40474, n39500, n8, Kp_23__N_861, 
        n42573;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n6_adj_4437, n26617, n27095, n42607, n42881, n40630, n42720, 
        n6_adj_4438, n44174, n3_adj_4439, n42871, n42811, n40538, 
        n3_adj_4440, n42524, n39548, n42714, n26784, n42791, n42490, 
        n39908, n42558, n26938, n40613, n39836, n42584;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n26056, n42640, n39616, n14_adj_4441, n13;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n42744, n42587, n26025, n40559, n39793, n27215, n42630, 
        n42631, n42859, n27436, n39606, n10_adj_4442, n26646, n42841, 
        n42593, n12_adj_4443, n42708, n42590, n42890, n36, n42847, 
        n42468, n34, n26, n40, n38, n39, n42805, n42462, n42729, 
        n37, n26687, n27551, n6_adj_4444, n39554, n42682, n26581, 
        n27203, n27451, n24, n39321, n17, n13_adj_4445, n27199, 
        n27588, n22, n26_adj_4446, n42862, n11, n48805, n46829, 
        n48691, n47462, n16, n8_adj_4447, n17_adj_4448, n42551, 
        n40481, n10_adj_4449, n26756, n14_adj_4450, n27071, n40557, 
        n42950, n42829, n42646, n40499, n40457, n6_adj_4451, n42322, 
        n42826, n42832, n31, n31_adj_4452, n42248, n7_c, n42296, 
        n40521, n18, Kp_23__N_1306, n42500, Kp_23__N_1330, n20_c, 
        n15_adj_4453, n39918, n23788, n1, n39598, n26809, n6_adj_4454, 
        n42334, n32, n31_adj_4455, n27137, n35, n42471, n26801, 
        n34_adj_4456, n38_adj_4457, n27196, n42548, n33, n42865, 
        n36_adj_4458, n25, n34_adj_4459, n20_adj_4460, n23, n7001, 
        n40_adj_4461, n7003, n7004, n7005, n38_adj_4462, n7006, 
        n39_adj_4463, n42637, n42302, n37_adj_4464, n7007, n15_adj_4465, 
        n44139, n27234, n22_adj_4466, n26_adj_4467, n44102, n7008, 
        n7009, n7010, n7011, n26496, n40566, n42685, n42433, n7012, 
        n7013, n44477, n2, n3_adj_4468, n7014, n7015, n26789, 
        n40472, n7016, n28, n42561, n8_adj_4469, n42281, n28731, 
        n7017, n7018, n7019, n7020, n7021, n7022, n42775, n1519, 
        n26_adj_4470, n6_adj_4471, n7023, n26667, n24724, n12_adj_4472, 
        n7024, n40494, n10_adj_4473, n42920, n40492, n27, n7025, 
        n26633, n27407, n16_adj_4474, n42941, n17_adj_4475, n27104, 
        n42567, n12_adj_4476, n27227, n42835, n39631, n42370, n42555, 
        n12_adj_4477, n6_adj_4478, n27246, n42319, n5, n42962, n42328, 
        n42902, n15_adj_4479, n42389, n14_adj_4480, n26968, n42361, 
        n42938, n12_adj_4481, n16_adj_4482, n17_adj_4483, Kp_23__N_1214, 
        n42689, n1668, n25_adj_4484, n10_adj_4485, n39516, n5_adj_4486;
    wire [0:0]n4888;
    
    wire n43197, n6_adj_4487, n6_adj_4488, n8_adj_4489, n10_adj_4490, 
        \FRAME_MATCHER.rx_data_ready_prev , n43569, n42620, n7002, n27685;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n44433, n43617, n43671, n6_adj_4491, n43611, n40620, n8_adj_4492, 
        n39556, n43826, n44504, n44257, n44269, n43861, n12_adj_4493, 
        n43516, n4_adj_4494, n18_adj_4495, n11_adj_4496, n44400, n20_adj_4497, 
        n44600, n25_adj_4498, n8_adj_4499, n45678, n26527, n28732, 
        n3_adj_4500, n42738, n28733, n45680, n28734, n42395, n10_adj_4501, 
        n27_adj_4502, n28735, n29, n42305, n42817, n42732, n42533, 
        n3_adj_4503, n28736, n28737, n3_adj_4504, n45831, n48823, 
        n46815, n45990, n48844, n28738, n20_adj_4505, n42959, n42693, 
        n12_adj_4506, n45832, n45830, n48577, n48769, n14_adj_4507, 
        n48775, n45991, n45945, n7_adj_4508, n45944;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n48829, n46817, n45984, n42274, n20_adj_4509, n45826, n45824, 
        n42260, n48763, n48595, n14_adj_4510, n48745, n45985, n45816, 
        n7_adj_4511, n45815, n48571, n46819, n45981, n20_adj_4512, 
        n45820, n45818, n48733, n48607, n14_adj_4513, n48739, n45982, 
        n45942, n7_adj_4514, n45941, n10_adj_4515, n42254, n28715, 
        n28716, n3_adj_4516, n3_adj_4517, n48802, n48847, n8_adj_4518, 
        n26713, Kp_23__N_1099, n27401, n27188, n27133, n42512, n10_adj_4519, 
        n42779, n27289, n10_adj_4520, Kp_23__N_1093, n41737, n41649, 
        n45843, Kp_23__N_1096, n45844, n45842, n28717, n48685, n48703, 
        n14_adj_4521, n28718, n46847, n41777, n41687, n48679, n47464, 
        n42345, n42794, n42493, n28719, n45837, n45838, n45836, 
        n48673, n48781, n14_adj_4522, n42430, n41775, n41689, n41773, 
        n43514, n7_adj_4523, n8_adj_4524, n7_adj_4525, n33842, n28720, 
        n7_adj_4526, n8_adj_4527, n41771, n41693, n7_adj_4528, n8_adj_4529, 
        n7_adj_4530, n8_adj_4531, n41769, n41695, n41767, n41697, 
        n41765, n41699, n41763, n41701, n41761, n41703, n41759, 
        n41667, n41757, n41705, n41755, n41707, n33222, n41709, 
        n41753, n41711, n41751, n41663, n41749, n41713, n41747, 
        n41715, n26855, Kp_23__N_1064, n6_adj_4532, n42410, n42748, 
        n41745, n41717, n41743, n41719, n41741, n41721, n33220, 
        n8_adj_4533, n41739, n41657, n41661, n10_adj_4534, n41655, 
        n48857, n28721, n42763, n28722, n42354, n42717, n10_adj_4535, 
        Kp_23__N_1090, n42705, Kp_23__N_936, n42465, n42782, n26643, 
        n42658, n10_adj_4536, n4_adj_4537, Kp_23__N_988, n6_adj_4538, 
        n48817, n46828, n6_adj_4539, n48667, n48841, n47468, n42545, 
        Kp_23__N_993, n27125, n42766, n7_adj_4540, n42376, n42449, 
        n6958, n43203, n4_adj_4541, n42364, n42337, n42325, n6_adj_4542, 
        Kp_23__N_969, n48796, n42899, n10_adj_4543, n42726, n8_adj_4544, 
        n1168, n12_adj_4545, n42711, n32_adj_4546, n22_adj_4547, n36_adj_4548, 
        n42407, n34_adj_4549, n35_adj_4550, n42509, n6_adj_4551, n33_adj_4552, 
        n39558, n39596, n6_adj_4553, n42436, n26531, n10_adj_4554, 
        n12_adj_4555, n44557, Kp_23__N_1195, n7_adj_4556, n28_adj_4557, 
        n14_adj_4558, n48790, n42808, n15_adj_4559, n26_adj_4560, 
        n27_adj_4561, n25_adj_4562, n43705, n2_adj_4563, n3_adj_4564, 
        n28_adj_4565, n12_adj_4566, n10_adj_4567, n11_adj_4568, n9_adj_4569, 
        n42439, n42316, n26_adj_4570, n42496, n42723, n27_adj_4571, 
        n25_adj_4572, n42293, n48826, n33839, n26661, n42442, n42675, 
        n42537, n42340, n28_adj_4573, n31_adj_4574, n10_adj_4575, 
        n42426, n42947, n48778, n48772, n48766, n48760, n48754, 
        n48748, n48742, n48736, n2_adj_4576, n2_adj_4577, n2_adj_4578, 
        n41301, n41307, n41309, n42392, n42518, n42911, n42379, 
        n42357, n42487, n41315, n41321, n41327, n41349, n42, n30, 
        n34_adj_4579, n41365, n41385, n40_adj_4580, n26553, n41, 
        n39_adj_4581, n48, n43, n37_adj_4582, n38_adj_4583, n40476, 
        n14_adj_4584, n15_adj_4585, n40334, n41405, n41425, n41445, 
        n63, n63_adj_4586, n41477, n29_adj_4587, n41505, n6_adj_4589, 
        n4_adj_4590, n3_adj_4591, n48730, n8_adj_4592, n28699, n48700, 
        n48694, n48688, n28700, n23_adj_4593, n26_adj_4594, n29_adj_4595, 
        n22_adj_4596, n28701, n41525, n41547, n45700, n28702, n28703, 
        n42616, n41567, n48682, n33873, n26421, n41587, n3_adj_4597, 
        n5_adj_4598, n6_adj_4599, n42196, n48676, n41615, n3_adj_4600, 
        n41641, n3_adj_4601, n2_adj_4602, n3_adj_4603, n28769, n28768, 
        n28767, n28766, n28765, n28764, n28763, n28762, n28761, 
        n28760, n28759, n28758, n28757, n28756, n28755, n28754, 
        n28704, n27964, n43482, n28216, n2_adj_4604, n28705, n28753, 
        n28752, n28751, n28750, n28749, n28748, n28747, n32_adj_4605, 
        n27_adj_4606, n26539, n28706, n48670, n48664, n48658, n28698, 
        n28697, n28696, n28695, n28694, n28693, n7_adj_4607, n48652, 
        n7_adj_4608, n28680, n2_adj_4609, n2_adj_4610, n42735, n10_adj_4611, 
        n2_adj_4612, n48646, n28679, n28678, n28677, n2_adj_4613, 
        n28676, n2_adj_4614, n48640;
    wire [31:0]\FRAME_MATCHER.state_31__N_2724 ;
    
    wire n161, n33239, n12_adj_4615, n44481, n40258, n10_adj_4616, 
        n39625, n6_adj_4617, n7_adj_4618, n1_adj_4619, n3_adj_4620, 
        n48838, n48634, n28675, n47460, n28673, n8_adj_4621, n28672, 
        n33827, n48820, n48814, n48628, n33639, n33209, n43918, 
        n7_adj_4622, n48622, n7_adj_4623, n48610, n33300, n48604, 
        n48592, n42506, n4_adj_4624, n48586, n7_adj_4625, n99, n42235, 
        n126;
    wire [31:0]\FRAME_MATCHER.state_31__N_2660 ;
    
    wire n12_adj_4626, n48580, n37565, n37564, n10_adj_4627, n12_adj_4628, 
        n28671, n28670, n7_adj_4629, n48574, n8_adj_4630, n42627, 
        n27378, n37563, n37562, n37561, n37560, n2_adj_4631, n1_adj_4632, 
        n88, n37559, tx_transmit_N_3513, n37558, n6_adj_4633, n37557, 
        n64, n74, n37556, n37555, n37554, n37553, n37552, n37551, 
        n37550, n37549, n37548, n37547, n37546, n48568, n37545, 
        n37544, n37543, n44470, n26495, n3813, n6_adj_4634, n10_adj_4635, 
        n4_adj_4636;
    wire [31:0]\FRAME_MATCHER.state_31__N_2692 ;
    
    wire n37542, n37541, n37540, n1_adj_4637, n37539, n37538, n39584, 
        n28661, n26268, n37537, n37536, n37535, n37534, n37533, 
        n28660, n28659, n28658, n28656, n28655, n28654, n28653, 
        n37532, n28570, n28569, n28568, n28567, n28566, n28565, 
        n28564, n28563, n28562, n28561, n28560, n28559, n28558, 
        n28557, n37531, n28556, n28555, n28554, n28553, n28552, 
        n28551, n28550, n28549, n28548, n28547, n42445, n28538, 
        n28537, n28536, n28535, n28534, n28533, n28532, n28531, 
        n42772, n42599, n40510, n44349, n27252, n10_adj_4639, n37530, 
        n6_adj_4640, n6_adj_4641, n43547, n42652, n6_adj_4642, n37529, 
        n37528, n42853, n43849, n10_adj_4643, n42536, n42823, n33835, 
        n8_adj_4644, n6_adj_4646, n6_adj_4647, n42163, n4_adj_4648, 
        n121, n39569, n42579, n6_adj_4649, n26289, n4_adj_4650, 
        n8_adj_4651, n26414, n44, n42_adj_4652, n43_adj_4653, n27276, 
        n12_adj_4654, n41_adj_4655, n40_adj_4656, n42874, n39_adj_4657, 
        n50, n45, n26477, n10_adj_4658, n16_adj_4659, n11_adj_4660, 
        n10_adj_4661, n14_adj_4662, n45674, n16_adj_4663, n17_adj_4664, 
        n26403, n16_adj_4665, n17_adj_4666, n42400, n18_adj_4667, 
        n10_adj_4668, n42893, n42331, n14_adj_4669, n19_adj_4670, 
        n42856, n6_adj_4671, n68, n42929, n66, n67, n42971, n39510, 
        n65, n42515, n44671, n72, n70, n42610, n71, n69, n80, 
        n73, n81, n39580, n8_adj_4672, n42820, n39652, n42481, 
        n14_adj_4673, n15_adj_4674, n42932, n40455, n42935, n14_adj_4675, 
        n6_adj_4676, n14_adj_4677, n6_adj_4678;
    
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n28303));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[20] [6]), .I1(n42503), .I2(GND_net), 
            .I3(GND_net), .O(n39859));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 select_658_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_658_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n28302));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_863 (.I0(n39586), .I1(n40632), .I2(GND_net), 
            .I3(GND_net), .O(n42655));
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h9999;
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n28301));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n28300));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n28299));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n28298));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n28297));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n28296));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut (.I0(n42687), .I1(n24648), .I2(\data_out_frame[25] [4]), 
            .I3(GND_net), .O(n44126));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_LUT4 select_658_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4405));
    defparam select_658_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n27647), .D(n44528));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [5]), 
            .I2(\data_out_frame[19] [0]), .I3(n4_c), .O(n42923));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut (.I0(n42923), .I1(n40485), .I2(GND_net), .I3(GND_net), 
            .O(n10));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut (.I0(n42968), .I1(n40535), .I2(n42785), .I3(n40513), 
            .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n39685), .I1(n14), .I2(n10), .I3(n27602), 
            .O(n26860));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n27647), .D(n44126));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_658_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4406));
    defparam select_658_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n27647), .D(n43493));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_865 (.I0(n27027), .I1(n42699), .I2(n42944), .I3(\data_out_frame[15] [1]), 
            .O(n14_adj_4407));
    defparam i6_4_lut_adj_865.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n27647), .D(n44255));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n27647), .D(n43687));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n27647), .D(n44708));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(CLK_c), 
            .E(n27647), .D(n40583));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n28295));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(CLK_c), 
           .D(n28294));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(CLK_c), 
           .D(n28293));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n27647), .D(n43608));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_866 (.I0(n27558), .I1(n26965), .I2(n27257), .I3(GND_net), 
            .O(n42769));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_866.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_867 (.I0(n9), .I1(n14_adj_4407), .I2(n26860), 
            .I3(n40489), .O(n39586));
    defparam i7_4_lut_adj_867.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n28292));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_868 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42477));
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[10] [5]), .I1(n42702), .I2(n42965), 
            .I3(\data_out_frame[6] [1]), .O(n10_adj_4408));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n42367), .I1(n10_adj_4408), .I2(\data_out_frame[5] [6]), 
            .I3(GND_net), .O(n42788));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_869 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26722));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_870 (.I0(\data_out_frame[15] [1]), .I1(n40489), 
            .I2(GND_net), .I3(GND_net), .O(n27309));
    defparam i1_2_lut_adj_870.LUT_INIT = 16'h9999;
    SB_LUT4 i5_3_lut_adj_871 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[11] [1]), .I3(GND_net), .O(n14_adj_4409));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_871.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_872 (.I0(n42838), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[10] [6]), .I3(n42564), .O(n15));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_872.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n27329), .I2(n14_adj_4409), .I3(n26511), 
            .O(n27374));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_873 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[14] [7]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n42965));
    defparam i2_3_lut_adj_873.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_874 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n27329));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_874.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_875 (.I0(\data_out_frame[9] [2]), .I1(n27507), 
            .I2(n27257), .I3(n26965), .O(n10_adj_4410));
    defparam i4_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_876 (.I0(n39567), .I1(n26912), .I2(GND_net), 
            .I3(GND_net), .O(n42844));
    defparam i1_2_lut_adj_876.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_877 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42403));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_877.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33659 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [0]), .I2(\data_out_frame[23] [0]), 
            .I3(byte_transmit_counter[1]), .O(n48832));
    defparam byte_transmit_counter_0__bdd_4_lut_33659.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_4_lut_adj_878 (.I0(n42905), .I1(\data_out_frame[14] [0]), 
            .I2(n6_c), .I3(n42760), .O(n42576));
    defparam i2_4_lut_adj_878.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_879 (.I0(n42576), .I1(n42403), .I2(n42844), .I3(n40525), 
            .O(n42741));   // verilog/coms.v(71[16:27])
    defparam i2_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_880 (.I0(\data_out_frame[15] [3]), .I1(n39574), 
            .I2(\data_out_frame[15] [2]), .I3(GND_net), .O(n42348));
    defparam i2_3_lut_adj_880.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_881 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[12] [7]), .I3(n42313), .O(n10_adj_4411));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_881.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut (.I0(n26748), .I1(\data_out_frame[13] [1]), .I2(n10_adj_4411), 
            .I3(n27558), .O(n42484));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4412));
    defparam select_658_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4413));
    defparam select_658_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n42529), .I1(n42769), .I2(\data_out_frame[13] [4]), 
            .I3(\data_out_frame[11] [3]), .O(n12));   // verilog/coms.v(85[17:70])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_882 (.I0(n26097), .I1(n12), .I2(n42878), .I3(\data_out_frame[11] [2]), 
            .O(n39506));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_883 (.I0(n27507), .I1(n42814), .I2(n42385), .I3(n42452), 
            .O(n12_adj_4414));   // verilog/coms.v(85[17:70])
    defparam i5_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_884 (.I0(\data_out_frame[9] [1]), .I1(n12_adj_4414), 
            .I2(\data_out_frame[13] [5]), .I3(n42529), .O(n26912));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_884.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n1516), .I3(n42458), .O(n26989));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4415));
    defparam select_658_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4416));
    defparam select_658_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_885 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[8] [7]), 
            .I2(n42769), .I3(n6_adj_4417), .O(n27084));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_885.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4418));
    defparam select_658_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n48808_bdd_4_lut (.I0(n48808), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n48811));
    defparam n48808_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_658_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4419));
    defparam select_658_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 n48850_bdd_4_lut (.I0(n48850), .I1(\data_out_frame[21][2] ), 
            .I2(\data_out_frame[20] [2]), .I3(byte_transmit_counter[1]), 
            .O(n48853));
    defparam n48850_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i30730_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45861));
    defparam i30730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30731_4_lut (.I0(n45861), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n45862));
    defparam i30731_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i30729_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45860));
    defparam i30729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2079252_i1_3_lut (.I0(n48583), .I1(n48589), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4420));
    defparam i2079252_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31876_2_lut (.I0(n48793), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46849));
    defparam i31876_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i32326_3_lut (.I0(n48757), .I1(n48835), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n47458));
    defparam i32326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30725_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n45856));
    defparam i30725_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i30723_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45854));
    defparam i30723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2080458_i1_3_lut (.I0(n48751), .I1(n48613), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4421));
    defparam i2080458_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31886_2_lut (.I0(n48799), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46834));
    defparam i31886_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_886 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[25] [6]), 
            .I2(n42754), .I3(n6_adj_4422), .O(n44033));
    defparam i4_4_lut_adj_886.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n23237));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0104;
    SB_LUT4 select_658_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4423));
    defparam select_658_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_887 (.I0(n2134), .I1(\data_out_frame[24] [0]), 
            .I2(n42417), .I3(n6_adj_4424), .O(n43653));
    defparam i4_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n24129));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n28291));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30768_3_lut (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[17] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45899));
    defparam i30768_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n27701), .D(n8825[1]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30769_3_lut (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[19] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45900));
    defparam i30769_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4425));
    defparam select_658_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(CLK_c), 
            .E(n27701), .D(n8825[2]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
            .E(n27701), .D(n8825[3]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
            .E(n27701), .D(n8825[4]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
            .E(n27701), .D(n8825[5]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
            .E(n27701), .D(n8825[6]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
            .E(n27701), .D(n8825[7]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_888 (.I0(n42613), .I1(n2134), .I2(n27282), .I3(n42850), 
            .O(n10_adj_4426));
    defparam i4_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_889 (.I0(n40529), .I1(n10_adj_4426), .I2(\data_out_frame[24] [1]), 
            .I3(GND_net), .O(n44014));
    defparam i5_3_lut_adj_889.LUT_INIT = 16'h9696;
    SB_LUT4 select_658_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4427));
    defparam select_658_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_890 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(n27084), .I3(\data_out_frame[16] [0]), .O(n27602));   // verilog/coms.v(71[16:62])
    defparam i3_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i30775_3_lut (.I0(\data_out_frame[22] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45906));
    defparam i30775_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_891 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26899));
    defparam i1_2_lut_adj_891.LUT_INIT = 16'h6666;
    SB_LUT4 i30774_3_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[21][1] ), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45905));
    defparam i30774_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_658_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4428));
    defparam select_658_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4429));
    defparam select_658_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_892 (.I0(\data_out_frame[15] [0]), .I1(n27602), 
            .I2(GND_net), .I3(GND_net), .O(n42309));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_892.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_893 (.I0(n40485), .I1(n42696), .I2(n42309), .I3(\data_out_frame[16] [7]), 
            .O(n39685));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_893.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(CLK_c), 
           .D(n28290));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_894 (.I0(\data_out_frame[5] [1]), .I1(n42413), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n27507));
    defparam i1_2_lut_3_lut_adj_894.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[5] [1]), .I1(n42413), .I2(\data_out_frame[11] [6]), 
            .I3(n42757), .O(n42905));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30718_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45849));
    defparam i30718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30719_4_lut (.I0(n45849), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n45850));
    defparam i30719_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 select_658_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4430));
    defparam select_658_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30717_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45848));
    defparam i30717_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2081664_i1_3_lut (.I0(n48697), .I1(n48649), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4431));
    defparam i2081664_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_895 (.I0(n27282), .I1(n42521), .I2(n40487), .I3(GND_net), 
            .O(n43490));
    defparam i2_3_lut_adj_895.LUT_INIT = 16'h6969;
    SB_LUT4 select_658_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4432));
    defparam select_658_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_896 (.I0(\data_out_frame[22] [0]), .I1(n42953), 
            .I2(n42884), .I3(\data_out_frame[24] [3]), .O(n43563));
    defparam i3_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_897 (.I0(n42887), .I1(n42799), .I2(\data_out_frame[22] [1]), 
            .I3(n42956), .O(n10_adj_4433));
    defparam i4_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4434));
    defparam select_658_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4435));
    defparam select_658_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_898 (.I0(n42649), .I1(\data_in_frame[14] [5]), 
            .I2(\data_in_frame[19] [0]), .I3(n42868), .O(n10_adj_4436));
    defparam i4_4_lut_adj_898.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_899 (.I0(\data_in_frame[16] [6]), .I1(n10_adj_4436), 
            .I2(n40264), .I3(GND_net), .O(n44109));
    defparam i5_3_lut_adj_899.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_900 (.I0(\data_in_frame[19] [7]), .I1(n40531), 
            .I2(n40474), .I3(GND_net), .O(n39500));
    defparam i2_3_lut_adj_900.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_901 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[19] [4]), .I3(\data_in_frame[19] [5]), .O(n8));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_902 (.I0(\data_in_frame[19] [6]), .I1(n8), .I2(\data_in_frame[19] [3]), 
            .I3(\data_in_frame[19] [2]), .O(Kp_23__N_861));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_903 (.I0(Kp_23__N_861), .I1(n40531), .I2(GND_net), 
            .I3(GND_net), .O(n42573));
    defparam i1_2_lut_adj_903.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4437));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_905 (.I0(n26617), .I1(n27095), .I2(n42607), .I3(n6_adj_4437), 
            .O(n42881));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_905.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_906 (.I0(n40630), .I1(\data_in_frame[15] [5]), 
            .I2(n42720), .I3(n6_adj_4438), .O(n44174));
    defparam i4_4_lut_adj_906.LUT_INIT = 16'h9669;
    SB_LUT4 select_658_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4439));
    defparam select_658_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_907 (.I0(\data_in_frame[16] [7]), .I1(n42871), 
            .I2(n42811), .I3(\data_in_frame[16] [6]), .O(n40538));
    defparam i3_4_lut_adj_907.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4440));
    defparam select_658_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_908 (.I0(n42524), .I1(n39548), .I2(n40538), .I3(GND_net), 
            .O(n42714));
    defparam i2_3_lut_adj_908.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_909 (.I0(\data_in_frame[17] [0]), .I1(n26784), 
            .I2(n42791), .I3(n42490), .O(n42871));
    defparam i3_4_lut_adj_909.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_910 (.I0(n39908), .I1(n42558), .I2(n26938), .I3(n40613), 
            .O(n42649));
    defparam i1_4_lut_adj_910.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_911 (.I0(n39836), .I1(n42584), .I2(\data_in_frame[14] [4]), 
            .I3(GND_net), .O(n39908));
    defparam i2_3_lut_adj_911.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_912 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[14] [2]), 
            .I2(n26056), .I3(\data_in_frame[16] [4]), .O(n42868));
    defparam i3_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_913 (.I0(n42640), .I1(\data_in_frame[12] [1]), 
            .I2(\data_in_frame[11] [7]), .I3(n39616), .O(n14_adj_4441));
    defparam i6_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[14] [3]), .I1(n13), .I2(n14_adj_4441), 
            .I3(GND_net), .O(n40613));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_914 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [6]), .O(n42744));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_915 (.I0(n40613), .I1(n42587), .I2(n26025), .I3(GND_net), 
            .O(n40559));
    defparam i2_3_lut_adj_915.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_in_frame[9] [0]), .I1(n39793), .I2(n27215), 
            .I3(n42630), .O(n42631));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_916 (.I0(\data_in_frame[17] [5]), .I1(n42859), 
            .I2(n27436), .I3(n39606), .O(n10_adj_4442));
    defparam i4_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_917 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [3]), 
            .I2(\data_in_frame[14] [1]), .I3(GND_net), .O(n42587));
    defparam i2_3_lut_adj_917.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_918 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n26646));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_918.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_919 (.I0(\data_in_frame[13] [3]), .I1(n42841), 
            .I2(\data_in_frame[10] [6]), .I3(n42593), .O(n12_adj_4443));   // verilog/coms.v(85[17:70])
    defparam i5_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_920 (.I0(\data_in_frame[13] [2]), .I1(n12_adj_4443), 
            .I2(\data_in_frame[15] [4]), .I3(n42708), .O(n39606));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_920.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_921 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42590));
    defparam i1_2_lut_adj_921.LUT_INIT = 16'h6666;
    SB_LUT4 i14_4_lut (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[9] [6]), 
            .I2(n39793), .I3(n42890), .O(n36));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[7] [4]), 
            .I2(n42847), .I3(n42468), .O(n34));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(\data_in_frame[10] [0]), .I1(n36), .I2(n26), 
            .I3(\data_in_frame[9] [4]), .O(n40));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[6] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(n26646), .O(n38));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_3_lut (.I0(\data_in_frame[3] [0]), .I1(n34), .I2(\data_in_frame[9] [5]), 
            .I3(GND_net), .O(n39));
    defparam i17_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut (.I0(n42805), .I1(n42462), .I2(n42729), .I3(\data_in_frame[5] [1]), 
            .O(n37));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n26056));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n28289));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_922 (.I0(\data_in_frame[8] [2]), .I1(n26687), .I2(n27551), 
            .I3(n6_adj_4444), .O(n42890));
    defparam i4_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\data_in_frame[9] [1]), .I1(n39554), .I2(GND_net), 
            .I3(GND_net), .O(n42682));
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_924 (.I0(n26581), .I1(n42682), .I2(\data_in_frame[9] [4]), 
            .I3(GND_net), .O(n42640));
    defparam i2_3_lut_adj_924.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut (.I0(n27203), .I1(n27451), .I2(\data_in_frame[9] [0]), 
            .I3(\data_in_frame[11] [7]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut (.I0(n39321), .I1(n42631), .I2(\data_in_frame[9] [6]), 
            .I3(GND_net), .O(n17));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_925 (.I0(\data_out_frame[19] [1]), .I1(n42309), 
            .I2(\data_out_frame[18] [7]), .I3(n26899), .O(n13_adj_4445));
    defparam i5_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_926 (.I0(n42682), .I1(n27199), .I2(\data_in_frame[12] [0]), 
            .I3(n27588), .O(n22));
    defparam i8_4_lut_adj_926.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_927 (.I0(n17), .I1(n24), .I2(\data_in_frame[13] [7]), 
            .I3(n42890), .O(n26_adj_4446));
    defparam i12_4_lut_adj_927.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(\data_in_frame[11] [5]), .I1(n26_adj_4446), .I2(n22), 
            .I3(\data_in_frame[9] [2]), .O(n26025));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_928 (.I0(\data_out_frame[7] [3]), .I1(n24129), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n42757));
    defparam i1_2_lut_3_lut_adj_928.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_929 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42862));
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_930 (.I0(n13_adj_4445), .I1(n11), .I2(n40535), 
            .I3(n39685), .O(n42699));
    defparam i7_4_lut_adj_930.LUT_INIT = 16'h9669;
    SB_LUT4 i31866_2_lut (.I0(n48805), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46829));
    defparam i31866_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_931 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[13] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42607));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_931.LUT_INIT = 16'h6666;
    SB_LUT4 i32330_3_lut (.I0(n48691), .I1(n48853), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n47462));
    defparam i32330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_932 (.I0(\data_in_frame[18] [3]), .I1(n42607), 
            .I2(\data_in_frame[14] [1]), .I3(n42862), .O(n16));
    defparam i6_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_933 (.I0(n26025), .I1(n42640), .I2(\data_in_frame[16] [1]), 
            .I3(n8_adj_4447), .O(n17_adj_4448));
    defparam i7_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17_adj_4448), .I1(\data_in_frame[16] [2]), .I2(n16), 
            .I3(\data_in_frame[11] [5]), .O(n42551));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_934 (.I0(n40481), .I1(n26056), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4449));
    defparam i2_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_935 (.I0(n42590), .I1(\data_in_frame[14] [0]), 
            .I2(n26756), .I3(n27203), .O(n14_adj_4450));
    defparam i6_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_936 (.I0(\data_in_frame[16] [3]), .I1(n14_adj_4450), 
            .I2(n10_adj_4449), .I3(n27071), .O(n40557));
    defparam i7_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\data_in_frame[17] [6]), .I1(n39606), 
            .I2(GND_net), .I3(GND_net), .O(n42950));
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_938 (.I0(n40557), .I1(n42551), .I2(\data_in_frame[18] [4]), 
            .I3(GND_net), .O(n42829));
    defparam i2_3_lut_adj_938.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_939 (.I0(\data_in_frame[11] [6]), .I1(n42646), 
            .I2(n40499), .I3(n40457), .O(n40481));
    defparam i3_4_lut_adj_939.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4451));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_941 (.I0(n42322), .I1(n40481), .I2(n42708), .I3(n6_adj_4451), 
            .O(n42826));   // verilog/coms.v(72[16:41])
    defparam i4_4_lut_adj_941.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_942 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42832));
    defparam i1_2_lut_adj_942.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_943 (.I0(\data_in_frame[16] [1]), .I1(n42832), 
            .I2(\data_in_frame[14] [0]), .I3(\data_in_frame[13] [5]), .O(n42322));   // verilog/coms.v(72[16:41])
    defparam i3_4_lut_adj_943.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42646));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_945 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27436));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_945.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_946 (.I0(n31), .I1(n31_adj_4452), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(n42248), .O(n7_c));
    defparam i1_2_lut_4_lut_adj_946.LUT_INIT = 16'hffca;
    SB_LUT4 i7_4_lut_adj_947 (.I0(\data_in_frame[13] [3]), .I1(n42296), 
            .I2(n40521), .I3(\data_in_frame[11] [1]), .O(n18));
    defparam i7_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_948 (.I0(Kp_23__N_1306), .I1(n18), .I2(n42500), 
            .I3(Kp_23__N_1330), .O(n20_c));
    defparam i9_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_949 (.I0(n15_adj_4453), .I1(n20_c), .I2(n42631), 
            .I3(n26581), .O(n39918));
    defparam i10_4_lut_adj_949.LUT_INIT = 16'h9669;
    SB_LUT4 i20323_2_lut_4_lut (.I0(n31), .I1(n31_adj_4452), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(n23788), .O(n1));
    defparam i20323_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\data_in_frame[16] [0]), .I1(n39918), 
            .I2(GND_net), .I3(GND_net), .O(n40630));
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_951 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[11] [6]), 
            .I2(\data_in_frame[12] [1]), .I3(GND_net), .O(n42847));
    defparam i2_3_lut_adj_951.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_952 (.I0(n39793), .I1(n39598), .I2(\data_in_frame[10] [7]), 
            .I3(n26809), .O(n42296));
    defparam i3_4_lut_adj_952.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42490));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\data_in_frame[12] [3]), .I1(n39321), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4454));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_955 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[10] [0]), 
            .I2(\data_in_frame[10] [2]), .I3(n6_adj_4454), .O(n42584));
    defparam i4_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_956 (.I0(\data_in_frame[11] [7]), .I1(n42334), 
            .I2(n42584), .I3(\data_in_frame[10] [3]), .O(n32));
    defparam i12_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[9] [3]), 
            .I2(n42490), .I3(n39554), .O(n31_adj_4455));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_957 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[12] [6]), 
            .I2(n27137), .I3(\data_in_frame[12] [4]), .O(n35));
    defparam i15_4_lut_adj_957.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_958 (.I0(n42471), .I1(\data_in_frame[10] [1]), 
            .I2(n42296), .I3(n26801), .O(n34_adj_4456));
    defparam i14_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_LUT4 i18_3_lut (.I0(n35), .I1(n31_adj_4455), .I2(n32), .I3(GND_net), 
            .O(n38_adj_4457));
    defparam i18_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13_4_lut_adj_959 (.I0(n27196), .I1(n42847), .I2(n27071), 
            .I3(n42548), .O(n33));
    defparam i13_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_960 (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[14] [7]), .I3(n42865), .O(n36_adj_4458));
    defparam i14_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_961 (.I0(n33), .I1(n40630), .I2(n38_adj_4457), 
            .I3(n34_adj_4456), .O(n25));
    defparam i3_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_962 (.I0(\data_in_frame[13] [3]), .I1(n27436), 
            .I2(n42646), .I3(n42322), .O(n34_adj_4459));
    defparam i12_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[15] [5]), 
            .I2(n42826), .I3(GND_net), .O(n20_adj_4460));
    defparam i6_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_963 (.I0(n42829), .I1(\data_in_frame[18] [5]), 
            .I2(n39918), .I3(n42950), .O(n23));
    defparam i9_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 i2022_2_lut_3_lut (.I0(n31_adj_4452), .I1(n23788), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n7001));
    defparam i2022_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i18_4_lut_adj_964 (.I0(n25), .I1(n36_adj_4458), .I2(n42590), 
            .I3(\data_in_frame[16] [6]), .O(n40_adj_4461));
    defparam i18_4_lut_adj_964.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n7001), .I3(GND_net), .O(n7003));
    defparam mux_2022_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n7001), .I3(GND_net), .O(n7004));
    defparam mux_2022_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n7001), .I3(GND_net), .O(n7005));
    defparam mux_2022_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut_adj_965 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[14] [4]), 
            .I2(n27095), .I3(\data_in_frame[14] [3]), .O(n38_adj_4462));
    defparam i16_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n7001), .I3(GND_net), .O(n7006));
    defparam mux_2022_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17_3_lut_adj_966 (.I0(\data_in_frame[15] [7]), .I1(n34_adj_4459), 
            .I2(\data_in_frame[15] [1]), .I3(GND_net), .O(n39_adj_4463));
    defparam i17_3_lut_adj_966.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut_adj_967 (.I0(n42637), .I1(n42302), .I2(n42587), 
            .I3(\data_in_frame[15] [3]), .O(n37_adj_4464));
    defparam i15_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n7001), .I3(GND_net), .O(n7007));
    defparam mux_2022_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_4_lut_adj_968 (.I0(n15_adj_4465), .I1(n44139), .I2(n40559), 
            .I3(n27234), .O(n22_adj_4466));
    defparam i8_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_969 (.I0(n23), .I1(n42868), .I2(n20_adj_4460), 
            .I3(n42811), .O(n26_adj_4467));
    defparam i12_4_lut_adj_969.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_970 (.I0(n37_adj_4464), .I1(n39_adj_4463), .I2(n38_adj_4462), 
            .I3(n40_adj_4461), .O(n44102));
    defparam i21_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_971 (.I0(n44102), .I1(n26_adj_4467), .I2(n22_adj_4466), 
            .I3(\data_in_frame[17] [7]), .O(n40474));
    defparam i13_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n7001), .I3(GND_net), .O(n7008));
    defparam mux_2022_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n7001), .I3(GND_net), .O(n7009));
    defparam mux_2022_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n7001), .I3(GND_net), .O(n7010));
    defparam mux_2022_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n7001), .I3(GND_net), .O(n7011));
    defparam mux_2022_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_972 (.I0(n31_adj_4452), .I1(n23788), .I2(\FRAME_MATCHER.state_c [2]), 
            .I3(n26496), .O(n27617));
    defparam i2_3_lut_4_lut_adj_972.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_adj_973 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[10] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42334));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_973.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_974 (.I0(n40566), .I1(n42685), .I2(n26801), .I3(n42433), 
            .O(n39836));
    defparam i3_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n7001), .I3(GND_net), .O(n7012));
    defparam mux_2022_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n7001), .I3(GND_net), .O(n7013));
    defparam mux_2022_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_975 (.I0(\data_in_frame[12] [4]), .I1(n26938), 
            .I2(\data_in_frame[10] [2]), .I3(n39836), .O(n44477));
    defparam i3_4_lut_adj_975.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2), .S(n3_adj_4468));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_2022_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n7001), .I3(GND_net), .O(n7014));
    defparam mux_2022_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n7001), .I3(GND_net), .O(n7015));
    defparam mux_2022_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_976 (.I0(\data_in_frame[14] [6]), .I1(n26938), 
            .I2(n44477), .I3(n26789), .O(n42791));
    defparam i3_4_lut_adj_976.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_977 (.I0(\data_in_frame[9] [0]), .I1(n39793), .I2(n27215), 
            .I3(GND_net), .O(n40472));
    defparam i2_3_lut_adj_977.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_978 (.I0(n39554), .I1(n26809), .I2(GND_net), 
            .I3(GND_net), .O(n40457));
    defparam i1_2_lut_adj_978.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2022_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n7001), .I3(GND_net), .O(n7016));
    defparam mux_2022_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_979 (.I0(n27084), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[14] [6]), .I3(n42484), .O(n28));
    defparam i12_4_lut_adj_979.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_980 (.I0(n26756), .I1(n42561), .I2(\data_in_frame[8] [0]), 
            .I3(GND_net), .O(n27551));
    defparam i2_3_lut_adj_980.LUT_INIT = 16'h9696;
    SB_LUT4 i15217_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n28731));
    defparam i15217_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1306));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42548));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h6666;
    SB_LUT4 mux_2022_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n7001), .I3(GND_net), .O(n7017));
    defparam mux_2022_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n7001), .I3(GND_net), .O(n7018));
    defparam mux_2022_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n7001), .I3(GND_net), .O(n7019));
    defparam mux_2022_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n7001), .I3(GND_net), .O(n7020));
    defparam mux_2022_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n7001), .I3(GND_net), .O(n7021));
    defparam mux_2022_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_2022_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n7001), .I3(GND_net), .O(n7022));
    defparam mux_2022_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_982 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26581));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_983 (.I0(n42775), .I1(\data_out_frame[14] [3]), 
            .I2(n1519), .I3(\data_out_frame[15] [4]), .O(n26_adj_4470));
    defparam i10_4_lut_adj_983.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_in_frame[9] [4]), .I1(n39598), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4471));
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_985 (.I0(n26581), .I1(n42548), .I2(Kp_23__N_1306), 
            .I3(n6_adj_4471), .O(n42630));
    defparam i4_4_lut_adj_985.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n7001), .I3(GND_net), .O(n7023));
    defparam mux_2022_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_986 (.I0(n26667), .I1(n27551), .I2(n40521), .I3(n24724), 
            .O(n12_adj_4472));
    defparam i5_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n7001), .I3(GND_net), .O(n7024));
    defparam mux_2022_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_987 (.I0(n26801), .I1(n12_adj_4472), .I2(n42593), 
            .I3(n40494), .O(n39793));
    defparam i6_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27137));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_989 (.I0(n8_adj_4447), .I1(n27137), .I2(n39793), 
            .I3(n42630), .O(n10_adj_4473));
    defparam i4_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_990 (.I0(n42920), .I1(n42348), .I2(n42741), 
            .I3(n40492), .O(n27));
    defparam i11_4_lut_adj_990.LUT_INIT = 16'h9669;
    SB_LUT4 mux_2022_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n7001), .I3(GND_net), .O(n7025));
    defparam mux_2022_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_991 (.I0(n26789), .I1(n27215), .I2(GND_net), 
            .I3(GND_net), .O(n26667));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_991.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_992 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42865));
    defparam i1_2_lut_adj_992.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_993 (.I0(n26633), .I1(\data_in_frame[17] [4]), 
            .I2(n42865), .I3(n27407), .O(n16_adj_4474));
    defparam i6_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_994 (.I0(n26667), .I1(n42859), .I2(n42941), .I3(\data_in_frame[13] [2]), 
            .O(n17_adj_4475));
    defparam i7_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_995 (.I0(n17_adj_4475), .I1(\data_in_frame[10] [4]), 
            .I2(n16_adj_4474), .I3(n26784), .O(n27104));
    defparam i9_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_996 (.I0(n42567), .I1(n42791), .I2(\data_in_frame[17] [2]), 
            .I3(\data_in_frame[13] [0]), .O(n12_adj_4476));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_997 (.I0(n27227), .I1(n12_adj_4476), .I2(n42835), 
            .I3(\data_in_frame[12] [5]), .O(n39548));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_997.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_998 (.I0(n42649), .I1(n42871), .I2(n42302), .I3(GND_net), 
            .O(n40264));
    defparam i2_3_lut_adj_998.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_999 (.I0(n39548), .I1(n27104), .I2(GND_net), 
            .I3(GND_net), .O(n39631));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1000 (.I0(n42370), .I1(n42555), .I2(\data_in_frame[18] [0]), 
            .I3(n40474), .O(n12_adj_4477));
    defparam i5_4_lut_adj_1000.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1001 (.I0(n44139), .I1(n12_adj_4477), .I2(n42832), 
            .I3(\data_in_frame[16] [0]), .O(n40531));
    defparam i6_4_lut_adj_1001.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1002 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n27407));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1003 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4478));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1003.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1004 (.I0(n27451), .I1(n27246), .I2(n42319), 
            .I3(n6_adj_4478), .O(n42433));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42567));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1006 (.I0(n26784), .I1(n42433), .I2(GND_net), 
            .I3(GND_net), .O(n24724));
    defparam i1_2_lut_adj_1006.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1007 (.I0(\data_in_frame[15] [0]), .I1(n5), .I2(GND_net), 
            .I3(GND_net), .O(n42835));
    defparam i1_2_lut_adj_1007.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1008 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26633));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1008.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(\data_in_frame[9] [7]), .I1(n27451), 
            .I2(GND_net), .I3(GND_net), .O(n42729));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1010 (.I0(n42962), .I1(\data_in_frame[10] [1]), 
            .I2(n42328), .I3(n42902), .O(n15_adj_4479));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1011 (.I0(n15_adj_4479), .I1(n42389), .I2(n14_adj_4480), 
            .I3(n26968), .O(n39616));   // verilog/coms.v(78[16:27])
    defparam i8_4_lut_adj_1011.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1012 (.I0(n39616), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n42558));
    defparam i2_3_lut_adj_1012.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42361));
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1014 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[14] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42938));
    defparam i1_2_lut_adj_1014.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1015 (.I0(n26789), .I1(n42938), .I2(n42361), 
            .I3(n42558), .O(n12_adj_4481));
    defparam i5_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1016 (.I0(n26633), .I1(n12_adj_4481), .I2(\data_in_frame[17] [1]), 
            .I3(n42835), .O(n42524));
    defparam i6_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1017 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[17] [3]), 
            .I2(n42841), .I3(n42361), .O(n16_adj_4482));
    defparam i6_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1018 (.I0(n26912), .I1(n39506), .I2(n26989), 
            .I3(GND_net), .O(n42920));
    defparam i1_2_lut_3_lut_adj_1018.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1019 (.I0(n24724), .I1(n42567), .I2(n42941), 
            .I3(n27215), .O(n17_adj_4483));
    defparam i7_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1020 (.I0(n17_adj_4483), .I1(\data_in_frame[10] [3]), 
            .I2(n16_adj_4482), .I3(\data_in_frame[15] [2]), .O(n27234));
    defparam i9_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1021 (.I0(Kp_23__N_1214), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n42561));
    defparam i2_3_lut_adj_1021.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42471));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(n26756), .I1(n27196), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1330));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1024 (.I0(n42965), .I1(n42689), .I2(n27374), 
            .I3(n1668), .O(n25_adj_4484));
    defparam i9_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1025 (.I0(n42720), .I1(\data_in_frame[13] [4]), 
            .I2(n42370), .I3(GND_net), .O(n42500));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1025.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1026 (.I0(n42881), .I1(n44174), .I2(\data_in_frame[15] [6]), 
            .I3(n42950), .O(n10_adj_4485));
    defparam i4_4_lut_adj_1026.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1027 (.I0(n42500), .I1(n10_adj_4485), .I2(\data_in_frame[18] [0]), 
            .I3(GND_net), .O(n39516));
    defparam i5_3_lut_adj_1027.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4486));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_DFFSR tx_transmit_3871 (.Q(\r_SM_Main_2__N_3616[0] ), .C(CLK_c), 
            .D(n4888[0]), .R(n43197));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1029 (.I0(n27234), .I1(n42524), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4487));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1030 (.I0(n39516), .I1(n44139), .I2(n27104), 
            .I3(GND_net), .O(n6_adj_4488));
    defparam i1_3_lut_adj_1030.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1031 (.I0(n42714), .I1(n8_adj_4489), .I2(n44139), 
            .I3(n27104), .O(n10_adj_4490));
    defparam i4_4_lut_adj_1031.LUT_INIT = 16'h9669;
    SB_LUT4 n48832_bdd_4_lut (.I0(n48832), .I1(\data_out_frame[21][0] ), 
            .I2(\data_out_frame[20] [0]), .I3(byte_transmit_counter[1]), 
            .O(n48835));
    defparam n48832_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_1032 (.I0(n25_adj_4484), .I1(n27), .I2(n26_adj_4470), 
            .I3(n28), .O(n40489));
    defparam i15_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n27647), .D(n43569));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1033 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n42620));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n27685), .D(n7002));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1034 (.I0(\data_in_frame[19] [6]), .I1(n39500), 
            .I2(\data_in_frame[20] [0]), .I3(n6_adj_4488), .O(n44433));
    defparam i4_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n27647), .D(n43617));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1035 (.I0(\data_out_frame[17] [1]), .I1(n1519), 
            .I2(n42788), .I3(n42785), .O(n43671));
    defparam i3_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(n40489), .I1(n42699), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4491));
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'h6666;
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n27647), .D(n43563));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut_adj_1037 (.I0(\data_in_frame[19] [3]), .I1(n42714), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[21] [4]), .O(n43611));
    defparam i2_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1038 (.I0(n40620), .I1(\data_in_frame[20] [7]), 
            .I2(n42573), .I3(GND_net), .O(n8_adj_4492));
    defparam i3_3_lut_adj_1038.LUT_INIT = 16'h6969;
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n27647), .D(n43490));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1039 (.I0(\data_out_frame[21][3] ), .I1(n43671), 
            .I2(n42620), .I3(n6_adj_4491), .O(n39556));
    defparam i4_4_lut_adj_1039.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1040 (.I0(n44174), .I1(\data_in_frame[18] [1]), 
            .I2(\data_in_frame[20] [3]), .I3(n42826), .O(n43826));
    defparam i2_4_lut_adj_1040.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1041 (.I0(n40557), .I1(\data_in_frame[18] [4]), 
            .I2(n40620), .I3(\data_in_frame[20] [6]), .O(n44504));
    defparam i3_4_lut_adj_1041.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1042 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[21] [2]), 
            .I2(n44109), .I3(GND_net), .O(n44257));
    defparam i2_3_lut_adj_1042.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut_adj_1043 (.I0(n39631), .I1(\data_in_frame[19] [4]), 
            .I2(\data_in_frame[21] [6]), .I3(\data_in_frame[19] [5]), .O(n44269));
    defparam i2_4_lut_adj_1043.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1044 (.I0(n42551), .I1(n42826), .I2(\data_in_frame[20] [4]), 
            .I3(GND_net), .O(n43861));
    defparam i2_3_lut_adj_1044.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1045 (.I0(n42524), .I1(n27104), .I2(n40538), 
            .I3(\data_in_frame[21] [0]), .O(n12_adj_4493));
    defparam i5_4_lut_adj_1045.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1046 (.I0(n5_adj_4486), .I1(n44139), .I2(\data_in_frame[19] [6]), 
            .I3(n27234), .O(n43516));
    defparam i3_4_lut_adj_1046.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1047 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[20] [5]), 
            .I2(n4_adj_4494), .I3(n42829), .O(n18_adj_4495));
    defparam i2_4_lut_adj_1047.LUT_INIT = 16'hde7b;
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n28288));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1048 (.I0(n44139), .I1(n42573), .I2(n27104), 
            .I3(n44109), .O(n11_adj_4496));
    defparam i4_4_lut_adj_1048.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1049 (.I0(\data_in_frame[21] [5]), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[19] [4]), .I3(n6_adj_4487), .O(n44400));
    defparam i4_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1050 (.I0(Kp_23__N_861), .I1(n44433), .I2(n10_adj_4490), 
            .I3(\data_in_frame[21] [1]), .O(n20_adj_4497));
    defparam i4_4_lut_adj_1050.LUT_INIT = 16'hdeed;
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n27647), .D(n44014));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n27647), .D(n43653));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1051 (.I0(\data_in_frame[20] [1]), .I1(n44174), 
            .I2(n39500), .I3(GND_net), .O(n44600));
    defparam i2_3_lut_adj_1051.LUT_INIT = 16'h6969;
    SB_LUT4 i9_4_lut_adj_1052 (.I0(n11_adj_4496), .I1(n18_adj_4495), .I2(n43516), 
            .I3(n12_adj_4493), .O(n25_adj_4498));
    defparam i9_4_lut_adj_1052.LUT_INIT = 16'hdfef;
    SB_LUT4 i30646_4_lut (.I0(n40538), .I1(n43611), .I2(n8_adj_4499), 
            .I3(\data_in_frame[21] [3]), .O(n45678));
    defparam i30646_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26527));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_LUT4 i15218_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n28732));
    defparam i15218_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n27647), .D(n44033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n28287));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i169 (.Q(\data_out_frame[21][0] ), .C(CLK_c), 
           .D(n28286));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_658_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4500));
    defparam select_658_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42738));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i170 (.Q(\data_out_frame[21][1] ), .C(CLK_c), 
           .D(n28285));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15219_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n28733));
    defparam i15219_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30648_4_lut (.I0(n43826), .I1(n44139), .I2(n8_adj_4492), 
            .I3(\data_in_frame[19] [0]), .O(n45680));
    defparam i30648_4_lut.LUT_INIT = 16'h2882;
    SB_LUT4 i15220_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n28734));
    defparam i15220_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1055 (.I0(n42395), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[4] [0]), .I3(n42738), .O(n10_adj_4501));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1056 (.I0(n43861), .I1(n44269), .I2(n44257), 
            .I3(n44504), .O(n27_adj_4502));
    defparam i11_4_lut_adj_1056.LUT_INIT = 16'hfbff;
    SB_LUT4 i15221_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n28735));
    defparam i15221_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1057 (.I0(n25_adj_4498), .I1(n44600), .I2(n20_adj_4497), 
            .I3(n44400), .O(n29));
    defparam i13_4_lut_adj_1057.LUT_INIT = 16'hfffb;
    SB_LUT4 i15_4_lut_adj_1058 (.I0(n29), .I1(n27_adj_4502), .I2(n45680), 
            .I3(n45678), .O(n31));
    defparam i15_4_lut_adj_1058.LUT_INIT = 16'hefff;
    SB_LUT4 i3_4_lut_adj_1059 (.I0(n42305), .I1(n42817), .I2(n42732), 
            .I3(n42533), .O(n1519));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(n1519), .I1(n1516), .I2(GND_net), .I3(GND_net), 
            .O(n27027));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42564));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'h6666;
    SB_LUT4 select_658_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4503));
    defparam select_658_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15222_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n28736));
    defparam i15222_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15223_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n28737));
    defparam i15223_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1062 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[11] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42385));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1062.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i171 (.Q(\data_out_frame[21][2] ), .C(CLK_c), 
           .D(n28284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i172 (.Q(\data_out_frame[21][3] ), .C(CLK_c), 
           .D(n28283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i173 (.Q(\data_out_frame[21][4] ), .C(CLK_c), 
           .D(n28282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(CLK_c), 
           .D(n28281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(CLK_c), 
           .D(n28280));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(CLK_c), 
           .D(n28279));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_658_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4504));
    defparam select_658_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(CLK_c), 
           .D(n28278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(CLK_c), 
           .D(n28277));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30700_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45831));
    defparam i30700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31864_2_lut (.I0(n48823), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46815));
    defparam i31864_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(CLK_c), 
           .D(n28276));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1063 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42533));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1064 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n42367));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1064.LUT_INIT = 16'h9696;
    SB_LUT4 i30859_4_lut (.I0(\data_out_frame[20] [5]), .I1(n46815), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[0]), .O(n45990));
    defparam i30859_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33669 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [3]), .I2(\data_out_frame[23] [3]), 
            .I3(byte_transmit_counter[1]), .O(n48844));
    defparam byte_transmit_counter_0__bdd_4_lut_33669.LUT_INIT = 16'he4aa;
    SB_LUT4 i15224_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42281), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n28738));
    defparam i15224_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i20_3_lut (.I0(\data_out_frame[22] [5]), 
            .I1(\data_out_frame[23] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4505));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_out_frame[11] [2]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42959));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1066 (.I0(\data_out_frame[8] [3]), .I1(n42693), 
            .I2(\data_out_frame[4] [0]), .I3(n42367), .O(n12_adj_4506));   // verilog/coms.v(85[17:63])
    defparam i5_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i30701_4_lut (.I0(n45831), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n45832));
    defparam i30701_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i30699_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45830));
    defparam i30699_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(CLK_c), 
           .D(n28275));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2085282_i1_3_lut (.I0(n48577), .I1(n48769), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4507));
    defparam i2085282_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30814_4_lut (.I0(n48775), .I1(n45991), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n45945));
    defparam i30814_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30813_3_lut (.I0(n7_adj_4508), .I1(n14_adj_4507), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n45944));
    defparam i30813_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(CLK_c), 
           .D(n28274));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30815_3_lut (.I0(n45944), .I1(n45945), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[5]));
    defparam i30815_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n28273));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i31861_2_lut (.I0(n48829), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46817));
    defparam i31861_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i30853_4_lut (.I0(\data_out_frame[20] [6]), .I1(n46817), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[0]), .O(n45984));
    defparam i30853_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 equal_299_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4469));   // verilog/coms.v(154[7:23])
    defparam equal_299_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42274), .I3(\FRAME_MATCHER.i [0]), .O(n42276));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i20_3_lut (.I0(\data_out_frame[22] [6]), 
            .I1(\data_out_frame[23] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4509));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30695_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n45826));
    defparam i30695_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1067 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42281), .I3(\FRAME_MATCHER.i [0]), .O(n42287));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1067.LUT_INIT = 16'hfbff;
    SB_LUT4 i30693_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45824));
    defparam i30693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1068 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42260), .I3(\FRAME_MATCHER.i [0]), .O(n42266));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1068.LUT_INIT = 16'hfbff;
    SB_LUT4 i2085885_i1_3_lut (.I0(n48763), .I1(n48595), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4510));
    defparam i2085885_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30685_4_lut (.I0(n48745), .I1(n45985), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n45816));
    defparam i30685_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30684_3_lut (.I0(n7_adj_4511), .I1(n14_adj_4510), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n45815));
    defparam i30684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30686_3_lut (.I0(n45815), .I1(n45816), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[6]));
    defparam i30686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31859_2_lut (.I0(n48571), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46819));
    defparam i31859_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i30850_4_lut (.I0(\data_out_frame[20] [7]), .I1(n46819), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[0]), .O(n45981));
    defparam i30850_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i20_3_lut (.I0(\data_out_frame[22] [7]), 
            .I1(\data_out_frame[23] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n20_adj_4512));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30689_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n45820));
    defparam i30689_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i30687_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45818));
    defparam i30687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2086488_i1_3_lut (.I0(n48733), .I1(n48607), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4513));
    defparam i2086488_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30811_4_lut (.I0(n48739), .I1(n45982), .I2(byte_transmit_counter[3]), 
            .I3(byte_transmit_counter[2]), .O(n45942));
    defparam i30811_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30810_3_lut (.I0(n7_adj_4514), .I1(n14_adj_4513), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n45941));
    defparam i30810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15201_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n28715));
    defparam i15201_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15202_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n28716));
    defparam i15202_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30812_3_lut (.I0(n45941), .I1(n45942), .I2(byte_transmit_counter[4]), 
            .I3(GND_net), .O(tx_data[7]));
    defparam i30812_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42468));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 select_658_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4516));
    defparam select_658_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4517));
    defparam select_658_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33634 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n48802));
    defparam byte_transmit_counter_0__bdd_4_lut_33634.LUT_INIT = 16'he4aa;
    SB_LUT4 n48844_bdd_4_lut (.I0(n48844), .I1(\data_out_frame[21][3] ), 
            .I2(\data_out_frame[20] [3]), .I3(byte_transmit_counter[1]), 
            .O(n48847));
    defparam n48844_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_adj_1070 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[0] [7]), 
            .I2(n8_adj_4518), .I3(n26713), .O(n27451));
    defparam i1_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1071 (.I0(\data_in_frame[4] [5]), .I1(Kp_23__N_1099), 
            .I2(n27401), .I3(n42468), .O(Kp_23__N_1214));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 equal_2186_i8_2_lut (.I0(Kp_23__N_1214), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4447));   // verilog/coms.v(236[9:81])
    defparam equal_2186_i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1072 (.I0(n27188), .I1(n12_adj_4506), .I2(n42305), 
            .I3(n42564), .O(n42313));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1073 (.I0(n26646), .I1(n27401), .I2(n27133), 
            .I3(n42512), .O(n10_adj_4519));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n28272));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_adj_1074 (.I0(\data_in_frame[4] [6]), .I1(n10_adj_4519), 
            .I2(\data_in_frame[7] [0]), .I3(GND_net), .O(n26756));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_adj_1074.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1075 (.I0(n42779), .I1(n27289), .I2(\data_in_frame[7] [2]), 
            .I3(n26968), .O(n10_adj_4520));
    defparam i4_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n28271));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1076 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_1093), 
            .I2(GND_net), .I3(GND_net), .O(n27199));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1076.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(CLK_c), 
            .D(n41737), .S(n41649));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30712_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45843));
    defparam i30712_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1077 (.I0(Kp_23__N_1096), .I1(\data_in_frame[8] [5]), 
            .I2(\data_in_frame[6] [3]), .I3(GND_net), .O(n42462));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1077.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\data_in_frame[5] [4]), .I1(\data_in_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42902));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_LUT4 i30713_4_lut (.I0(n45843), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n45844));
    defparam i30713_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i30711_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45842));
    defparam i30711_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42693));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i15203_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n28717));
    defparam i15203_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2082870_i1_3_lut (.I0(n48685), .I1(n48703), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4521));
    defparam i2082870_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15204_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n28718));
    defparam i15204_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n48802_bdd_4_lut (.I0(n48802), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n48805));
    defparam n48802_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i31786_2_lut (.I0(n48811), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46847));
    defparam i31786_2_lut.LUT_INIT = 16'h2222;
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(CLK_c), 
            .D(n41777), .S(n41687));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i32332_3_lut (.I0(n48679), .I1(n48847), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n47464));
    defparam i32332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1080 (.I0(n42345), .I1(n42902), .I2(n42794), 
            .I3(n42493), .O(n39598));
    defparam i3_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1081 (.I0(\data_in_frame[6] [4]), .I1(n42462), 
            .I2(Kp_23__N_1093), .I3(GND_net), .O(n27215));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1081.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27246));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_LUT4 i15205_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n28719));
    defparam i15205_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30706_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45837));
    defparam i30706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30707_4_lut (.I0(n45837), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n45838));
    defparam i30707_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i30705_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n45836));
    defparam i30705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2084076_i1_3_lut (.I0(n48673), .I1(n48781), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4522));
    defparam i2084076_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1083 (.I0(\data_in_frame[5] [0]), .I1(n42744), 
            .I2(\data_in_frame[7] [1]), .I3(GND_net), .O(n42430));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1083.LUT_INIT = 16'h9696;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(CLK_c), 
            .D(n41775), .S(n41689));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(CLK_c), 
            .D(n41773), .S(n43514));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(CLK_c), 
            .D(n7_adj_4523), .S(n8_adj_4524));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(CLK_c), 
            .D(n7_adj_4525), .S(n33842));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15206_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n28720));
    defparam i15206_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(CLK_c), 
            .D(n7_adj_4526), .S(n8_adj_4527));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(CLK_c), 
            .D(n41771), .S(n41693));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(CLK_c), 
            .D(n7_adj_4528), .S(n8_adj_4529));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(CLK_c), 
            .D(n7_adj_4530), .S(n8_adj_4531));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(CLK_c), 
            .D(n41769), .S(n41695));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(CLK_c), 
            .D(n41767), .S(n41697));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(CLK_c), 
            .D(n41765), .S(n41699));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(CLK_c), 
            .D(n41763), .S(n41701));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(CLK_c), 
            .D(n41761), .S(n41703));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(CLK_c), 
            .D(n41759), .S(n41667));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(CLK_c), 
            .D(n41757), .S(n41705));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(CLK_c), 
            .D(n41755), .S(n41707));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(CLK_c), 
            .D(n33222), .S(n41709));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(CLK_c), 
            .D(n41753), .S(n41711));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(CLK_c), 
            .D(n41751), .S(n41663));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(CLK_c), 
            .D(n41749), .S(n41713));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(CLK_c), 
            .D(n41747), .S(n41715));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1084 (.I0(\data_in_frame[5] [6]), .I1(n26855), 
            .I2(Kp_23__N_1064), .I3(n6_adj_4532), .O(n40494));
    defparam i4_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1085 (.I0(\data_in_frame[8] [2]), .I1(n27246), 
            .I2(n42410), .I3(n42748), .O(n26784));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_in_frame[8] [0]), .I1(n40494), 
            .I2(GND_net), .I3(GND_net), .O(n40566));
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(CLK_c), 
            .D(n41745), .S(n41717));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(CLK_c), 
            .D(n41743), .S(n41719));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(CLK_c), 
            .D(n41741), .S(n41721));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(CLK_c), 
            .D(n33220), .S(n8_adj_4533));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(CLK_c), 
            .D(n41739), .S(n41657));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n41661), .S(n10_adj_4534));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state_c [1]), .C(CLK_c), 
            .D(n41655), .S(n48857));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15207_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n28721));
    defparam i15207_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1087 (.I0(\data_in_frame[6] [7]), .I1(n42763), 
            .I2(n42430), .I3(\data_in_frame[4] [5]), .O(n27196));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i15208_3_lut_4_lut (.I0(n10_adj_4515), .I1(n42254), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n28722));
    defparam i15208_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1088 (.I0(n42354), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(n42717), .O(n10_adj_4535));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1089 (.I0(\data_in_frame[4] [0]), .I1(n10_adj_4535), 
            .I2(\data_in_frame[1] [4]), .I3(GND_net), .O(Kp_23__N_1090));   // verilog/coms.v(78[16:27])
    defparam i5_3_lut_adj_1089.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1090 (.I0(n42319), .I1(n42705), .I2(\data_in_frame[1] [6]), 
            .I3(GND_net), .O(Kp_23__N_936));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1090.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1091 (.I0(\data_in_frame[5] [3]), .I1(n26968), 
            .I2(GND_net), .I3(GND_net), .O(n42493));
    defparam i1_2_lut_adj_1091.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_in_frame[5] [1]), .I1(n42744), 
            .I2(GND_net), .I3(GND_net), .O(n42465));
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1093 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42782));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1094 (.I0(n26643), .I1(\data_in_frame[7] [6]), 
            .I2(n26855), .I3(GND_net), .O(n26801));
    defparam i2_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1095 (.I0(n42493), .I1(\data_in_frame[5] [2]), 
            .I2(\data_in_frame[7] [4]), .I3(n42658), .O(n10_adj_4536));
    defparam i4_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1096 (.I0(n27289), .I1(n10_adj_4536), .I2(n4_adj_4537), 
            .I3(GND_net), .O(n26809));
    defparam i5_3_lut_adj_1096.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1097 (.I0(n26968), .I1(n42782), .I2(\data_in_frame[0] [7]), 
            .I3(Kp_23__N_988), .O(n6_adj_4538));   // verilog/coms.v(85[17:70])
    defparam i1_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1098 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[4] [7]), 
            .I2(n42465), .I3(n6_adj_4538), .O(n39554));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i31892_2_lut (.I0(n48817), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n46828));
    defparam i31892_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i4_4_lut_adj_1099 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[4] [3]), .I3(n6_adj_4539), .O(Kp_23__N_1099));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i32336_3_lut (.I0(n48667), .I1(n48841), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n47468));
    defparam i32336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1100 (.I0(\data_in_frame[2] [0]), .I1(n42545), 
            .I2(Kp_23__N_993), .I3(n27125), .O(Kp_23__N_1096));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1101 (.I0(Kp_23__N_1096), .I1(Kp_23__N_1099), .I2(GND_net), 
            .I3(GND_net), .O(n42766));
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1102 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42389));
    defparam i1_2_lut_adj_1102.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1103 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4540));   // verilog/coms.v(85[17:63])
    defparam i2_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1104 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42376));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1064));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1105 (.I0(n26855), .I1(\data_in_frame[1] [4]), 
            .I2(n42376), .I3(\data_in_frame[5] [6]), .O(n42410));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1106 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42717));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1106.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42805));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42449));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(CLK_c), 
            .E(n27701), .D(n8825[0]), .R(n28149));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(CLK_c), .E(n43203), .D(n6958), 
            .R(n4_adj_4541));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n42512));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42364));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42337));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1112 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42354));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1112.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1113 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(n42325), .I3(n6_adj_4542), .O(Kp_23__N_969));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42325));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_993));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1115 (.I0(\data_in_frame[1] [4]), .I1(n42962), 
            .I2(GND_net), .I3(GND_net), .O(n42345));
    defparam i1_2_lut_adj_1115.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33629 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n48796));
    defparam byte_transmit_counter_0__bdd_4_lut_33629.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1116 (.I0(n42899), .I1(n42313), .I2(\data_out_frame[10] [0]), 
            .I3(n42959), .O(n10_adj_4543));
    defparam i4_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n26713));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42794));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42779));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1120 (.I0(n42726), .I1(n10_adj_4543), .I2(n7_adj_4540), 
            .I3(n8_adj_4544), .O(n40492));
    defparam i5_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1121 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_988), .I3(\data_in_frame[0] [5]), .O(n26968));
    defparam i1_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1122 (.I0(\data_in_frame[5] [4]), .I1(n42658), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n26643));
    defparam i2_3_lut_adj_1122.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1123 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42545));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1123.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1124 (.I0(n26965), .I1(\data_out_frame[4] [7]), 
            .I2(n1168), .I3(GND_net), .O(n26097));   // verilog/coms.v(71[16:69])
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1125 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[12] [3]), .I3(\data_out_frame[12] [1]), 
            .O(n12_adj_4545));
    defparam i5_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n28270));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_1126 (.I0(n42711), .I1(n26968), .I2(n42328), 
            .I3(n42779), .O(n32_adj_4546));   // verilog/coms.v(78[16:27])
    defparam i12_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1127 (.I0(n42763), .I1(n32_adj_4546), .I2(n22_adj_4547), 
            .I3(\data_in_frame[5] [1]), .O(n36_adj_4548));   // verilog/coms.v(78[16:27])
    defparam i16_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1128 (.I0(\data_in_frame[4] [4]), .I1(n27133), 
            .I2(\data_in_frame[5] [2]), .I3(n42407), .O(n34_adj_4549));   // verilog/coms.v(78[16:27])
    defparam i14_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n28269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n28268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n28267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n28266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n28265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n28264));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n28263));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_1129 (.I0(Kp_23__N_969), .I1(n42354), .I2(n42744), 
            .I3(\data_in_frame[2] [1]), .O(n35_adj_4550));   // verilog/coms.v(78[16:27])
    defparam i15_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1130 (.I0(\data_out_frame[12] [2]), .I1(n12_adj_4545), 
            .I2(\data_out_frame[6] [3]), .I3(n26527), .O(n42509));
    defparam i6_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n28262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n28261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n28260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n28259));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n28258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n28257));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n28256));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1131 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4551));
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_1132 (.I0(n42717), .I1(n42410), .I2(n42705), 
            .I3(n26713), .O(n33_adj_4552));   // verilog/coms.v(78[16:27])
    defparam i13_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n33_adj_4552), .I1(n35_adj_4550), .I2(n34_adj_4549), 
            .I3(n36_adj_4548), .O(n39558));   // verilog/coms.v(78[16:27])
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1133 (.I0(\data_out_frame[7] [1]), .I1(n42757), 
            .I2(n26097), .I3(n6_adj_4551), .O(n39567));
    defparam i4_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(\data_in_frame[8] [1]), .I1(n39558), 
            .I2(GND_net), .I3(GND_net), .O(n39596));
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1135 (.I0(\data_in_frame[4] [5]), .I1(\data_in_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4553));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n28255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n28254));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n28253));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1136 (.I0(n42512), .I1(n42449), .I2(n42805), 
            .I3(n6_adj_4553), .O(n42436));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1137 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[16] [4]), .I3(GND_net), .O(n26531));
    defparam i2_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1138 (.I0(Kp_23__N_993), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[1] [5]), .I3(n42364), .O(n10_adj_4554));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1139 (.I0(\data_in_frame[3] [7]), .I1(n10_adj_4554), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(Kp_23__N_1093));   // verilog/coms.v(73[16:42])
    defparam i5_3_lut_adj_1139.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1140 (.I0(n27401), .I1(Kp_23__N_1093), .I2(n42436), 
            .I3(n39596), .O(n12_adj_4555));
    defparam i5_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1141 (.I0(Kp_23__N_936), .I1(n12_adj_4555), .I2(n42766), 
            .I3(Kp_23__N_1090), .O(n44557));
    defparam i6_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 equal_2186_i7_2_lut (.I0(Kp_23__N_1195), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4556));   // verilog/coms.v(236[9:81])
    defparam equal_2186_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i12_4_lut_adj_1142 (.I0(n39554), .I1(n26809), .I2(n44557), 
            .I3(n26801), .O(n28_adj_4557));
    defparam i12_4_lut_adj_1142.LUT_INIT = 16'hf7ff;
    SB_LUT4 i5_3_lut_adj_1143 (.I0(n39567), .I1(\data_out_frame[8] [4]), 
            .I2(n42509), .I3(GND_net), .O(n14_adj_4558));
    defparam i5_3_lut_adj_1143.LUT_INIT = 16'h9696;
    SB_LUT4 n48796_bdd_4_lut (.I0(n48796), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n48799));
    defparam n48796_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33624 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27][0] ), 
            .I3(byte_transmit_counter[1]), .O(n48790));
    defparam byte_transmit_counter_0__bdd_4_lut_33624.LUT_INIT = 16'he4aa;
    SB_LUT4 n48790_bdd_4_lut (.I0(n48790), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n48793));
    defparam n48790_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1144 (.I0(n42808), .I1(\data_out_frame[12] [0]), 
            .I2(n40492), .I3(n42693), .O(n15_adj_4559));
    defparam i6_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n28252));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i10_4_lut_adj_1145 (.I0(n26789), .I1(n27196), .I2(n40566), 
            .I3(n26784), .O(n26_adj_4560));
    defparam i10_4_lut_adj_1145.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1146 (.I0(n27215), .I1(n5), .I2(n39598), .I3(n7_adj_4556), 
            .O(n27_adj_4561));
    defparam i11_4_lut_adj_1146.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1147 (.I0(n27203), .I1(n26756), .I2(n42685), 
            .I3(n8_adj_4447), .O(n25_adj_4562));
    defparam i9_4_lut_adj_1147.LUT_INIT = 16'hffef;
    SB_LUT4 i15_4_lut_adj_1148 (.I0(n25_adj_4562), .I1(n27_adj_4561), .I2(n26_adj_4560), 
            .I3(n28_adj_4557), .O(n31_adj_4452));
    defparam i15_4_lut_adj_1148.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1149 (.I0(n15_adj_4559), .I1(\data_out_frame[4] [1]), 
            .I2(n14_adj_4558), .I3(\data_out_frame[4] [2]), .O(n43705));
    defparam i8_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(CLK_c), 
            .D(n2_adj_4563), .S(n3_adj_4564));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i12_4_lut_adj_1150 (.I0(\data_out_frame[8] [0]), .I1(n27027), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[6] [2]), .O(n28_adj_4565));
    defparam i12_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1151 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4566));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_1151.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut_adj_1152 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4567));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_1152.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_1153 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4568));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_1153.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1154 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_4569));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_1154.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1155 (.I0(n9_adj_4569), .I1(n11_adj_4568), .I2(n10_adj_4567), 
            .I3(n12_adj_4566), .O(n23788));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1155.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1156 (.I0(n42439), .I1(n42316), .I2(\data_out_frame[13] [7]), 
            .I3(n42726), .O(n26_adj_4570));
    defparam i10_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1157 (.I0(n42496), .I1(n42723), .I2(n42738), 
            .I3(n43705), .O(n27_adj_4571));
    defparam i11_4_lut_adj_1157.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1158 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(n42760), .I3(n42509), .O(n25_adj_4572));
    defparam i9_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1159 (.I0(\FRAME_MATCHER.state [0]), .I1(n23788), 
            .I2(GND_net), .I3(GND_net), .O(n42248));
    defparam i1_2_lut_adj_1159.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1160 (.I0(n25_adj_4572), .I1(n27_adj_4571), .I2(n26_adj_4570), 
            .I3(n28_adj_4565), .O(n42293));
    defparam i15_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 n48826_bdd_4_lut (.I0(n48826), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n48829));
    defparam n48826_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i33270_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n7_c), .I2(\FRAME_MATCHER.state_c [2]), 
            .I3(n33839), .O(n27685));
    defparam i33270_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i2_3_lut_4_lut_adj_1161 (.I0(n26661), .I1(n27133), .I2(n42436), 
            .I3(\data_in_frame[6] [0]), .O(n27588));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 mux_2022_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n7001), .I3(GND_net), .O(n7002));
    defparam mux_2022_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1162 (.I0(n26661), .I1(n27133), .I2(\data_in_frame[4] [7]), 
            .I3(GND_net), .O(n42763));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1162.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1163 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n27125));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1163.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1164 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n27133));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1165 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n4_adj_4537));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_1165.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_969), 
            .I2(GND_net), .I3(GND_net), .O(n42442));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1167 (.I0(\data_out_frame[20] [2]), .I1(n42675), 
            .I2(n42537), .I3(\data_out_frame[24] [4]), .O(n42887));
    defparam i3_4_lut_adj_1167.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1168 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42340));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1169 (.I0(\FRAME_MATCHER.state_c [29]), .I1(\FRAME_MATCHER.state_c [26]), 
            .I2(\FRAME_MATCHER.state_c [19]), .I3(\FRAME_MATCHER.state_c [11]), 
            .O(n28_adj_4573));   // verilog/coms.v(212[5:16])
    defparam i10_4_lut_adj_1169.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1170 (.I0(\FRAME_MATCHER.state_c [31]), .I1(\FRAME_MATCHER.state_c [21]), 
            .I2(\FRAME_MATCHER.state_c [24]), .I3(\FRAME_MATCHER.state_c [15]), 
            .O(n31_adj_4574));   // verilog/coms.v(212[5:16])
    defparam i13_4_lut_adj_1170.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1171 (.I0(\FRAME_MATCHER.state_c [25]), .I1(\FRAME_MATCHER.state_c [28]), 
            .I2(\FRAME_MATCHER.state_c [14]), .I3(\FRAME_MATCHER.state_c [10]), 
            .O(n10_adj_4575));
    defparam i4_4_lut_adj_1171.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1172 (.I0(\data_out_frame[20] [1]), .I1(n42426), 
            .I2(\data_out_frame[19] [6]), .I3(\data_out_frame[22] [2]), 
            .O(n42953));
    defparam i3_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1173 (.I0(\data_out_frame[22] [4]), .I1(n42953), 
            .I2(n42947), .I3(n42887), .O(n43569));
    defparam i3_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33619 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n48778));
    defparam byte_transmit_counter_0__bdd_4_lut_33619.LUT_INIT = 16'he4aa;
    SB_LUT4 n48778_bdd_4_lut (.I0(n48778), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n48781));
    defparam n48778_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33609 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(byte_transmit_counter[1]), .O(n48772));
    defparam byte_transmit_counter_0__bdd_4_lut_33609.LUT_INIT = 16'he4aa;
    SB_LUT4 n48772_bdd_4_lut (.I0(n48772), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(byte_transmit_counter[1]), 
            .O(n48775));
    defparam n48772_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33604 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n48766));
    defparam byte_transmit_counter_0__bdd_4_lut_33604.LUT_INIT = 16'he4aa;
    SB_LUT4 n48766_bdd_4_lut (.I0(n48766), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n48769));
    defparam n48766_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33599 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n48760));
    defparam byte_transmit_counter_0__bdd_4_lut_33599.LUT_INIT = 16'he4aa;
    SB_LUT4 n48760_bdd_4_lut (.I0(n48760), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n48763));
    defparam n48760_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33594 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n48754));
    defparam byte_transmit_counter_0__bdd_4_lut_33594.LUT_INIT = 16'he4aa;
    SB_LUT4 n48754_bdd_4_lut (.I0(n48754), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n48757));
    defparam n48754_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33589 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n48748));
    defparam byte_transmit_counter_0__bdd_4_lut_33589.LUT_INIT = 16'he4aa;
    SB_LUT4 n48748_bdd_4_lut (.I0(n48748), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n48751));
    defparam n48748_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33584 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(byte_transmit_counter[1]), .O(n48742));
    defparam byte_transmit_counter_0__bdd_4_lut_33584.LUT_INIT = 16'he4aa;
    SB_LUT4 n48742_bdd_4_lut (.I0(n48742), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(byte_transmit_counter[1]), 
            .O(n48745));
    defparam n48742_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33579 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n48736));
    defparam byte_transmit_counter_0__bdd_4_lut_33579.LUT_INIT = 16'he4aa;
    SB_LUT4 n48736_bdd_4_lut (.I0(n48736), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n48739));
    defparam n48736_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4576), .S(n3_adj_4440));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4577), .S(n3_adj_4439));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4578), .S(n3_adj_4435));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n41301), .S(n3_adj_4434));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n41307), .S(n3_adj_4432));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n41309), .S(n3_adj_4430));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1174 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n26748));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1175 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(n1168), .I3(\data_out_frame[4] [5]), .O(n26965));
    defparam i1_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42392));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1177 (.I0(\data_out_frame[6] [3]), .I1(n42518), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n27188));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1177.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42878));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_out_frame[9] [1]), .I1(n27188), 
            .I2(GND_net), .I3(GND_net), .O(n42911));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1180 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42305));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1180.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1181 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n42732));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1182 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n42817));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1182.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1183 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n42379));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1183.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42357));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1185 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42838));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1185.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1186 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n42452));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_adj_1186.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1187 (.I0(\data_out_frame[5] [5]), .I1(n42487), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[5] [3]), .O(n1168));   // verilog/coms.v(71[16:62])
    defparam i3_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1188 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n42413));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1188.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1189 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n42529));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1189.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n41315), .S(n3_adj_4429));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n41321), .S(n3_adj_4428));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n41327), .S(n3_adj_4427));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n41349), .S(n3_adj_4425));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i17_4_lut (.I0(n42529), .I1(n27257), .I2(n42413), .I3(\data_out_frame[8] [0]), 
            .O(n42));   // verilog/coms.v(73[16:42])
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4564));
    defparam select_658_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1190 (.I0(\FRAME_MATCHER.state_c [17]), .I1(\FRAME_MATCHER.state_c [12]), 
            .I2(\FRAME_MATCHER.state_c [8]), .I3(\FRAME_MATCHER.state_c [16]), 
            .O(n30));   // verilog/coms.v(212[5:16])
    defparam i12_4_lut_adj_1190.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1191 (.I0(n31_adj_4574), .I1(\FRAME_MATCHER.state_c [18]), 
            .I2(n28_adj_4573), .I3(\FRAME_MATCHER.state_c [22]), .O(n34_adj_4579));   // verilog/coms.v(212[5:16])
    defparam i16_4_lut_adj_1191.LUT_INIT = 16'hfffe;
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n41365), .S(n3_adj_4423));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n41385), .S(n3_adj_4419));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_1192 (.I0(n42357), .I1(n42379), .I2(\data_out_frame[9] [3]), 
            .I3(n42817), .O(n40_adj_4580));   // verilog/coms.v(73[16:42])
    defparam i15_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1193 (.I0(n26553), .I1(\data_out_frame[6] [3]), 
            .I2(n42487), .I3(n42838), .O(n41));   // verilog/coms.v(73[16:42])
    defparam i16_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1194 (.I0(n42911), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[9] [4]), .I3(n42878), .O(n39_adj_4581));   // verilog/coms.v(73[16:42])
    defparam i14_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(n39_adj_4581), .I1(n41), .I2(n40_adj_4580), 
            .I3(n42), .O(n48));   // verilog/coms.v(73[16:42])
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1195 (.I0(n42392), .I1(\data_out_frame[6] [6]), 
            .I2(n42814), .I3(n26965), .O(n43));   // verilog/coms.v(73[16:42])
    defparam i18_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n43), .I1(n48), .I2(n37_adj_4582), .I3(n38_adj_4583), 
            .O(n40476));   // verilog/coms.v(73[16:42])
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_out_frame[11] [7]), .I1(n40476), 
            .I2(GND_net), .I3(GND_net), .O(n42899));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1197 (.I0(\data_out_frame[10] [0]), .I1(n40476), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n42723));
    defparam i2_3_lut_adj_1197.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1198 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n14_adj_4584));
    defparam i5_3_lut_adj_1198.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1199 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[9] [7]), 
            .I2(n42723), .I3(n42899), .O(n15_adj_4585));
    defparam i6_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1200 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n10_adj_4575), 
            .I2(\FRAME_MATCHER.state_c [13]), .I3(GND_net), .O(n40334));
    defparam i5_3_lut_adj_1200.LUT_INIT = 16'hfefe;
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n41405), .S(n3_adj_4418));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n41425), .S(n3_adj_4416));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n41445), .S(n3_adj_4415));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19788_3_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(n63), .I2(n63_adj_4586), 
            .I3(GND_net), .O(n122));   // verilog/coms.v(139[4] 141[7])
    defparam i19788_3_lut.LUT_INIT = 16'hb3b3;
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n41477), .S(n3_adj_4413));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11_4_lut_adj_1201 (.I0(\FRAME_MATCHER.state_c [20]), .I1(\FRAME_MATCHER.state_c [23]), 
            .I2(\FRAME_MATCHER.state_c [27]), .I3(\FRAME_MATCHER.state_c [30]), 
            .O(n29_adj_4587));   // verilog/coms.v(212[5:16])
    defparam i11_4_lut_adj_1201.LUT_INIT = 16'hfffe;
    SB_LUT4 select_686_Select_2_i7_3_lut (.I0(\FRAME_MATCHER.state_31__N_2660[2] ), 
            .I1(n26494), .I2(n4452), .I3(GND_net), .O(n7));
    defparam select_686_Select_2_i7_3_lut.LUT_INIT = 16'h3232;
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n41505), .S(n3_adj_4412));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19764_2_lut (.I0(\FRAME_MATCHER.state_31__N_2660[2] ), .I1(n3303), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2788[2] ));   // verilog/coms.v(227[6] 229[9])
    defparam i19764_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1202 (.I0(\FRAME_MATCHER.state_c [4]), .I1(\FRAME_MATCHER.state_c [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4589));
    defparam i2_2_lut_adj_1202.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1203 (.I0(n29_adj_4587), .I1(n40334), .I2(n34_adj_4579), 
            .I3(n30), .O(n4_adj_4590));   // verilog/coms.v(212[5:16])
    defparam i1_4_lut_adj_1203.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1204 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n4_adj_4590), 
            .I2(n6_adj_4589), .I3(\FRAME_MATCHER.state_c [6]), .O(n33839));   // verilog/coms.v(212[5:16])
    defparam i2_4_lut_adj_1204.LUT_INIT = 16'hfffe;
    SB_LUT4 select_658_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4591));
    defparam select_658_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33574 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n48730));
    defparam byte_transmit_counter_0__bdd_4_lut_33574.LUT_INIT = 16'he4aa;
    SB_LUT4 n48730_bdd_4_lut (.I0(n48730), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n48733));
    defparam n48730_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15185_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n28699));
    defparam i15185_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33569 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n48700));
    defparam byte_transmit_counter_0__bdd_4_lut_33569.LUT_INIT = 16'he4aa;
    SB_LUT4 n48700_bdd_4_lut (.I0(n48700), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n48703));
    defparam n48700_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33545 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n48694));
    defparam byte_transmit_counter_0__bdd_4_lut_33545.LUT_INIT = 16'he4aa;
    SB_LUT4 n48694_bdd_4_lut (.I0(n48694), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n48697));
    defparam n48694_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33540 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n48688));
    defparam byte_transmit_counter_0__bdd_4_lut_33540.LUT_INIT = 16'he4aa;
    SB_LUT4 n48688_bdd_4_lut (.I0(n48688), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n48691));
    defparam n48688_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15186_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n28700));
    defparam i15186_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1205 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_969), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[2] [1]), .O(n23_adj_4593));
    defparam i6_4_lut_adj_1205.LUT_INIT = 16'h2184;
    SB_LUT4 i9_3_lut (.I0(n23788), .I1(\data_in_frame[1] [4]), .I2(\data_in_frame[1] [5]), 
            .I3(GND_net), .O(n26_adj_4594));
    defparam i9_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i12_4_lut_adj_1206 (.I0(n23_adj_4593), .I1(n26661), .I2(\data_in_frame[2] [7]), 
            .I3(n42337), .O(n29_adj_4595));
    defparam i12_4_lut_adj_1206.LUT_INIT = 16'h2002;
    SB_LUT4 i5_4_lut_adj_1207 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n42340), .I3(n42442), .O(n22_adj_4596));
    defparam i5_4_lut_adj_1207.LUT_INIT = 16'h1248;
    SB_LUT4 i15187_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n28701));
    defparam i15187_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n41525), .S(n3_adj_4406));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n41547), .S(n3_adj_4405));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30668_3_lut (.I0(n4_adj_4537), .I1(\data_in_frame[2] [0]), 
            .I2(n42442), .I3(GND_net), .O(n45700));
    defparam i30668_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i15188_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n28702));
    defparam i15188_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15189_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n28703));
    defparam i15189_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1208 (.I0(n15_adj_4585), .I1(n42379), .I2(n14_adj_4584), 
            .I3(n24129), .O(n42616));
    defparam i8_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n41567), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33535 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n48682));
    defparam byte_transmit_counter_0__bdd_4_lut_33535.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_adj_1209 (.I0(n43197), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n33873), .I3(GND_net), .O(n26421));
    defparam i1_3_lut_adj_1209.LUT_INIT = 16'haeae;
    SB_LUT4 n48682_bdd_4_lut (.I0(n48682), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n48685));
    defparam n48682_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n41587), .S(n3_adj_4597));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33092_4_lut (.I0(n26421), .I1(n33873), .I2(n5_adj_4598), 
            .I3(n6_adj_4599), .O(n42196));
    defparam i33092_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33530 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n48676));
    defparam byte_transmit_counter_0__bdd_4_lut_33530.LUT_INIT = 16'he4aa;
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n41615), .S(n3_adj_4600));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n41641), .S(n3_adj_4601));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4602), .S(n3_adj_4603));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n28251));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_adj_1210 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_c));
    defparam i2_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n28783));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n28782));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n28781));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n28780));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n28779));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n28778));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n28777));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n28776));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n28775));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n28774));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n28773));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n28772));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n28771));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n28770));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n28769));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n28768));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n28767));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n28766));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n28765));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n28764));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n28763));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n28762));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n28761));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n28760));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n28759));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n28758));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n28757));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n28756));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n28755));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n28754));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n28250));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n28249));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n28248));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n28247));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n28246));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n28245));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n28244));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n28243));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n28242));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n28241));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n28240));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n28239));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n28238));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n28237));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n28236));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n28234));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n28233));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n28232));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n28226));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n28225));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n28224));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n28223));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n28222));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n28221));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(CLK_c), 
           .D(n41665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n28219));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n28218));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15190_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n28704));
    defparam i15190_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(CLK_c), .E(n42196), .D(n27964), 
            .R(n43482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n28217));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n28216));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4604), .S(n3_adj_4591));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15191_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n28705));
    defparam i15191_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n28753));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n28752));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n28751));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n28750));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n28749));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n28748));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n28747));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_1211 (.I0(n29_adj_4595), .I1(n26646), .I2(n26_adj_4594), 
            .I3(n27125), .O(n32_adj_4605));
    defparam i15_4_lut_adj_1211.LUT_INIT = 16'h0020;
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n28215));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n28214));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n28213));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n28212));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n28211));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n28210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n28209));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n28208));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n28207));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n28206));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n28205));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n28204));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n28202));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n28746));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48676_bdd_4_lut (.I0(n48676), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n48679));
    defparam n48676_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n28745));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n28744));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n28743));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n28742));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n28741));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n28740));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i10_4_lut_adj_1212 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [6]), 
            .I2(n27133), .I3(\data_in_frame[1] [2]), .O(n27_adj_4606));
    defparam i10_4_lut_adj_1212.LUT_INIT = 16'h0800;
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n28739));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1213 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n42395));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n28738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n28737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n28736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n28735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n28734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n28733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n28732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n28731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n28730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n28729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n28728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n28727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n28726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n28725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n28724));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n28723));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n28722));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n28721));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26539));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i15192_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42260), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n28706));
    defparam i15192_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n28720));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33525 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n48670));
    defparam byte_transmit_counter_0__bdd_4_lut_33525.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n28719));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48670_bdd_4_lut (.I0(n48670), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n48673));
    defparam n48670_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n28718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n28717));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33520 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(byte_transmit_counter[1]), .O(n48664));
    defparam byte_transmit_counter_0__bdd_4_lut_33520.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n28716));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48664_bdd_4_lut (.I0(n48664), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(byte_transmit_counter[1]), 
            .O(n48667));
    defparam n48664_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n28715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n28714));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n47468), .I2(n46828), .I3(byte_transmit_counter[4]), .O(n48658));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n28713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n28712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n28711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n28710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n28709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n28708));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n28707));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n28706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n28705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n28704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n28703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n28702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n28701));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n28700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n28699));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n28698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n28697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n28696));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n28695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n28694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n28693));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48658_bdd_4_lut (.I0(n48658), .I1(n14_adj_4522), .I2(n7_adj_4607), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n48658_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33510 (.I0(byte_transmit_counter[3]), 
            .I1(n47464), .I2(n46847), .I3(byte_transmit_counter[4]), .O(n48652));
    defparam byte_transmit_counter_3__bdd_4_lut_33510.LUT_INIT = 16'he4aa;
    SB_LUT4 n48652_bdd_4_lut (.I0(n48652), .I1(n14_adj_4521), .I2(n7_adj_4608), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n48652_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n28680));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4609), .S(n3_adj_4517));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4610), .S(n3_adj_4516));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1215 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(\data_out_frame[7] [5]), .O(n42496));
    defparam i3_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1216 (.I0(n42395), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[12] [2]), .I3(n42735), .O(n10_adj_4611));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_4612), .S(n3_adj_4504));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33515 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n48646));
    defparam byte_transmit_counter_0__bdd_4_lut_33515.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n28679));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n28678));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n28677));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4613), .S(n3_adj_4503));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n48646_bdd_4_lut (.I0(n48646), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n48649));
    defparam n48646_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n28676));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4614), .S(n3_adj_4500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n28169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n28168));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n27685), .D(n7025));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n27685), .D(n7024));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n27685), .D(n7023));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n27685), .D(n7022));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n27685), .D(n7021));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n27685), .D(n7020));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n27685), .D(n7019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n27685), .D(n7018));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n27685), .D(n7017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i217 (.Q(\data_out_frame[27][0] ), .C(CLK_c), 
           .D(n28166));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n27685), .D(n7016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n28164));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n27685), .D(n7015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n27685), .D(n7014));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n27685), .D(n7013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n27685), .D(n7012));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n27685), .D(n7011));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n27685), .D(n7010));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n27685), .D(n7009));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n27685), .D(n7008));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n27685), .D(n7007));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n27685), .D(n7006));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n27685), .D(n7005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n27685), .D(n7004));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n27685), .D(n7003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n28163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n28162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n28161));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33505 (.I0(byte_transmit_counter[3]), 
            .I1(n47462), .I2(n46829), .I3(byte_transmit_counter[4]), .O(n48640));
    defparam byte_transmit_counter_3__bdd_4_lut_33505.LUT_INIT = 16'he4aa;
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n28160));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i16_4_lut_adj_1217 (.I0(n27_adj_4606), .I1(n32_adj_4605), .I2(n45700), 
            .I3(n22_adj_4596), .O(\FRAME_MATCHER.state_31__N_2724 [3]));
    defparam i16_4_lut_adj_1217.LUT_INIT = 16'h0800;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1218 (.I0(n33239), .I1(n10_adj_4515), .I2(GND_net), 
            .I3(GND_net), .O(n42281));
    defparam i1_2_lut_adj_1218.LUT_INIT = 16'hdddd;
    SB_LUT4 i5_4_lut_adj_1219 (.I0(\data_out_frame[7] [7]), .I1(n42496), 
            .I2(\data_out_frame[5] [7]), .I3(n26539), .O(n12_adj_4615));
    defparam i5_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[22] [7]), .I1(n44481), .I2(n40258), 
            .I3(GND_net), .O(n10_adj_4616));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1220 (.I0(\data_out_frame[22] [7]), .I1(n44481), 
            .I2(n39625), .I3(GND_net), .O(n6_adj_4617));
    defparam i1_2_lut_3_lut_adj_1220.LUT_INIT = 16'h6969;
    SB_LUT4 n48640_bdd_4_lut (.I0(n48640), .I1(n14_adj_4431), .I2(n7_adj_4618), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n48640_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1221 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [4]), .I3(GND_net), .O(n41739));
    defparam i1_2_lut_3_lut_adj_1221.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33664 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [4]), .I2(\data_out_frame[23] [4]), 
            .I3(byte_transmit_counter[1]), .O(n48838));
    defparam byte_transmit_counter_0__bdd_4_lut_33664.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1222 (.I0(n33239), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n42274));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1222.LUT_INIT = 16'hffdf;
    SB_LUT4 i19724_2_lut_3_lut (.I0(n1_adj_4619), .I1(n3_adj_4620), .I2(\FRAME_MATCHER.state_c [5]), 
            .I3(GND_net), .O(n33220));
    defparam i19724_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_3_lut_adj_1223 (.I0(n39558), .I1(n27588), .I2(n27451), 
            .I3(GND_net), .O(n42685));
    defparam i2_2_lut_3_lut_adj_1223.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1224 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [6]), .I3(GND_net), .O(n41741));
    defparam i1_2_lut_3_lut_adj_1224.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n45905), .I2(n45906), .I3(byte_transmit_counter[2]), .O(n48634));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n28675));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1225 (.I0(\data_out_frame[5] [3]), .I1(n12_adj_4615), 
            .I2(\data_out_frame[12] [3]), .I3(\data_out_frame[9] [7]), .O(n42458));
    defparam i6_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1226 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [7]), .I3(GND_net), .O(n41743));
    defparam i1_2_lut_3_lut_adj_1226.LUT_INIT = 16'he0e0;
    SB_LUT4 n48634_bdd_4_lut (.I0(n48634), .I1(n45900), .I2(n45899), .I3(byte_transmit_counter[2]), 
            .O(n47460));
    defparam n48634_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n28673));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1227 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [8]), .I3(GND_net), .O(n41745));
    defparam i1_2_lut_3_lut_adj_1227.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1228 (.I0(n39558), .I1(n27588), .I2(\data_in_frame[3] [5]), 
            .I3(GND_net), .O(n6_adj_4532));
    defparam i1_2_lut_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [9]), .I3(GND_net), .O(n41747));
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1230 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [10]), .I3(GND_net), .O(n41749));
    defparam i1_2_lut_3_lut_adj_1230.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1231 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [11]), .I3(GND_net), .O(n41751));
    defparam i1_2_lut_3_lut_adj_1231.LUT_INIT = 16'he0e0;
    SB_LUT4 i15165_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n28679));
    defparam i15165_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1232 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [12]), .I3(GND_net), .O(n41753));
    defparam i1_2_lut_3_lut_adj_1232.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n28672));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1233 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n19799));   // verilog/coms.v(214[11:56])
    defparam i2_3_lut_adj_1233.LUT_INIT = 16'hfefe;
    SB_LUT4 i19725_2_lut_3_lut (.I0(n1_adj_4619), .I1(n3_adj_4620), .I2(\FRAME_MATCHER.state_c [13]), 
            .I3(GND_net), .O(n33222));
    defparam i19725_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i20325_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n33827));
    defparam i20325_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1234 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n33827), .I3(byte_transmit_counter[2]), .O(n34010));
    defparam i2_4_lut_adj_1234.LUT_INIT = 16'h8880;
    SB_LUT4 n48820_bdd_4_lut (.I0(n48820), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n48823));
    defparam n48820_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33644 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n48814));
    defparam byte_transmit_counter_0__bdd_4_lut_33644.LUT_INIT = 16'he4aa;
    SB_LUT4 n48814_bdd_4_lut (.I0(n48814), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n48817));
    defparam n48814_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33495 (.I0(byte_transmit_counter[3]), 
            .I1(n47460), .I2(n46834), .I3(byte_transmit_counter[4]), .O(n48628));
    defparam byte_transmit_counter_3__bdd_4_lut_33495.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33639 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n48808));
    defparam byte_transmit_counter_0__bdd_4_lut_33639.LUT_INIT = 16'he4aa;
    SB_LUT4 i3_4_lut_adj_1235 (.I0(n34010), .I1(n33639), .I2(n33209), 
            .I3(n19799), .O(n43918));
    defparam i3_4_lut_adj_1235.LUT_INIT = 16'hfffb;
    SB_LUT4 n48628_bdd_4_lut (.I0(n48628), .I1(n14_adj_4421), .I2(n7_adj_4622), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n48628_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1378_i1_3_lut (.I0(n43918), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n33873), .I3(GND_net), .O(n4888[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_1378_i1_3_lut.LUT_INIT = 16'h5c5c;
    SB_LUT4 i1_2_lut_3_lut_adj_1236 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [14]), .I3(GND_net), .O(n41755));
    defparam i1_2_lut_3_lut_adj_1236.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_33486 (.I0(byte_transmit_counter[3]), 
            .I1(n47458), .I2(n46849), .I3(byte_transmit_counter[4]), .O(n48622));
    defparam byte_transmit_counter_3__bdd_4_lut_33486.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1237 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [15]), .I3(GND_net), .O(n41757));
    defparam i1_2_lut_3_lut_adj_1237.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1238 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [16]), .I3(GND_net), .O(n41759));
    defparam i1_2_lut_3_lut_adj_1238.LUT_INIT = 16'he0e0;
    SB_LUT4 n48622_bdd_4_lut (.I0(n48622), .I1(n14_adj_4420), .I2(n7_adj_4623), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n48622_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15166_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n28680));
    defparam i15166_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1239 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [17]), .I3(GND_net), .O(n41761));
    defparam i1_2_lut_3_lut_adj_1239.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1240 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [18]), .I3(GND_net), .O(n41763));
    defparam i1_2_lut_3_lut_adj_1240.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33500 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n48610));
    defparam byte_transmit_counter_0__bdd_4_lut_33500.LUT_INIT = 16'he4aa;
    SB_LUT4 n48610_bdd_4_lut (.I0(n48610), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n48613));
    defparam n48610_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19803_2_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33300));
    defparam i19803_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33472 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n48604));
    defparam byte_transmit_counter_0__bdd_4_lut_33472.LUT_INIT = 16'he4aa;
    SB_LUT4 n48604_bdd_4_lut (.I0(n48604), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n48607));
    defparam n48604_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1241 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [19]), .I3(GND_net), .O(n41765));
    defparam i1_2_lut_3_lut_adj_1241.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1242 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [20]), .I3(GND_net), .O(n41767));
    defparam i1_2_lut_3_lut_adj_1242.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1243 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [21]), .I3(GND_net), .O(n41769));
    defparam i1_2_lut_3_lut_adj_1243.LUT_INIT = 16'he0e0;
    SB_LUT4 i15179_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n28693));
    defparam i15179_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1244 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [22]), .I3(GND_net), .O(n7_adj_4530));
    defparam i1_2_lut_3_lut_adj_1244.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1245 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [23]), .I3(GND_net), .O(n7_adj_4528));
    defparam i1_2_lut_3_lut_adj_1245.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [24]), .I3(GND_net), .O(n41771));
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1247 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [25]), .I3(GND_net), .O(n7_adj_4526));
    defparam i1_2_lut_3_lut_adj_1247.LUT_INIT = 16'he0e0;
    SB_LUT4 i15180_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n28694));
    defparam i15180_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33467 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n48592));
    defparam byte_transmit_counter_0__bdd_4_lut_33467.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1248 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [26]), .I3(GND_net), .O(n7_adj_4525));
    defparam i1_2_lut_3_lut_adj_1248.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1249 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [27]), .I3(GND_net), .O(n7_adj_4523));
    defparam i1_2_lut_3_lut_adj_1249.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1250 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [28]), .I3(GND_net), .O(n41773));
    defparam i1_2_lut_3_lut_adj_1250.LUT_INIT = 16'he0e0;
    SB_LUT4 i15181_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n28695));
    defparam i15181_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1251 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [29]), .I3(GND_net), .O(n41775));
    defparam i1_2_lut_3_lut_adj_1251.LUT_INIT = 16'he0e0;
    SB_LUT4 n48592_bdd_4_lut (.I0(n48592), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n48595));
    defparam n48592_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1252 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [30]), .I3(GND_net), .O(n41777));
    defparam i1_2_lut_3_lut_adj_1252.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1253 (.I0(n1_adj_4619), .I1(n3_adj_4620), 
            .I2(\FRAME_MATCHER.state_c [31]), .I3(GND_net), .O(n41737));
    defparam i1_2_lut_3_lut_adj_1253.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1254 (.I0(n42506), .I1(n42799), .I2(n27084), 
            .I3(n42884), .O(n4_adj_4624));
    defparam i1_2_lut_4_lut_adj_1254.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1255 (.I0(n42506), .I1(n42799), .I2(n27084), 
            .I3(\data_out_frame[19] [6]), .O(n27282));
    defparam i1_2_lut_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i15182_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n28696));
    defparam i15182_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33458 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n48586));
    defparam byte_transmit_counter_0__bdd_4_lut_33458.LUT_INIT = 16'he4aa;
    SB_LUT4 n48586_bdd_4_lut (.I0(n48586), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n48589));
    defparam n48586_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15183_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n28697));
    defparam i15183_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_658_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4603));
    defparam select_658_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1256 (.I0(n63), .I1(n63_adj_4586), 
            .I2(n7_adj_4625), .I3(n99), .O(n42235));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_4_lut_adj_1256.LUT_INIT = 16'h8880;
    SB_LUT4 i1_3_lut_4_lut (.I0(n63), .I1(n63_adj_4586), .I2(n126), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(\FRAME_MATCHER.state_31__N_2660 [1]));   // verilog/coms.v(139[7:80])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf8f0;
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(n63), .I1(n63_adj_4586), .I2(n126), 
            .I3(GND_net), .O(n23516));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'h0808;
    SB_LUT4 select_658_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4601));
    defparam select_658_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1258 (.I0(\data_out_frame[5] [4]), .I1(n42905), 
            .I2(\data_out_frame[12] [0]), .I3(n42616), .O(n12_adj_4626));
    defparam i5_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4600));
    defparam select_658_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_658_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4468));
    defparam select_658_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1259 (.I0(\data_out_frame[11] [7]), .I1(n12_adj_4626), 
            .I2(\data_out_frame[14] [2]), .I3(n42735), .O(n42689));
    defparam i6_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33453 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n48580));
    defparam byte_transmit_counter_0__bdd_4_lut_33453.LUT_INIT = 16'he4aa;
    SB_LUT4 i15184_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42260), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n28698));
    defparam i15184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n48580_bdd_4_lut (.I0(n48580), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n48583));
    defparam n48580_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n28159));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1260 (.I0(\data_in_frame[6] [2]), .I1(Kp_23__N_1090), 
            .I2(\data_in_frame[8] [3]), .I3(n42748), .O(n26789));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n37565), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n28158));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n37564), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_4_lut_adj_1261 (.I0(\data_in[2] [7]), .I1(n10_adj_4627), 
            .I2(\data_in[3] [4]), .I3(\data_in[1] [5]), .O(n12_adj_4628));
    defparam i1_2_lut_4_lut_adj_1261.LUT_INIT = 16'hffdf;
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n28671));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n28670));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in[2] [7]), .I1(n10_adj_4627), .I2(\data_in[3] [4]), 
            .I3(\data_in[2] [4]), .O(n7_adj_4629));
    defparam i2_2_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i3_4_lut_adj_1262 (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state_31__N_2724 [3]), 
            .I2(n23237), .I3(n33839), .O(n23622));
    defparam i3_4_lut_adj_1262.LUT_INIT = 16'h0080;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33448 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n48574));
    defparam byte_transmit_counter_0__bdd_4_lut_33448.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1263 (.I0(\data_in_frame[6] [2]), .I1(Kp_23__N_1090), 
            .I2(n26687), .I3(n27199), .O(n42593));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1264 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n33239), .O(n42254));
    defparam i2_3_lut_4_lut_adj_1264.LUT_INIT = 16'hf7ff;
    SB_LUT4 equal_2186_i5_2_lut_3_lut_4_lut (.I0(\data_in_frame[6] [2]), .I1(Kp_23__N_1090), 
            .I2(\data_in_frame[8] [4]), .I3(n27199), .O(n5));   // verilog/coms.v(74[16:43])
    defparam equal_2186_i5_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2898_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4630));
    defparam i2898_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1265 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42260), .I3(\FRAME_MATCHER.i [0]), .O(n42267));
    defparam i1_2_lut_3_lut_4_lut_adj_1265.LUT_INIT = 16'hf7ff;
    SB_LUT4 i32709_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n33873), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4541));
    defparam i32709_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45862), .I3(n45860), .O(n7_adj_4623));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i33425_4_lut (.I0(n43197), .I1(\FRAME_MATCHER.state [3]), .I2(n6958), 
            .I3(n33873), .O(n43203));
    defparam i33425_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45856), .I3(n45854), .O(n7_adj_4622));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i32755_2_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6958));   // verilog/coms.v(145[4] 299[11])
    defparam i32755_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1266 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42281), .I3(\FRAME_MATCHER.i [0]), .O(n42288));
    defparam i1_2_lut_3_lut_4_lut_adj_1266.LUT_INIT = 16'hf7ff;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[18] [0]), 
            .I2(n42627), .I3(n10_adj_4433), .O(n43617));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_CARRY add_3971_8 (.CI(n37564), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n37565));
    SB_LUT4 i2_3_lut_4_lut_adj_1267 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[18] [0]), 
            .I2(n27378), .I3(n42506), .O(n42426));
    defparam i2_3_lut_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45850), .I3(n45848), .O(n7_adj_4618));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n37563), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_7 (.CI(n37563), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n37564));
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n37562), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_6 (.CI(n37562), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n37563));
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n37561), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_5 (.CI(n37561), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n37562));
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n37560), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_4_lut_adj_1268 (.I0(n2_adj_4631), .I1(n1_adj_4632), 
            .I2(n1_adj_4619), .I3(\FRAME_MATCHER.state [3]), .O(n88));
    defparam i1_3_lut_4_lut_adj_1268.LUT_INIT = 16'hfe00;
    SB_CARRY add_3971_4 (.CI(n37560), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n37561));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n37559), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_3 (.CI(n37559), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n37560));
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3513), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 n48574_bdd_4_lut (.I0(n48574), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n48577));
    defparam n48574_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3513), 
            .CO(n37559));
    SB_LUT4 add_43_33_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [31]), 
            .I2(GND_net), .I3(n37558), .O(n2_adj_4563)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45832), .I3(n45830), .O(n7_adj_4508));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n28669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n28157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n28668));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n28667));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_32_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [30]), 
            .I2(GND_net), .I3(n37557), .O(n2_adj_4576)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n28666));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_32 (.CI(n37557), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n37558));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45826), .I3(n45824), .O(n7_adj_4511));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i32_3_lut_4_lut (.I0(n26912), .I1(n39506), .I2(n39574), .I3(n64), 
            .O(n74));
    defparam i32_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 equal_286_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4621));   // verilog/coms.v(154[7:23])
    defparam equal_286_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_2_lut_3_lut_adj_1269 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4592));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_adj_1269.LUT_INIT = 16'hfefe;
    SB_LUT4 add_43_31_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [29]), 
            .I2(GND_net), .I3(n37556), .O(n2_adj_4577)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n37556), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n37557));
    SB_LUT4 add_43_30_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [28]), 
            .I2(GND_net), .I3(n37555), .O(n2_adj_4578)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_30 (.CI(n37555), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n37556));
    SB_LUT4 add_43_29_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(n37554), .O(n41301)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_29 (.CI(n37554), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n37555));
    SB_LUT4 add_43_28_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [26]), 
            .I2(GND_net), .I3(n37553), .O(n41307)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_28 (.CI(n37553), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n37554));
    SB_LUT4 add_43_27_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [25]), 
            .I2(GND_net), .I3(n37552), .O(n41309)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_27 (.CI(n37552), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n37553));
    SB_LUT4 add_43_26_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [24]), 
            .I2(GND_net), .I3(n37551), .O(n41315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_26 (.CI(n37551), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n37552));
    SB_LUT4 add_43_25_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [23]), 
            .I2(GND_net), .I3(n37550), .O(n41321)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_25 (.CI(n37550), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n37551));
    SB_LUT4 add_43_24_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [22]), 
            .I2(GND_net), .I3(n37549), .O(n41327)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_24 (.CI(n37549), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n37550));
    SB_LUT4 add_43_23_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [21]), 
            .I2(GND_net), .I3(n37548), .O(n41349)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n37548), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n37549));
    SB_LUT4 add_43_22_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [20]), 
            .I2(GND_net), .I3(n37547), .O(n41365)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_22 (.CI(n37547), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n37548));
    SB_LUT4 add_43_21_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [19]), 
            .I2(GND_net), .I3(n37546), .O(n41385)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_21 (.CI(n37546), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n37547));
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33443 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n48568));
    defparam byte_transmit_counter_0__bdd_4_lut_33443.LUT_INIT = 16'he4aa;
    SB_LUT4 add_43_20_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [18]), 
            .I2(GND_net), .I3(n37545), .O(n41405)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n37545), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n37546));
    SB_LUT4 add_43_19_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [17]), 
            .I2(GND_net), .I3(n37544), .O(n41425)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_19 (.CI(n37544), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n37545));
    SB_LUT4 add_43_18_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [16]), 
            .I2(GND_net), .I3(n37543), .O(n41445)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n28665));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1270 (.I0(n44470), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n26495), .I3(n3813), .O(n42244));   // verilog/coms.v(157[9:60])
    defparam i1_3_lut_4_lut_adj_1270.LUT_INIT = 16'hff0d;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45838), .I3(n45836), .O(n7_adj_4607));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i2_4_lut_adj_1271 (.I0(\FRAME_MATCHER.state_31__N_2660 [1]), .I1(n3303), 
            .I2(n43094), .I3(n26482), .O(n6_adj_4634));
    defparam i2_4_lut_adj_1271.LUT_INIT = 16'h0aee;
    SB_CARRY add_43_18 (.CI(n37543), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n37544));
    SB_LUT4 i5_3_lut_4_lut_adj_1272 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [7]), 
            .I2(n10_adj_4635), .I3(n42576), .O(n44481));
    defparam i5_3_lut_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1273 (.I0(n44470), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n42235), .I3(n26495), .O(n2_adj_4631));   // verilog/coms.v(157[9:60])
    defparam i1_3_lut_4_lut_adj_1273.LUT_INIT = 16'h00d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1274 (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n33839), .I3(GND_net), .O(n4_adj_4636));   // verilog/coms.v(263[5:27])
    defparam i1_2_lut_3_lut_adj_1274.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1275 (.I0(n44470), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.state_31__N_2660 [1]), .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2692 [1]));   // verilog/coms.v(157[9:60])
    defparam i1_2_lut_3_lut_adj_1275.LUT_INIT = 16'hf2f2;
    SB_LUT4 add_43_17_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [15]), 
            .I2(GND_net), .I3(n37542), .O(n41477)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1276 (.I0(n62), .I1(n6_adj_4634), .I2(\FRAME_MATCHER.state_31__N_2692 [1]), 
            .I3(n26495), .O(n48857));
    defparam i3_4_lut_adj_1276.LUT_INIT = 16'hddfd;
    SB_CARRY add_43_17 (.CI(n37542), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n37543));
    SB_LUT4 add_43_16_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [14]), 
            .I2(GND_net), .I3(n37541), .O(n41505)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_16 (.CI(n37541), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n37542));
    SB_LUT4 add_43_15_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [13]), 
            .I2(GND_net), .I3(n37540), .O(n41525)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1277 (.I0(n1_adj_4632), .I1(n2_adj_4631), 
            .I2(n1_adj_4637), .I3(\FRAME_MATCHER.state_c [5]), .O(n8_adj_4533));
    defparam i1_2_lut_4_lut_adj_1277.LUT_INIT = 16'hfe00;
    SB_LUT4 n48568_bdd_4_lut (.I0(n48568), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n48571));
    defparam n48568_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1278 (.I0(n1_adj_4632), .I1(n2_adj_4631), 
            .I2(n1_adj_4637), .I3(\FRAME_MATCHER.state_c [22]), .O(n8_adj_4531));
    defparam i1_2_lut_4_lut_adj_1278.LUT_INIT = 16'hfe00;
    SB_CARRY add_43_15 (.CI(n37540), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n37541));
    SB_LUT4 i1_2_lut_4_lut_adj_1279 (.I0(n1_adj_4632), .I1(n2_adj_4631), 
            .I2(n1_adj_4637), .I3(\FRAME_MATCHER.state_c [25]), .O(n8_adj_4527));
    defparam i1_2_lut_4_lut_adj_1279.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1280 (.I0(n1_adj_4632), .I1(n2_adj_4631), 
            .I2(n1_adj_4637), .I3(\FRAME_MATCHER.state_c [26]), .O(n33842));
    defparam i1_2_lut_4_lut_adj_1280.LUT_INIT = 16'hfe00;
    SB_LUT4 add_43_14_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [12]), 
            .I2(GND_net), .I3(n37539), .O(n41547)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n28664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n28663));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_14 (.CI(n37539), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n37540));
    SB_LUT4 add_43_13_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [11]), 
            .I2(GND_net), .I3(n37538), .O(n41567)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1281 (.I0(\data_out_frame[18] [5]), .I1(n42293), 
            .I2(n26531), .I3(n40535), .O(n39584));
    defparam i3_4_lut_adj_1281.LUT_INIT = 16'h9669;
    SB_CARRY add_43_13 (.CI(n37538), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n37539));
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n28662));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n28661));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33137_3_lut_4_lut (.I0(n26268), .I1(n33639), .I2(n33209), 
            .I3(n62), .O(n27701));   // verilog/coms.v(212[5:16])
    defparam i33137_3_lut_4_lut.LUT_INIT = 16'h04ff;
    SB_LUT4 add_43_12_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(n37537), .O(n41587)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_12 (.CI(n37537), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n37538));
    SB_LUT4 i1_3_lut_4_lut_adj_1282 (.I0(n26268), .I1(n33639), .I2(n23516), 
            .I3(n19), .O(n1_adj_4619));   // verilog/coms.v(212[5:16])
    defparam i1_3_lut_4_lut_adj_1282.LUT_INIT = 16'h4000;
    SB_LUT4 add_43_11_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [9]), 
            .I2(GND_net), .I3(n37536), .O(n41615)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_11 (.CI(n37536), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n37537));
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[7] [4]), .I3(\data_out_frame[5] [2]), .O(n42735));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_10_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [8]), 
            .I2(GND_net), .I3(n37535), .O(n41641)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n37535), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n37536));
    SB_LUT4 add_43_9_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n37534), .O(n2_adj_4602)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_9 (.CI(n37534), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n37535));
    SB_LUT4 add_43_8_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n37533), .O(n2_adj_4604)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n28660));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n28659));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n28658));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_8 (.CI(n37533), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n37534));
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n28656));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n28655));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n28654));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n28653));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n28652));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n28651));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n28650));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n28618));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n28617));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n28616));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n28615));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_7_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n37532), .O(n2_adj_4609)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n28612));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_7 (.CI(n37532), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n37533));
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n28604));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n28603));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n28602));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n28601));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n28600));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n28599));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n28598));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n28597));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n28596));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n28595));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n28594));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n28593));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n28592));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n28591));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n28590));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n28589));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n28588));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n28587));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n28586));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n28585));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n28584));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n28583));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n28582));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n28581));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n28580));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n28579));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n28578));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n28577));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n28576));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n28575));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n28574));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n28573));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n28572));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n28571));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n28570));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n28569));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n28568));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n28567));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n28566));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n28565));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n28564));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n28563));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n28562));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n28561));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n28560));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n28559));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n28558));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n28557));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_6_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n37531), .O(n2_adj_4610)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n28556));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n28555));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n28554));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n28553));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n28552));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n28551));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n28550));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n28549));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n28548));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n28547));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_adj_1283 (.I0(\FRAME_MATCHER.state_31__N_2660 [1]), .I1(n20), 
            .I2(n3813), .I3(GND_net), .O(n41655));
    defparam i1_3_lut_adj_1283.LUT_INIT = 16'ha8a8;
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n28546));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n28545));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n28544));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n28543));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_out_frame[21][1] ), .I1(n26860), 
            .I2(GND_net), .I3(GND_net), .O(n42445));
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n28542));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n28541));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n28540));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n28539));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i20138_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(GND_net), .O(n33639));
    defparam i20138_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n28538));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n28537));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n28536));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n28535));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n28534));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n28533));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n28532));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n28531));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n28530));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n28529));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n28528));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n28527));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n28526));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n28525));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n28524));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n28523));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n28522));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n28521));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n28520));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n28519));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45844), .I3(n45842), .O(n7_adj_4608));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n28518));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1285 (.I0(\FRAME_MATCHER.state_c [2]), 
            .I1(\FRAME_MATCHER.state [0]), .I2(n26268), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n26482));
    defparam i2_2_lut_3_lut_4_lut_adj_1285.LUT_INIT = 16'hfff7;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n28517));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1286 (.I0(\data_out_frame[23] [1]), .I1(\data_out_frame[21][1] ), 
            .I2(n26860), .I3(\data_out_frame[18] [4]), .O(n42772));
    defparam i2_3_lut_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n28516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n28515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n28514));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n28510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n28509));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n28508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n28507));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n28506));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n28505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n28501));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n28500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n28499));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n28498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n28497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n28496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n28495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n28494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n28493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n28492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n28491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n28490));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n28489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n28488));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n28487));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n28483));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n45820), .I3(n45818), .O(n7_adj_4514));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_CARRY add_43_6 (.CI(n37531), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n37532));
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n28482));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1287 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [1]), .I3(GND_net), .O(n42599));
    defparam i1_2_lut_3_lut_adj_1287.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1288 (.I0(n40510), .I1(n44349), .I2(\data_out_frame[25] [3]), 
            .I3(\data_out_frame[25] [2]), .O(n44255));
    defparam i2_3_lut_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1289 (.I0(\data_out_frame[25] [5]), .I1(n42445), 
            .I2(n27252), .I3(\data_out_frame[23] [4]), .O(n10_adj_4639));
    defparam i4_4_lut_adj_1289.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_5_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n37530), .O(n2_adj_4612)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[13] [0]), .I3(GND_net), .O(n6_adj_4640));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1291 (.I0(\FRAME_MATCHER.state_c [2]), .I1(n88), 
            .I2(\FRAME_MATCHER.state_31__N_2724 [3]), .I3(n26496), .O(n10_adj_4534));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1291.LUT_INIT = 16'hccdc;
    SB_LUT4 i5_3_lut_adj_1292 (.I0(\data_out_frame[23] [3]), .I1(n10_adj_4639), 
            .I2(n39556), .I3(GND_net), .O(n42687));
    defparam i5_3_lut_adj_1292.LUT_INIT = 16'h9696;
    SB_CARRY add_43_5 (.CI(n37530), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n37531));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1293 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[5] [2]), .O(n42487));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i15139_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n28653));
    defparam i15139_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15140_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n28654));
    defparam i15140_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1294 (.I0(\FRAME_MATCHER.state_c [4]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41657));
    defparam i1_2_lut_adj_1294.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1295 (.I0(\data_out_frame[18] [2]), .I1(n39625), 
            .I2(\data_out_frame[22] [5]), .I3(n40258), .O(n43547));
    defparam i2_3_lut_4_lut_adj_1295.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1296 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[20] [2]), 
            .I2(\data_out_frame[24] [6]), .I3(n42537), .O(n42652));
    defparam i2_3_lut_4_lut_adj_1296.LUT_INIT = 16'h9669;
    SB_LUT4 i15141_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n28655));
    defparam i15141_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15142_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n28656));
    defparam i15142_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1297 (.I0(n27084), .I1(n26912), .I2(\data_out_frame[17] [7]), 
            .I3(\data_out_frame[15] [6]), .O(n42627));
    defparam i1_2_lut_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1298 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41721));
    defparam i1_2_lut_adj_1298.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1299 (.I0(n26912), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n27378));
    defparam i1_2_lut_3_lut_adj_1299.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1300 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[15] [4]), 
            .I2(n39506), .I3(n27374), .O(n6_adj_4642));
    defparam i2_2_lut_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_4_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n37529), .O(n2_adj_4613)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n28479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n28478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n28477));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n28476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n28475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n28474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n28473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n28472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n28471));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state_c [2]), .C(CLK_c), 
           .D(n48873));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n28469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n28468));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n28467));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n28466));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n28465));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n28464));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1301 (.I0(n39586), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42754));
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n28463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n28462));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n28457));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n28456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n28455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n28454));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n28453));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n28452));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n28451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n28450));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n28449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n28448));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n28447));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i880_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1668));   // verilog/coms.v(85[17:28])
    defparam i880_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n28446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n28445));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n28444));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n28443));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n28442));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n28441));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n28440));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_4 (.CI(n37529), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n37530));
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n28439));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n28438));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n28433));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15144_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n28658));
    defparam i15144_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n28432));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n28428));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1302 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[6] [5]), 
            .I2(\data_in_frame[6] [4]), .I3(n42766), .O(n42941));
    defparam i1_2_lut_3_lut_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n28426));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15145_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n28659));
    defparam i15145_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n28425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n28424));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n28423));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n28422));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n28421));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n28420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n28419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n28418));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n28417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n28416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n28415));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n28414));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n28413));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n28412));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n28411));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n28410));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n28409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n28408));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15146_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n28660));
    defparam i15146_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n28407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n28406));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n28405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n28404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n28403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n28402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n28401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n28400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n28399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n28398));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1303 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n42518));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1303.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n28397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n28396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n28395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n28394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n28393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n28392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n28391));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30860_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n45990), .I3(n20_adj_4505), .O(n45991));
    defparam i30860_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n28390));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1304 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26553));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1304.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n28389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n28384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n28383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n28382));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_3_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n37528), .O(n2_adj_4614)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n28381));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n28380));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n28379));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15147_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42260), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n28661));
    defparam i15147_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n28378));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n28377));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n28376));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n28375));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n28374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n28373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n28372));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_3 (.CI(n37528), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n37529));
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n28371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n28370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n28369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n28368));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1305 (.I0(n42518), .I1(n42808), .I2(\data_out_frame[10] [6]), 
            .I3(GND_net), .O(n42316));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1305.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n28367));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n28366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n28365));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1306 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41719));
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h8888;
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n28364));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n28363));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n28362));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n28361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n28360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n28359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n28358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n28357));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n28356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n28355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n28354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n28353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n28352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n28351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n28350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n28349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n28348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n28347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n28346));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_2_lut (.I0(n6_adj_4633), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n28345));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n28344));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n28343));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n37528));
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n28342));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n28341));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n28340));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n28335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n28331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n28329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n28328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n28327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n28326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n28325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n28324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n28323));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n28322));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n28321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n28320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n28319));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(CLK_c), 
           .D(n28317));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n28316));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1307 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[22] [3]), .I3(GND_net), .O(n42956));
    defparam i1_2_lut_3_lut_adj_1307.LUT_INIT = 16'h9696;
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n28314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(CLK_c), 
           .D(n28313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(CLK_c), 
           .D(n28312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n28311));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1308 (.I0(n42316), .I1(\data_out_frame[4] [2]), 
            .I2(n42702), .I3(n6_adj_4640), .O(n39574));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n28310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n28309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n28308));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n28156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n28307));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n28306));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n28305));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(CLK_c), 
           .D(n28304));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1309 (.I0(n39574), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42853));
    defparam i1_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\data_out_frame[21][4] ), .I1(\data_out_frame[23] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n42417));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h6666;
    SB_LUT4 i30854_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n45984), .I3(n20_adj_4509), .O(n45985));
    defparam i30854_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_3_lut_adj_1311 (.I0(\data_out_frame[18] [6]), .I1(n43849), 
            .I2(n39584), .I3(GND_net), .O(n27252));
    defparam i1_2_lut_3_lut_adj_1311.LUT_INIT = 16'h6969;
    SB_LUT4 i3_3_lut_4_lut (.I0(\data_in[0] [6]), .I1(\data_in[0] [3]), 
            .I2(\data_in[1] [0]), .I3(\data_in[3] [0]), .O(n99));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_adj_1312 (.I0(\FRAME_MATCHER.state_c [8]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41717));
    defparam i1_2_lut_adj_1312.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_3_lut_adj_1313 (.I0(\data_out_frame[18] [6]), .I1(n43849), 
            .I2(\data_out_frame[21][0] ), .I3(GND_net), .O(n10_adj_4643));
    defparam i2_2_lut_3_lut_adj_1313.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1314 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [4]), 
            .I2(n42968), .I3(\data_out_frame[16] [6]), .O(n42696));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1315 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[20] [7]), .I3(n40513), .O(n43849));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1315.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1316 (.I0(\data_out_frame[20] [3]), .I1(n42536), 
            .I2(\data_out_frame[24] [5]), .I3(n42823), .O(n42947));
    defparam i2_3_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1317 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41715));
    defparam i1_2_lut_adj_1317.LUT_INIT = 16'h8888;
    SB_LUT4 i30851_3_lut_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[1]), 
            .I2(n45981), .I3(n20_adj_4512), .O(n45982));
    defparam i30851_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1318 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(n27125), .O(n42407));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1318.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1319 (.I0(\FRAME_MATCHER.state_c [1]), .I1(n26268), 
            .I2(n60), .I3(n33835), .O(n3846));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1319.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41713));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1321 (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n26268), .I3(\FRAME_MATCHER.state_c [1]), .O(n26495));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_4_lut_adj_1321.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_2_lut_4_lut_adj_1322 (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n26268), .I3(n26482), .O(n33835));   // verilog/coms.v(254[5:25])
    defparam i2_2_lut_4_lut_adj_1322.LUT_INIT = 16'hfb00;
    SB_LUT4 i1_2_lut_4_lut_adj_1323 (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n26268), .I3(\FRAME_MATCHER.state_c [1]), .O(n26494));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_4_lut_adj_1323.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut_adj_1324 (.I0(n42458), .I1(n42775), .I2(\data_out_frame[17] [0]), 
            .I3(\data_out_frame[16] [6]), .O(n42944));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1324.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1325 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41663));
    defparam i1_2_lut_adj_1325.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1326 (.I0(n42458), .I1(n42775), .I2(n42689), 
            .I3(GND_net), .O(n40513));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1326.LUT_INIT = 16'h9696;
    SB_LUT4 i32809_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(n33300), 
            .I2(n26421), .I3(n33839), .O(n43482));
    defparam i32809_3_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i1_2_lut_adj_1327 (.I0(\FRAME_MATCHER.state_c [12]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41711));
    defparam i1_2_lut_adj_1327.LUT_INIT = 16'h8888;
    SB_LUT4 i15156_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n28670));
    defparam i15156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(\FRAME_MATCHER.state_c [13]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41709));
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1329 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41707));
    defparam i1_2_lut_adj_1329.LUT_INIT = 16'h8888;
    SB_LUT4 i28170_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(n33300), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n33839), .O(n43197));
    defparam i28170_3_lut_4_lut.LUT_INIT = 16'hffe0;
    SB_LUT4 i1_2_lut_adj_1330 (.I0(\FRAME_MATCHER.state [3]), .I1(n33839), 
            .I2(GND_net), .I3(GND_net), .O(n26268));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_adj_1330.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1331 (.I0(n33839), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i2_2_lut_adj_1331.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n60));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'heeee;
    SB_LUT4 i19714_2_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3616[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n33209));
    defparam i19714_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut_adj_1333 (.I0(n60), .I1(n6), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n62));
    defparam i3_3_lut_adj_1333.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1334 (.I0(n39586), .I1(\data_out_frame[23] [4]), 
            .I2(n42687), .I3(GND_net), .O(n6_adj_4646));
    defparam i1_2_lut_3_lut_adj_1334.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(\FRAME_MATCHER.state_c [15]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41705));
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1336 (.I0(n27196), .I1(n27203), .I2(n39554), 
            .I3(n26809), .O(n40521));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_4_lut_adj_1336.LUT_INIT = 16'h6996;
    SB_LUT4 i15157_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n28671));
    defparam i15157_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15158_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n28672));
    defparam i15158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15159_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n28673));
    defparam i15159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1337 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[17] [2]), 
            .I2(n42853), .I3(n6_adj_4647), .O(n40529));
    defparam i4_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41667));
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h8888;
    SB_LUT4 i15161_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n28675));
    defparam i15161_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1339 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[16] [7]), .I3(n42944), .O(n6_adj_4647));
    defparam i1_2_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1340 (.I0(\FRAME_MATCHER.state_c [17]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41703));
    defparam i1_2_lut_adj_1340.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1341 (.I0(\FRAME_MATCHER.state_c [2]), 
            .I1(\FRAME_MATCHER.state_c [1]), .I2(\FRAME_MATCHER.state [0]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n42163));
    defparam i1_2_lut_3_lut_4_lut_adj_1341.LUT_INIT = 16'h0100;
    SB_LUT4 i15162_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n28676));
    defparam i15162_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(\FRAME_MATCHER.state_c [18]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41701));
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h8888;
    SB_LUT4 i15163_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n28677));
    defparam i15163_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\FRAME_MATCHER.state_c [19]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41699));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1344 (.I0(\FRAME_MATCHER.state_c [1]), .I1(n33839), 
            .I2(n42163), .I3(GND_net), .O(n27647));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_adj_1344.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_adj_1345 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41697));
    defparam i1_2_lut_adj_1345.LUT_INIT = 16'h8888;
    SB_LUT4 i15164_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42260), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n28678));
    defparam i15164_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1346 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n7233));
    defparam i1_2_lut_3_lut_adj_1346.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_adj_1347 (.I0(\FRAME_MATCHER.state_c [21]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41695));
    defparam i1_2_lut_adj_1347.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1348 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[10] [4]), .I3(\data_out_frame[6] [0]), .O(n42702));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1348.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1349 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[12] [7]), 
            .I2(\data_out_frame[12] [6]), .I3(GND_net), .O(n42808));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1349.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1350 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4529));
    defparam i1_2_lut_adj_1350.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1351 (.I0(\FRAME_MATCHER.state [3]), .I1(n3813), 
            .I2(n23516), .I3(n3_adj_4620), .O(n41661));
    defparam i1_3_lut_4_lut_adj_1351.LUT_INIT = 16'haa80;
    SB_LUT4 i1_2_lut_adj_1352 (.I0(\FRAME_MATCHER.state_c [24]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41693));
    defparam i1_2_lut_adj_1352.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_4_lut_adj_1353 (.I0(\FRAME_MATCHER.state [3]), .I1(n33839), 
            .I2(\FRAME_MATCHER.state [0]), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n26496));   // verilog/coms.v(231[5:23])
    defparam i2_2_lut_4_lut_adj_1353.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_4_lut_adj_1354 (.I0(n42471), .I1(n42561), .I2(Kp_23__N_1195), 
            .I3(n26617), .O(n42708));
    defparam i1_2_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_4_lut (.I0(n42471), .I1(n42561), .I2(Kp_23__N_1195), 
            .I3(n40499), .O(n15_adj_4453));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\FRAME_MATCHER.state_c [27]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4524));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1356 (.I0(n3813), .I1(n26495), .I2(n44470), .I3(\FRAME_MATCHER.i [31]), 
            .O(n4_adj_4648));
    defparam i1_4_lut_adj_1356.LUT_INIT = 16'hbbab;
    SB_LUT4 i2_4_lut_adj_1357 (.I0(\FRAME_MATCHER.state_c [28]), .I1(n23516), 
            .I2(n43068), .I3(n4_adj_4648), .O(n43514));   // verilog/coms.v(95[12:19])
    defparam i2_4_lut_adj_1357.LUT_INIT = 16'h8808;
    SB_LUT4 i1_2_lut_4_lut_adj_1358 (.I0(n42471), .I1(n42561), .I2(Kp_23__N_1195), 
            .I3(\data_in_frame[11] [3]), .O(n42370));
    defparam i1_2_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_4_lut_4_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state_31__N_2724 [3]), .I3(\FRAME_MATCHER.state_c [1]), 
            .O(n6_adj_4599));
    defparam i2_4_lut_4_lut_4_lut.LUT_INIT = 16'h8988;
    SB_LUT4 i1_3_lut_4_lut_adj_1359 (.I0(\data_in_frame[18] [7]), .I1(n40264), 
            .I2(\data_in_frame[16] [5]), .I3(n39631), .O(n15_adj_4465));
    defparam i1_3_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i14640_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n33839), 
            .I2(n33639), .I3(n27701), .O(n28149));   // verilog/coms.v(212[5:16])
    defparam i14640_2_lut_3_lut_4_lut.LUT_INIT = 16'hef00;
    SB_LUT4 i1_2_lut_adj_1360 (.I0(\FRAME_MATCHER.state_c [29]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41689));
    defparam i1_2_lut_adj_1360.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1361 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n33839), .I2(n33639), .I3(n19), .O(n20));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1361.LUT_INIT = 16'h1000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1362 (.I0(n99), .I1(n121), .I2(n42251), 
            .I3(n122), .O(\FRAME_MATCHER.state_31__N_2660[2] ));   // verilog/coms.v(95[12:19])
    defparam i1_2_lut_3_lut_4_lut_adj_1362.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1363 (.I0(n2_adj_4631), .I1(n1_adj_4632), 
            .I2(n3813), .I3(n23516), .O(n6_adj_4641));
    defparam i1_2_lut_3_lut_4_lut_adj_1363.LUT_INIT = 16'hfeee;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(\data_in_frame[18] [7]), .I1(n40264), 
            .I2(n39631), .I3(n40531), .O(n8_adj_4489));
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1365 (.I0(\data_in_frame[18] [7]), .I1(n40264), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[19] [1]), .O(n8_adj_4499));
    defparam i3_3_lut_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(n27196), .I1(n27203), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n27095));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n33839), .O(n33873));
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'hfffe;
    SB_LUT4 i19742_2_lut_3_lut (.I0(n33835), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n33239));
    defparam i19742_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_4_lut_adj_1368 (.I0(n39554), .I1(n27203), .I2(\data_in_frame[9] [4]), 
            .I3(\data_in_frame[11] [5]), .O(n42637));
    defparam i1_2_lut_4_lut_adj_1368.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1369 (.I0(n39554), .I1(n27203), .I2(\data_in_frame[9] [4]), 
            .I3(\data_in_frame[9] [5]), .O(n40499));
    defparam i1_2_lut_4_lut_adj_1369.LUT_INIT = 16'h6996;
    SB_LUT4 i15049_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n28563));
    defparam i15049_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15050_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n28564));
    defparam i15050_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15051_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n28565));
    defparam i15051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15052_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n28566));
    defparam i15052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15053_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n28567));
    defparam i15053_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1370 (.I0(n40529), .I1(n42417), .I2(\data_out_frame[25] [6]), 
            .I3(n6_adj_4646), .O(n44528));
    defparam i4_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1371 (.I0(n39569), .I1(n42579), .I2(\data_out_frame[19] [4]), 
            .I3(\data_out_frame[21][4] ), .O(n42850));
    defparam i1_2_lut_4_lut_adj_1371.LUT_INIT = 16'h9669;
    SB_LUT4 i15054_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n28568));
    defparam i15054_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1372 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41687));
    defparam i1_2_lut_adj_1372.LUT_INIT = 16'h8888;
    SB_LUT4 i15055_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n28569));
    defparam i15055_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15056_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42274), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n28570));
    defparam i15056_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i32750_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n27964));
    defparam i32750_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_4_lut_4_lut_adj_1373 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(n1), .I3(\FRAME_MATCHER.state_c [1]), .O(n5_adj_4598));
    defparam i1_4_lut_4_lut_adj_1373.LUT_INIT = 16'h6273;
    SB_LUT4 i14702_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n28216));
    defparam i14702_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15249_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n28763));
    defparam i15249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15250_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n28764));
    defparam i15250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1374 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4649));
    defparam i2_2_lut_adj_1374.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1375 (.I0(\FRAME_MATCHER.i [0]), .I1(n6_adj_4649), 
            .I2(n26289), .I3(\FRAME_MATCHER.i [1]), .O(n44470));
    defparam i3_4_lut_adj_1375.LUT_INIT = 16'hfefc;
    SB_LUT4 i1_2_lut_adj_1376 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4650));   // verilog/coms.v(231[5:23])
    defparam i1_2_lut_adj_1376.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_1377 (.I0(n33835), .I1(n4_adj_4636), .I2(n62), 
            .I3(n33300), .O(n8_adj_4651));
    defparam i3_4_lut_adj_1377.LUT_INIT = 16'ha080;
    SB_LUT4 i4_4_lut_adj_1378 (.I0(n26268), .I1(n8_adj_4651), .I2(n4_adj_4650), 
            .I3(n33639), .O(n3813));
    defparam i4_4_lut_adj_1378.LUT_INIT = 16'h88c8;
    SB_LUT4 i1_2_lut_4_lut_adj_1379 (.I0(n39569), .I1(n42579), .I2(\data_out_frame[19] [4]), 
            .I3(\data_out_frame[23] [7]), .O(n40487));
    defparam i1_2_lut_4_lut_adj_1379.LUT_INIT = 16'h9669;
    SB_LUT4 i15251_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n28765));
    defparam i15251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15252_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n28766));
    defparam i15252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15253_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n28767));
    defparam i15253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1380 (.I0(\FRAME_MATCHER.i [4]), .I1(n26414), .I2(GND_net), 
            .I3(GND_net), .O(n26289));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1380.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1381 (.I0(n26989), .I1(\data_out_frame[15] [0]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n42785));
    defparam i1_2_lut_3_lut_adj_1381.LUT_INIT = 16'h9696;
    SB_LUT4 i15254_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n28768));
    defparam i15254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15255_3_lut_4_lut (.I0(n8_adj_4592), .I1(n42281), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n28769));
    defparam i15255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i12_2_lut_4_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[5] [5]), .I3(n26511), .O(n37_adj_4582));   // verilog/coms.v(73[16:42])
    defparam i12_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1382 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n42254), .I3(\FRAME_MATCHER.i [3]), .O(n42255));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1382.LUT_INIT = 16'hfeff;
    SB_LUT4 equal_304_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4515));   // verilog/coms.v(154[7:23])
    defparam equal_304_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 n48838_bdd_4_lut (.I0(n48838), .I1(\data_out_frame[21][4] ), 
            .I2(\data_out_frame[20] [4]), .I3(byte_transmit_counter[1]), 
            .O(n48841));
    defparam n48838_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i28037_4_lut (.I0(n8_adj_4592), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n26289), .I3(\FRAME_MATCHER.i [3]), .O(n3303));
    defparam i28037_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_3_lut_adj_1383 (.I0(n3303), .I1(n26482), .I2(n42235), .I3(GND_net), 
            .O(n1_adj_4632));
    defparam i1_3_lut_adj_1383.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_4_lut_adj_1384 (.I0(n1168), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[5] [0]), .I3(\data_out_frame[4] [6]), .O(n27257));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1385 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n33239), .I3(\FRAME_MATCHER.i [3]), .O(n42260));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1385.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n26511));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1387 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[4] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[6] [5]), .O(n42814));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1388 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n42325), .I3(n27125), .O(n27401));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1389 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[4] [2]), 
            .I2(n26643), .I3(GND_net), .O(n22_adj_4547));   // verilog/coms.v(78[16:27])
    defparam i2_2_lut_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 i15041_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n28555));
    defparam i15041_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1390 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[1] [1]), .O(n42658));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1391 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n42711));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1391.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1392 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[3] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[3] [5]), .O(n42328));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1393 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [4]), .I3(n42962), .O(Kp_23__N_988));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1394 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[1] [3]), .O(n42962));   // verilog/coms.v(96[12:25])
    defparam i2_3_lut_4_lut_adj_1394.LUT_INIT = 16'h6996;
    SB_LUT4 i15042_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n28556));
    defparam i15042_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(n3813), .I1(n23516), .I2(GND_net), 
            .I3(GND_net), .O(n1_adj_4637));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h8888;
    SB_LUT4 i32806_2_lut (.I0(n34010), .I1(n19799), .I2(GND_net), .I3(GND_net), 
            .O(tx_transmit_N_3513));
    defparam i32806_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_3_lut_adj_1396 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n26661));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1396.LUT_INIT = 16'h9696;
    SB_LUT4 i15043_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n28557));
    defparam i15043_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18_4_lut_adj_1397 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut_adj_1397.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n6_adj_4542));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'h9696;
    SB_LUT4 i15044_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n28558));
    defparam i15044_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1399 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_4652));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut_adj_1399.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1400 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_4653));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut_adj_1400.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1401 (.I0(\data_in_frame[3] [7]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[4] [0]), .O(n42705));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1402 (.I0(n40583), .I1(n42299), .I2(GND_net), 
            .I3(GND_net), .O(n27276));
    defparam i1_2_lut_adj_1402.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1403 (.I0(n39556), .I1(n40529), .I2(\data_out_frame[25] [7]), 
            .I3(n42850), .O(n6_adj_4422));
    defparam i1_2_lut_4_lut_adj_1403.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1404 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n26855));
    defparam i1_2_lut_3_lut_adj_1404.LUT_INIT = 16'h9696;
    SB_LUT4 i15045_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n28559));
    defparam i15045_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15046_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n28560));
    defparam i15046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15047_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n28561));
    defparam i15047_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1405 (.I0(n39556), .I1(n40529), .I2(\data_out_frame[25] [7]), 
            .I3(n40487), .O(n6_adj_4424));
    defparam i1_2_lut_4_lut_adj_1405.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1406 (.I0(\data_out_frame[19] [7]), .I1(n42652), 
            .I2(n42947), .I3(n43547), .O(n12_adj_4654));
    defparam i5_4_lut_adj_1406.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1407 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_4655));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut_adj_1407.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1408 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_4656));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut_adj_1408.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1409 (.I0(n42426), .I1(n12_adj_4654), .I2(n42874), 
            .I3(n27276), .O(n43608));
    defparam i6_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1410 (.I0(\data_in_frame[6] [5]), .I1(\data_in_frame[6] [4]), 
            .I2(Kp_23__N_1096), .I3(Kp_23__N_1099), .O(Kp_23__N_1195));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i15048_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42274), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n28562));
    defparam i15048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15033_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n28547));
    defparam i15033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15034_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n28548));
    defparam i15034_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4657));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15035_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n28549));
    defparam i15035_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24_4_lut_adj_1411 (.I0(n41_adj_4655), .I1(n43_adj_4653), .I2(n42_adj_4652), 
            .I3(n44), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut_adj_1411.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1412 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut_adj_1412.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39_adj_4657), .I3(n40_adj_4656), 
            .O(n26414));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(n27133), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n6_adj_4539));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1414 (.I0(n26477), .I1(\data_in[3] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4658));
    defparam i1_2_lut_adj_1414.LUT_INIT = 16'heeee;
    SB_LUT4 i15036_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n28550));
    defparam i15036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1415 (.I0(\data_in[1] [2]), .I1(\data_in[3] [2]), 
            .I2(\data_in[2] [5]), .I3(n10_adj_4658), .O(n16_adj_4659));
    defparam i7_4_lut_adj_1415.LUT_INIT = 16'hff7f;
    SB_LUT4 i2_4_lut_adj_1416 (.I0(\data_in[2] [6]), .I1(\data_in[0] [5]), 
            .I2(\data_in[0] [1]), .I3(\data_in[2] [0]), .O(n11_adj_4660));
    defparam i2_4_lut_adj_1416.LUT_INIT = 16'hbfff;
    SB_LUT4 i1_2_lut_4_lut_adj_1417 (.I0(n26713), .I1(n42345), .I2(\data_in_frame[3] [0]), 
            .I3(n42340), .O(n27289));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n42319));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1419 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[10] [3]), .I3(\data_out_frame[10] [4]), 
            .O(n8_adj_4544));   // verilog/coms.v(85[17:63])
    defparam i3_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i15037_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n28551));
    defparam i15037_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1420 (.I0(n11_adj_4660), .I1(n16_adj_4659), .I2(\data_in[1] [6]), 
            .I3(\data_in[1] [3]), .O(n42251));
    defparam i8_4_lut_adj_1420.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1421 (.I0(n121), .I1(n42251), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4625));
    defparam i1_2_lut_adj_1421.LUT_INIT = 16'heeee;
    SB_LUT4 i2_2_lut_adj_1422 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4661));
    defparam i2_2_lut_adj_1422.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_4_lut_adj_1423 (.I0(\data_in_frame[6] [1]), .I1(n42319), 
            .I2(n42705), .I3(\data_in_frame[1] [6]), .O(n42748));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1424 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4662));
    defparam i6_4_lut_adj_1424.LUT_INIT = 16'hfeff;
    SB_LUT4 i5_3_lut_4_lut_adj_1425 (.I0(\data_in_frame[5] [1]), .I1(n42744), 
            .I2(n10_adj_4520), .I3(n26661), .O(n27203));
    defparam i5_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1426 (.I0(\data_in[3] [6]), .I1(n14_adj_4662), 
            .I2(n10_adj_4661), .I3(\data_in[2] [1]), .O(n26477));
    defparam i7_4_lut_adj_1426.LUT_INIT = 16'hfffd;
    SB_LUT4 i3_3_lut_4_lut_adj_1427 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[5] [5]), 
            .I2(\data_in_frame[1] [3]), .I3(n42389), .O(n8_adj_4518));
    defparam i3_3_lut_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i30642_2_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n45674));
    defparam i30642_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15038_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n28552));
    defparam i15038_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15039_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n28553));
    defparam i15039_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15040_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42274), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n28554));
    defparam i15040_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15241_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n28755));
    defparam i15241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1428 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4627));
    defparam i4_4_lut_adj_1428.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_3_lut_4_lut_adj_1429 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[11] [6]), 
            .O(n42726));
    defparam i2_3_lut_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1430 (.I0(\data_out_frame[6] [1]), .I1(n10_adj_4501), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[10] [2]), .O(n1516));   // verilog/coms.v(85[17:70])
    defparam i5_3_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1431 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [2]), 
            .I2(\data_out_frame[11] [1]), .I3(GND_net), .O(n42439));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1431.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1432 (.I0(n7_adj_4629), .I1(\data_in[2] [2]), .I2(\data_in[1] [4]), 
            .I3(\data_in[1] [5]), .O(n121));
    defparam i4_4_lut_adj_1432.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_1433 (.I0(\data_out_frame[19] [3]), .I1(n43671), 
            .I2(GND_net), .I3(GND_net), .O(n42579));
    defparam i1_2_lut_adj_1433.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1434 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[22] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n42874));
    defparam i1_2_lut_adj_1434.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1435 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4663));
    defparam i6_4_lut_adj_1435.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_4_lut_adj_1436 (.I0(\data_in_frame[20] [2]), .I1(n42500), 
            .I2(n10_adj_4485), .I3(\data_in_frame[18] [0]), .O(n4_adj_4494));
    defparam i1_2_lut_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1437 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4664));
    defparam i7_4_lut_adj_1437.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1438 (.I0(n17_adj_4664), .I1(\data_in[1] [6]), 
            .I2(n16_adj_4663), .I3(\data_in[3] [7]), .O(n26403));
    defparam i9_4_lut_adj_1438.LUT_INIT = 16'hfbff;
    SB_LUT4 i15242_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n28756));
    defparam i15242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1439 (.I0(n99), .I1(n121), .I2(GND_net), .I3(GND_net), 
            .O(n32652));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1439.LUT_INIT = 16'heeee;
    SB_LUT4 i15243_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n28757));
    defparam i15243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1440 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n32652), .O(n16_adj_4665));
    defparam i6_4_lut_adj_1440.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_1441 (.I0(\data_in_frame[9] [2]), .I1(n26756), 
            .I2(n27196), .I3(GND_net), .O(n42720));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1442 (.I0(n26403), .I1(\data_in[3] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[2] [3]), .O(n17_adj_4666));
    defparam i7_4_lut_adj_1442.LUT_INIT = 16'hbfff;
    SB_LUT4 i2_3_lut_adj_1443 (.I0(\data_out_frame[22] [0]), .I1(\data_out_frame[23] [6]), 
            .I2(\data_out_frame[24] [0]), .I3(GND_net), .O(n42613));
    defparam i2_3_lut_adj_1443.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1444 (.I0(n42348), .I1(\data_out_frame[17] [4]), 
            .I2(n27374), .I3(GND_net), .O(n42400));
    defparam i2_3_lut_adj_1444.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1445 (.I0(n17_adj_4666), .I1(\data_in[3] [5]), 
            .I2(n16_adj_4665), .I3(\data_in[3] [1]), .O(n63_adj_4586));
    defparam i9_4_lut_adj_1445.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_4_lut_adj_1446 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[5] [6]), 
            .I2(\data_in_frame[9] [7]), .I3(n27451), .O(n14_adj_4480));   // verilog/coms.v(78[16:27])
    defparam i5_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1447 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n42841));
    defparam i1_2_lut_3_lut_adj_1447.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1448 (.I0(n40472), .I1(n42630), .I2(n10_adj_4473), 
            .I3(\data_in_frame[15] [3]), .O(n42859));
    defparam i5_3_lut_4_lut_adj_1448.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1449 (.I0(n42449), .I1(n42766), .I2(\data_in_frame[8] [4]), 
            .I3(GND_net), .O(n26687));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1449.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(\data_in_frame[10] [3]), .I1(n26784), 
            .I2(n42433), .I3(GND_net), .O(n26938));
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1451 (.I0(n26789), .I1(n27215), .I2(\data_in_frame[12] [7]), 
            .I3(\data_in_frame[10] [6]), .O(n27227));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1452 (.I0(n42637), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[13] [6]), .I3(\data_in_frame[15] [7]), .O(n42555));
    defparam i2_3_lut_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i15244_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n28758));
    defparam i15244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15245_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n28759));
    defparam i15245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1453 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n26801), .I3(n26809), .O(n39321));
    defparam i2_3_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1454 (.I0(n26477), .I1(\data_in[1] [0]), .I2(\data_in[0] [6]), 
            .I3(\data_in[1] [4]), .O(n18_adj_4667));
    defparam i7_4_lut_adj_1454.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1455 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[11] [4]), .I3(GND_net), .O(n27071));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1455.LUT_INIT = 16'h9696;
    SB_LUT4 i15246_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n28760));
    defparam i15246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1456 (.I0(n1516), .I1(\data_out_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4668));
    defparam i2_2_lut_adj_1456.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1457 (.I0(\data_out_frame[19] [5]), .I1(n42893), 
            .I2(n42853), .I3(n42331), .O(n14_adj_4669));
    defparam i6_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1458 (.I0(\data_out_frame[19] [4]), .I1(n14_adj_4669), 
            .I2(n10_adj_4668), .I3(n42400), .O(n2134));
    defparam i7_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1459 (.I0(\data_out_frame[20] [0]), .I1(n42400), 
            .I2(n6_adj_4642), .I3(\data_out_frame[17] [6]), .O(n42675));
    defparam i1_4_lut_adj_1459.LUT_INIT = 16'h9669;
    SB_LUT4 i15247_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n28761));
    defparam i15247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15248_3_lut_4_lut (.I0(n8_adj_4621), .I1(n42281), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n28762));
    defparam i15248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1460 (.I0(n26403), .I1(\data_in[0] [3]), .I2(\data_in[3] [0]), 
            .I3(\data_in[2] [2]), .O(n19_adj_4670));
    defparam i8_4_lut_adj_1460.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1461 (.I0(n19_adj_4670), .I1(\data_in[2] [4]), 
            .I2(n18_adj_4667), .I3(n12_adj_4628), .O(n63));
    defparam i10_4_lut_adj_1461.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_4_lut_adj_1462 (.I0(n27329), .I1(n10_adj_4410), .I2(\data_out_frame[11] [4]), 
            .I3(n42293), .O(n42856));
    defparam i1_2_lut_4_lut_adj_1462.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1463 (.I0(\data_out_frame[10] [0]), .I1(n10_adj_4611), 
            .I2(\data_out_frame[10] [1]), .I3(n42616), .O(n40535));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1464 (.I0(n26756), .I1(Kp_23__N_1214), .I2(\data_in_frame[8] [7]), 
            .I3(\data_in_frame[9] [1]), .O(n26617));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1465 (.I0(n45674), .I1(\data_in[0] [6]), .I2(\data_in[3] [0]), 
            .I3(n7_adj_4625), .O(n126));
    defparam i4_4_lut_adj_1465.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1466 (.I0(\data_out_frame[7] [3]), .I1(n24129), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[9] [5]), .O(n42760));
    defparam i1_2_lut_3_lut_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1467 (.I0(\data_out_frame[15] [1]), .I1(n1519), 
            .I2(GND_net), .I3(GND_net), .O(n42331));
    defparam i1_2_lut_adj_1467.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1468 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4671));
    defparam i1_2_lut_adj_1468.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1469 (.I0(n42484), .I1(n42331), .I2(n42788), 
            .I3(n6_adj_4671), .O(n39569));
    defparam i4_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1470 (.I0(\data_out_frame[10] [0]), .I1(n10_adj_4611), 
            .I2(\data_out_frame[10] [1]), .I3(\data_out_frame[14] [4]), 
            .O(n42775));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1471 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[8] [1]), 
            .I2(n39558), .I3(GND_net), .O(n6_adj_4444));
    defparam i1_2_lut_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1472 (.I0(\data_out_frame[19] [5]), .I1(n39569), 
            .I2(GND_net), .I3(GND_net), .O(n42799));
    defparam i1_2_lut_adj_1472.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1473 (.I0(n42484), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[15] [3]), .I3(\data_out_frame[17] [5]), 
            .O(n42506));
    defparam i4_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_3_lut (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[7] [3]), 
            .I2(n42430), .I3(GND_net), .O(n26));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1474 (.I0(n42675), .I1(n2134), .I2(\data_out_frame[24] [2]), 
            .I3(n27282), .O(n42884));
    defparam i3_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1475 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [7]), 
            .I2(\data_in_frame[14] [5]), .I3(GND_net), .O(n42302));
    defparam i1_2_lut_3_lut_adj_1475.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1476 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[24] [1]), 
            .I2(n4_adj_4624), .I3(\data_out_frame[22] [1]), .O(n42521));
    defparam i2_4_lut_adj_1476.LUT_INIT = 16'h9669;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[22] [2]), .I1(\data_out_frame[23] [7]), 
            .I2(n42772), .I3(n42521), .O(n64));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[20] [7]), .I3(\data_out_frame[17] [3]), 
            .O(n68));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1477 (.I0(n42929), .I1(n40525), .I2(n42655), 
            .I3(\data_out_frame[24] [5]), .O(n66));
    defparam i24_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1478 (.I0(n27329), .I1(n10_adj_4410), .I2(\data_out_frame[11] [4]), 
            .I3(n39567), .O(n40525));
    defparam i1_2_lut_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i15017_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n28531));
    defparam i15017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1479 (.I0(\data_in_frame[10] [7]), .I1(n10_adj_4442), 
            .I2(n26667), .I3(n42334), .O(n44139));
    defparam i5_3_lut_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1480 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[23] [2]), .I3(\data_out_frame[17] [6]), 
            .O(n67));
    defparam i25_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_4_lut (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[9] [7]), 
            .I2(n42630), .I3(GND_net), .O(n13));
    defparam i5_4_lut_4_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i23_4_lut_adj_1481 (.I0(n42971), .I1(\data_out_frame[14] [4]), 
            .I2(n42613), .I3(n39510), .O(n65));
    defparam i23_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n42579), .I1(\data_out_frame[18] [2]), .I2(n42515), 
            .I3(n44671), .O(n72));
    defparam i30_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i19920_4_lut (.I0(n8_adj_4630), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n26414), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i19920_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i28_4_lut (.I0(\data_out_frame[24] [4]), .I1(n42458), .I2(\data_out_frame[17] [7]), 
            .I3(n42956), .O(n70));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n42923), .I1(n42616), .I2(n42687), .I3(n42610), 
            .O(n71));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1482 (.I0(n4452), .I1(n26494), .I2(n23516), .I3(GND_net), 
            .O(n3_adj_4620));
    defparam i1_3_lut_adj_1482.LUT_INIT = 16'h1010;
    SB_LUT4 i27_4_lut (.I0(\data_out_frame[17] [1]), .I1(n42599), .I2(\data_out_frame[17] [4]), 
            .I3(n42417), .O(n69));
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1483 (.I0(n39836), .I1(n42584), .I2(\data_in_frame[14] [4]), 
            .I3(n42524), .O(n42811));
    defparam i1_2_lut_4_lut_adj_1483.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1484 (.I0(n42637), .I1(\data_in_frame[11] [4]), 
            .I2(n42862), .I3(n42881), .O(n6_adj_4438));
    defparam i1_2_lut_4_lut_adj_1484.LUT_INIT = 16'h6996;
    SB_LUT4 i15018_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n28532));
    defparam i15018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_2_lut_4_lut (.I0(n26912), .I1(n39506), .I2(n26989), .I3(n26531), 
            .O(n11));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1485 (.I0(n40613), .I1(n42587), .I2(n26025), 
            .I3(\data_in_frame[18] [5]), .O(n40620));
    defparam i1_2_lut_4_lut_adj_1485.LUT_INIT = 16'h9669;
    SB_LUT4 i38_4_lut (.I0(n65), .I1(n67), .I2(n66), .I3(n68), .O(n80));
    defparam i38_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut (.I0(n40489), .I1(\data_out_frame[25] [6]), .I2(n42293), 
            .I3(\data_out_frame[15] [5]), .O(n73));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1486 (.I0(\FRAME_MATCHER.state_c [31]), .I1(n6_adj_4641), 
            .I2(GND_net), .I3(GND_net), .O(n41649));
    defparam i1_2_lut_adj_1486.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1487 (.I0(n26912), .I1(n39506), .I2(\data_out_frame[15] [1]), 
            .I3(n40489), .O(n40485));
    defparam i1_2_lut_3_lut_4_lut_adj_1487.LUT_INIT = 16'h9669;
    SB_LUT4 i39_4_lut (.I0(n69), .I1(n71), .I2(n70), .I3(n72), .O(n81));
    defparam i39_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i41_4_lut (.I0(n81), .I1(n73), .I2(n80), .I3(n74), .O(n40583));
    defparam i41_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1488 (.I0(\data_out_frame[15] [4]), .I1(n39506), 
            .I2(n27374), .I3(GND_net), .O(n39580));
    defparam i2_3_lut_adj_1488.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33649 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n48820));
    defparam byte_transmit_counter_0__bdd_4_lut_33649.LUT_INIT = 16'he4aa;
    SB_LUT4 i15019_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n28533));
    defparam i15019_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15020_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n28534));
    defparam i15020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15021_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n28535));
    defparam i15021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15022_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n28536));
    defparam i15022_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15023_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n28537));
    defparam i15023_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1489 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[17] [6]), 
            .I2(n42627), .I3(n39580), .O(n44671));
    defparam i3_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(n44671), .I1(n42536), .I2(GND_net), 
            .I3(GND_net), .O(n42537));
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1491 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[24] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42971));
    defparam i1_2_lut_adj_1491.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(\data_out_frame[22] [4]), .I1(\data_out_frame[22] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42929));
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h6666;
    SB_LUT4 i15024_3_lut_4_lut (.I0(n8_adj_4469), .I1(n42274), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n28538));
    defparam i15024_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15233_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n28747));
    defparam i15233_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_adj_1493 (.I0(n42652), .I1(n39584), .I2(n42929), 
            .I3(GND_net), .O(n8_adj_4672));
    defparam i3_3_lut_adj_1493.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1494 (.I0(\data_out_frame[25] [0]), .I1(n42503), 
            .I2(n8_adj_4672), .I3(n42820), .O(n42299));
    defparam i1_4_lut_adj_1494.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1495 (.I0(n39652), .I1(n42299), .I2(\data_out_frame[25] [1]), 
            .I3(GND_net), .O(n44708));
    defparam i2_3_lut_adj_1495.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1496 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n42481));
    defparam i1_2_lut_adj_1496.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_33654 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n48826));
    defparam byte_transmit_counter_0__bdd_4_lut_33654.LUT_INIT = 16'he4aa;
    SB_LUT4 i15234_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n28748));
    defparam i15234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_adj_1497 (.I0(n40525), .I1(\data_out_frame[18] [1]), 
            .I2(n39685), .I3(GND_net), .O(n14_adj_4673));
    defparam i5_3_lut_adj_1497.LUT_INIT = 16'h6969;
    SB_LUT4 i15235_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n28749));
    defparam i15235_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1498 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[13] [6]), 
            .I2(n42481), .I3(n42696), .O(n15_adj_4674));
    defparam i6_4_lut_adj_1498.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1499 (.I0(n15_adj_4674), .I1(n42477), .I2(n14_adj_4673), 
            .I3(n27309), .O(n42536));
    defparam i8_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i15236_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n28750));
    defparam i15236_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15237_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n28751));
    defparam i15237_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15238_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n28752));
    defparam i15238_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1500 (.I0(\data_out_frame[20] [3]), .I1(n42536), 
            .I2(GND_net), .I3(GND_net), .O(n42932));
    defparam i1_2_lut_adj_1500.LUT_INIT = 16'h6666;
    SB_LUT4 i15239_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n28753));
    defparam i15239_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15240_3_lut_4_lut (.I0(n8_adj_4644), .I1(n42281), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n28754));
    defparam i15240_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1501 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42274), .I3(\FRAME_MATCHER.i [0]), .O(n42277));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1501.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1502 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42260), .I3(\FRAME_MATCHER.i [0]), .O(n42264));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1502.LUT_INIT = 16'hfdff;
    SB_LUT4 equal_301_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4644));   // verilog/coms.v(154[7:23])
    defparam equal_301_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(\data_out_frame[18] [2]), .I1(n39625), 
            .I2(GND_net), .I3(GND_net), .O(n40455));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1504 (.I0(\data_out_frame[20] [5]), .I1(n42932), 
            .I2(\data_out_frame[24] [7]), .I3(n27252), .O(n42820));
    defparam i3_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n42610));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1506 (.I0(n42935), .I1(n39859), .I2(n42820), 
            .I3(n40455), .O(n14_adj_4675));
    defparam i6_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1507 (.I0(n43547), .I1(n14_adj_4675), .I2(n10_adj_4616), 
            .I3(\data_out_frame[18] [4]), .O(n39652));
    defparam i7_4_lut_adj_1507.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1508 (.I0(n39652), .I1(n42610), .I2(n40510), 
            .I3(GND_net), .O(n43687));
    defparam i2_3_lut_adj_1508.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1509 (.I0(\data_out_frame[15] [6]), .I1(n42741), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4676));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1509.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1510 (.I0(n39506), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[16] [0]), .I3(n6_adj_4676), .O(n40258));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1511 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n42281), .I3(\FRAME_MATCHER.i [0]), .O(n42285));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1511.LUT_INIT = 16'hfdff;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[22] [2]), .I2(\data_out_frame[23] [2]), 
            .I3(byte_transmit_counter[1]), .O(n48850));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1512 (.I0(\data_out_frame[20] [4]), .I1(\data_out_frame[23] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42935));
    defparam i1_2_lut_adj_1512.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1513 (.I0(\data_out_frame[18] [2]), .I1(n40258), 
            .I2(GND_net), .I3(GND_net), .O(n42823));
    defparam i1_2_lut_adj_1513.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1514 (.I0(\data_out_frame[16] [1]), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[16] [3]), .I3(GND_net), .O(n42968));
    defparam i1_2_lut_3_lut_adj_1514.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1515 (.I0(\data_out_frame[10] [7]), .I1(n42959), 
            .I2(\data_out_frame[9] [1]), .I3(n27188), .O(n6_adj_4417));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_4_lut_adj_1515.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1516 (.I0(n42823), .I1(\data_out_frame[22] [6]), 
            .I2(\data_out_frame[23] [1]), .I3(\data_out_frame[20] [5]), 
            .O(n14_adj_4677));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1516.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1517 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[21][2] ), 
            .O(n9));
    defparam i1_2_lut_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1518 (.I0(n42935), .I1(n14_adj_4677), .I2(n10_adj_4643), 
            .I3(\data_out_frame[20] [6]), .O(n40510));   // verilog/coms.v(78[16:27])
    defparam i7_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1519 (.I0(n40510), .I1(n44349), .I2(GND_net), 
            .I3(GND_net), .O(n39510));
    defparam i1_2_lut_adj_1519.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_4_lut_adj_1520 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[8] [6]), .O(n27558));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4678));
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1522 (.I0(n42844), .I1(n42599), .I2(n42856), 
            .I3(n6_adj_4678), .O(n39625));
    defparam i4_4_lut_adj_1522.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1523 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n42893));
    defparam i1_2_lut_3_lut_adj_1523.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1524 (.I0(n40632), .I1(\data_out_frame[20] [5]), 
            .I2(n42772), .I3(n6_adj_4617), .O(n44349));
    defparam i4_4_lut_adj_1524.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1525 (.I0(\data_out_frame[25] [3]), .I1(\data_out_frame[25] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42515));
    defparam i1_2_lut_adj_1525.LUT_INIT = 16'h6666;
    SB_LUT4 i13_3_lut_4_lut (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[4] [6]), .O(n38_adj_4583));   // verilog/coms.v(74[16:27])
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 select_658_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n3846), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4597));
    defparam select_658_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1526 (.I0(n24648), .I1(n42515), .I2(n44349), 
            .I3(GND_net), .O(n43493));
    defparam i2_3_lut_adj_1526.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1527 (.I0(\data_out_frame[21][0] ), .I1(n39586), 
            .I2(n40632), .I3(\data_out_frame[23] [3]), .O(n24648));
    defparam i2_3_lut_4_lut_adj_1527.LUT_INIT = 16'h9669;
    SB_LUT4 i20334_1_lut (.I0(n33835), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_4633));
    defparam i20334_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_3_lut_adj_1528 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[20] [6]), 
            .I2(n42503), .I3(GND_net), .O(n40632));
    defparam i1_2_lut_3_lut_adj_1528.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1529 (.I0(n26722), .I1(n42689), .I2(n42293), 
            .I3(n42856), .O(n10_adj_4635));
    defparam i4_4_lut_adj_1529.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1530 (.I0(n4_adj_4636), .I1(n42248), .I2(n31), 
            .I3(\FRAME_MATCHER.state_c [1]), .O(n44019));
    defparam i3_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1531 (.I0(n44481), .I1(\data_out_frame[18] [4]), 
            .I2(\data_out_frame[18] [6]), .I3(n43849), .O(n42503));
    defparam i3_4_lut_adj_1531.LUT_INIT = 16'h6996;
    uart_tx tx (.r_Bit_Index({Open_32, Open_33, \r_Bit_Index[0] }), .GND_net(GND_net), 
            .n27840(n27840), .r_SM_Main({r_SM_Main}), .n28123(n28123), 
            .\r_SM_Main_2__N_3616[0] (\r_SM_Main_2__N_3616[0] ), .\r_SM_Main_2__N_3613[1] (\r_SM_Main_2__N_3613[1] ), 
            .CLK_c(CLK_c), .tx_o(tx_o), .tx_data({tx_data}), .VCC_net(VCC_net), 
            .n28387(n28387), .n28235(n28235), .tx_active(tx_active), .n18934(n18934), 
            .n4(n4), .n48874(n48874), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.\r_Bit_Index[0] (\r_Bit_Index[0]_adj_3 ), .GND_net(GND_net), 
            .n27844(n27844), .r_SM_Main({r_SM_Main_adj_10}), .n28125(n28125), 
            .CLK_c(CLK_c), .\r_SM_Main_2__N_3542[2] (\r_SM_Main_2__N_3542[2] ), 
            .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), .n4(n4_adj_7), .n4_adj_1(n4_adj_8), 
            .VCC_net(VCC_net), .n4_adj_2(n4_adj_9), .n26398(n26398), .n26390(n26390), 
            .n33332(n33332), .n28431(n28431), .n41875(n41875), .rx_data_ready(rx_data_ready), 
            .n28203(n28203), .rx_data({rx_data}), .n28201(n28201), .n28200(n28200), 
            .n28199(n28199), .n28198(n28198), .n28197(n28197), .n28196(n28196), 
            .n42166(n42166), .n28437(n28437)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (r_Bit_Index, GND_net, n27840, r_SM_Main, n28123, \r_SM_Main_2__N_3616[0] , 
            \r_SM_Main_2__N_3613[1] , CLK_c, tx_o, tx_data, VCC_net, 
            n28387, n28235, tx_active, n18934, n4, n48874, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output [2:0]r_Bit_Index;
    input GND_net;
    output n27840;
    output [2:0]r_SM_Main;
    output n28123;
    input \r_SM_Main_2__N_3616[0] ;
    output \r_SM_Main_2__N_3613[1] ;
    input CLK_c;
    output tx_o;
    input [7:0]tx_data;
    input VCC_net;
    input n28387;
    input n28235;
    output tx_active;
    output n18934;
    output n4;
    input n48874;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n45869, n45870, n45873, n45872;
    wire [2:0]r_Bit_Index_c;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]n307;
    
    wire n33888, n21050, n21051, o_Tx_Serial_N_3644, n3;
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n28017, n38379, n38378, n38377, n38376, n38375, n38374, 
        n38373, n25940, n38372, n48718, n3_adj_4404, n44061, n10;
    
    SB_LUT4 i30738_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45869));
    defparam i30738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30739_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45870));
    defparam i30739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30742_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45873));
    defparam i30742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30741_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n45872));
    defparam i30741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2363_3_lut (.I0(r_Bit_Index_c[2]), .I1(r_Bit_Index_c[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i2363_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i14609_3_lut (.I0(n27840), .I1(n33888), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28123));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14609_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2356_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i2356_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n33888));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7660_4_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(n33888), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3613[1] ), .O(n21050));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7660_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7661_3_lut (.I0(n21050), .I1(\r_SM_Main_2__N_3613[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n21051));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7661_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3644), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFESR r_Clock_Count_2201__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n1), 
            .D(n41[1]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n1), 
            .D(n41[2]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n1), 
            .D(n41[3]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n1), 
            .D(n41[4]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n1), 
            .D(n41[5]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n1), 
            .D(n41[6]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n1), 
            .D(n41[7]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_2201__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n1), 
            .D(n41[8]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 r_Clock_Count_2201_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n38379), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2201_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n38378), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_9 (.CI(n38378), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n38379));
    SB_LUT4 r_Clock_Count_2201_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n38377), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_8 (.CI(n38377), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n38378));
    SB_LUT4 r_Clock_Count_2201_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n38376), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_7 (.CI(n38376), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n38377));
    SB_LUT4 r_Clock_Count_2201_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n38375), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_6 (.CI(n38375), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n38376));
    SB_LUT4 r_Clock_Count_2201_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n38374), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_5 (.CI(n38374), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n38375));
    SB_LUT4 r_Clock_Count_2201_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n38373), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n25940), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n21051), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_CARRY r_Clock_Count_2201_add_4_4 (.CI(n38373), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n38374));
    SB_LUT4 r_Clock_Count_2201_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n38372), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_3 (.CI(n38372), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n38373));
    SB_LUT4 r_Clock_Count_2201_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2201_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2201_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n38372));
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(CLK_c), .E(n27840), 
            .D(n307[1]), .R(n28123));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(CLK_c), .E(n27840), 
            .D(n307[2]), .R(n28123));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_2201__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n1), 
            .D(n41[0]), .R(n28017));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index_c[1]), .I1(n45872), 
            .I2(n45873), .I3(r_Bit_Index_c[2]), .O(n48718));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n48718_bdd_4_lut (.I0(n48718), .I1(n45870), .I2(n45869), .I3(r_Bit_Index_c[2]), 
            .O(o_Tx_Serial_N_3644));
    defparam n48718_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n28387));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n28235));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i5553_2_lut (.I0(\r_SM_Main_2__N_3616[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n18934));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5553_2_lut.LUT_INIT = 16'h2222;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4404), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n25940), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n25940), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n25940), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n25940), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n25940), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n25940), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n25940), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[3]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[2]), .O(n44061));
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[5]), .I2(n44061), 
            .I3(r_Clock_Count[8]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[6]), .I1(n10), .I2(r_Clock_Count[7]), 
            .I3(GND_net), .O(\r_SM_Main_2__N_3613[1] ));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i32705_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3613[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n28017));
    defparam i32705_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n48874));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3613[1] ), .O(n27840));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3616[0] ), 
            .I3(r_SM_Main[1]), .O(n25940));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i9721_2_lut_3_lut (.I0(\r_SM_Main_2__N_3613[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4404));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i9721_2_lut_3_lut.LUT_INIT = 16'h7878;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (\r_Bit_Index[0] , GND_net, n27844, r_SM_Main, n28125, 
            CLK_c, \r_SM_Main_2__N_3542[2] , r_Rx_Data, RX_N_10, n4, 
            n4_adj_1, VCC_net, n4_adj_2, n26398, n26390, n33332, 
            n28431, n41875, rx_data_ready, n28203, rx_data, n28201, 
            n28200, n28199, n28198, n28197, n28196, n42166, n28437) /* synthesis syn_module_defined=1 */ ;
    output \r_Bit_Index[0] ;
    input GND_net;
    output n27844;
    output [2:0]r_SM_Main;
    output n28125;
    input CLK_c;
    output \r_SM_Main_2__N_3542[2] ;
    output r_Rx_Data;
    input RX_N_10;
    output n4;
    output n4_adj_1;
    input VCC_net;
    output n4_adj_2;
    output n26398;
    output n26390;
    output n33332;
    input n28431;
    input n41875;
    output rx_data_ready;
    input n28203;
    output [7:0]rx_data;
    input n28201;
    input n28200;
    input n28199;
    input n28198;
    input n28197;
    input n28196;
    input n42166;
    input n28437;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]n326;
    
    wire n33882;
    wire [7:0]n37;
    
    wire n27778;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n28026, n33968;
    wire [2:0]r_SM_Main_2__N_3548;
    
    wire n1, n3, r_Rx_Data_R, n46844, n38371, n38370, n38369, 
        n38368, n33898, n38367, n38366, n38365, n26318, n45668, 
        n26292, n6, n46896, n46894, n6_adj_4403;
    
    SB_LUT4 i2341_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i2341_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i14611_3_lut (.I0(n27844), .I1(n33882), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28125));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14611_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2334_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i2334_2_lut.LUT_INIT = 16'h6666;
    SB_DFFESR r_Clock_Count_2199__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n27778), 
            .D(n37[1]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n27778), 
            .D(n37[2]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n27778), 
            .D(n37[3]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n27778), 
            .D(n37[4]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n27778), 
            .D(n37[5]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_2199__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n27778), 
            .D(n37[6]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n33882));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_DFFESR r_Clock_Count_2199__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n27778), 
            .D(n37[7]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n33882), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n33968));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n33968), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n27844), 
            .D(n326[1]), .R(n28125));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_334_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_334_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n27844), 
            .D(n326[2]), .R(n28125));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 equal_332_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_332_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i31799_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3548[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n46844));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i31799_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_Clock_Count_2199_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n38371), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_2199_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n38370), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_8 (.CI(n38370), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n38371));
    SB_LUT4 r_Clock_Count_2199_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n38369), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_7 (.CI(n38369), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n38370));
    SB_LUT4 r_Clock_Count_2199_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n38368), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n46844), .I1(\r_SM_Main_2__N_3542[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n33898));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_CARRY r_Clock_Count_2199_add_4_6 (.CI(n38368), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n38369));
    SB_LUT4 r_Clock_Count_2199_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n38367), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_5 (.CI(n38367), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n38368));
    SB_LUT4 r_Clock_Count_2199_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n38366), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_4 (.CI(n38366), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n38367));
    SB_LUT4 r_Clock_Count_2199_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n38365), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_3 (.CI(n38365), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n38366));
    SB_LUT4 r_Clock_Count_2199_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_2199_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_2199_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n38365));
    SB_LUT4 equal_330_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_330_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut (.I0(n26318), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n26398));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR r_Clock_Count_2199__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n27778), 
            .D(n37[0]), .R(n28026));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i1_2_lut_adj_861 (.I0(n26318), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n26390));
    defparam i1_2_lut_adj_861.LUT_INIT = 16'hbbbb;
    SB_LUT4 i19834_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33332));
    defparam i19834_2_lut.LUT_INIT = 16'h8888;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(CLK_c), .D(n28431));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n41875));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n28203));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n28201));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n28200));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n28199));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n33898), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n28198));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n28197));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n28196));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n42166));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i4_4_lut (.I0(n45668), .I1(n26292), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[1]), .O(r_SM_Main_2__N_3548[0]));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20381_4_lut (.I0(r_Clock_Count[0]), .I1(n26292), .I2(n6), 
            .I3(r_Clock_Count[1]), .O(\r_SM_Main_2__N_3542[2] ));
    defparam i20381_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i30636_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(GND_net), .I3(GND_net), .O(n45668));
    defparam i30636_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[5]), .O(n26292));   // verilog/uart_rx.v(68[17:52])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i31998_4_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[1]), .I2(n26292), 
            .I3(r_Clock_Count[3]), .O(n46896));
    defparam i31998_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i32006_3_lut (.I0(n46896), .I1(r_SM_Main[0]), .I2(n45668), 
            .I3(GND_net), .O(n46894));
    defparam i32006_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n46894), .I2(\r_SM_Main_2__N_3542[2] ), 
            .I3(r_SM_Main[1]), .O(n28026));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_2_lut_adj_862 (.I0(r_SM_Main_2__N_3548[0]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4403));
    defparam i2_2_lut_adj_862.LUT_INIT = 16'h4444;
    SB_LUT4 i32694_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4403), 
            .I3(r_Rx_Data), .O(n27778));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i32694_4_lut.LUT_INIT = 16'h4555;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n28437));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3542[2] ), .O(n26318));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3542[2] ), .O(n27844));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    
endmodule
