// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Fri Jan 31 00:11:14 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(122[22:39])
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(123[21:45])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(125[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(126[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(127[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(128[22:24])
    
    wire n4;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(130[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(131[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(132[22:35])
    
    wire n28284, n28118, n28283;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(162[22:33])
    
    wire n27990, n33251, n5629, n5630;
    wire [7:0]data;   // verilog/TinyFPGA_B.v(206[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(230[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(238[15:20])
    wire [22:0]pwm_setpoint_22__N_11;
    
    wire RX_N_10;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n4_adj_4865;
    wire [31:0]motor_state_23__N_82;
    wire [25:0]encoder0_position_scaled_23__N_34;
    wire [23:0]displacement_23__N_58;
    
    wire n28282, n587, n588, n589, n590, n591, n592, n593, n594, 
        n595, n596, n597, n598, n599, n600, n601, n602, n603, 
        n604, n605, n606, n607, n608, n609, n610, n611, n612, 
        n613, n614, n615, n616, n617, n618, n619, n18735, n18734, 
        n18733, n18732, n18731, n18730, n18729, \ID_READOUT_FSM.state_2__N_207 , 
        n36603;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n27903, n33396, n28117, n18728, n18727, n7, n4_adj_4866, 
        n18726, n28281, n27989, n18725, n18724, n18723, n18722, 
        n18721, n18720, n18719, n18718, n18717, n18716, n18715, 
        n18714, n18713, n28116, n28280, n28279, n28278, n1, n28115, 
        n28277, n28276, n28275, n28114, n27902, n27988, n28274, 
        n18712, n36784, n36788, n27987, n28273, n24676, n27746, 
        n24674, n36714, n27901, n27658, n28113, n15, n27986, n27642, 
        n18703, n18702, n18701, n18700, n18699, n18698, n18697, 
        n18696, n28112, n28272, n27985, n28111, n28271, n20, n36733, 
        n425, n18693, n18692, n18, n27657;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n28110, n15_adj_4867, n24712, n28270, n28269, n16, n23704, 
        n3, n4_adj_4868, n5, n6, n7_adj_4869, n8, n9, n10, n11, 
        n12, n13, n14, n15_adj_4870, n16_adj_4871, n17, n18_adj_4872, 
        n19, n20_adj_4873, n21, n22, n23, n24, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n28109, n27641, n10125, n27984, n28108, n28268;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n34118, n123, n37, n36, n30, n29, n28, n27, n26, 
        n25_adj_4874, n36620, n24_adj_4875, n23_adj_4876, n22_adj_4877, 
        n21_adj_4878, n34, n33, n32, n31, n30_adj_4879, n7_adj_4880, 
        n28267, n37939, n28107, n27983, n17_adj_4881, n28266, n27982, 
        n16_adj_4882, n36615, n16_adj_4883, n12_adj_4884, n10_adj_4885, 
        n36611, n28265, n28264, n37934, n27981, n28106, n28263, 
        n28262, n28261, n28260, n28105, n28104, n27980, n27979, 
        n27978, n28103, n28259, n27745, n27977, n28258, n28257, 
        n28256, n28255, n28102, n28101, n28254, n28100, n27976, 
        n28099, n36605, n27744, n28253, n28252, n28098, n27743, 
        n28097, n28251, n27742, n28250, n28096, n24606, n28249, 
        n28095, n28248, n28247, n28246, n28245, n28094, n28244, 
        n28243, n27741, n28093, n28092, n28091, n28090, n28089, 
        n33723, n28242, n28088, n27656, n27740, n28241, n28240, 
        n28087, n28239, n28086, n24634, n28085, n24570, n28084, 
        n27640, n28238, n24624, n27739, n24622, n28237, n27738, 
        n27737, n23776, n24616, n28236, n28235, n36550, n27736, 
        n27735, n28234, n27734, n28233, n5_adj_4886, n28232, n27733, 
        n27732, n36468, n26386, n28231, n28230, n28229, n28075, 
        n28228, n28074, n28227, n27731, n36470, n27730, n28073, 
        n27655, n28226, n28072, n28225, n28224, n28223, n28071, 
        n28070, n28222, n27729, n28221, n28069, n28220, n28068, 
        n28067, n28066, n28219, n27728, n28218, n3303, n28217, 
        n30964, n31596, n4452, n33948, n28216, n28065, n28215, 
        n31590, n66, n27654, n28214, n28064, n28213, n27639, n36300, 
        n22_adj_4887, n20_adj_4888, n18_adj_4889, n13_adj_4890, n28212, 
        n28211, n28063, n24596, n28210, n28209, n14_adj_4891, n10_adj_4892, 
        n28062, n4_adj_4893, n28061, n18691, n18690, n18689, \FRAME_MATCHER.i_31__N_2461 , 
        n36789, n35957, n7_adj_4894, n35956, n35954, n24470, n28208, 
        n32395, n28060, n24425, n24181, n24598, n19204, n19202, 
        n19201, n19200, n19199, n19198, n19197, n19194, n19193, 
        n19192, n19191, n19190, n19189, n19188, n28207, n19185, 
        n28059, n24688, n30803, n19175, n19174, n19173, n19172, 
        n19171, n19170, n19169, n19168, n19167, n19166, n19165, 
        n19164, n19163, n19162, n19161, n19160, n19159, n19158, 
        n19157, n19156, n19155, n19154, n19153, n19152, n19151, 
        n19149, n19148, n19147, n19146, n19145, n19144, n18688, 
        n1172, n18687, n18686, n18685, n18684, n18683, n18682, 
        n18681, n18680, n18679, n18678, n18677, n18676, n18675, 
        n18674, n25_adj_4895, n24_adj_4896, n23_adj_4897, n22_adj_4898, 
        n21_adj_4899, n20_adj_4900, n19_adj_4901, n18_adj_4902, n17_adj_4903, 
        n16_adj_4904, n15_adj_4905, n14_adj_4906, n13_adj_4907, n12_adj_4908, 
        n11_adj_4909, n10_adj_4910, n9_adj_4911, n8_adj_4912, n7_adj_4913, 
        n6_adj_4914, n5_adj_4915, n4_adj_4916, n3_adj_4917, n2, n18673, 
        n19143, n3568, n19142, n19141, n28058, n19140, n19139, 
        n19138, n19137, n19136, n18672, n19135, n19134, n19133, 
        n28206, n19132, n19131, n19130, n19129, n19128, n19127, 
        n19126, n19125, n19124, n19123, n19122, n19121, n19120, 
        n19119, n19118, n19117, n19116, n19115, n19114, n19113, 
        n6_adj_4918, n19112, n19111, n19110, n19109, n19108, n19107, 
        n19106, n19105, n19104, n19103, n5_adj_4919, n19102, n19101, 
        n19100, n19099, n19098, n19097, n19096, n19095, n19094, 
        n19093, n19092, n19091, n6_adj_4920, n19090, n19089, n19088, 
        n19087, n19086, n19085, n19084, n4_adj_4921, n19083, n19082, 
        n19081, n19080, n19079, n19078, n19077, n19076, n28205, 
        n19075, n19074, n19073, n19072, n19071, n19070, n19069, 
        n19068, n19067, n19066, n19065, n19064, n19063, n19062, 
        n19061, n19060, n19059, n19058, n19057, n19056, n28057, 
        n28204, n28203, n28202, n27653, n27652, n19055, n19054, 
        n5627, n19053, n19052, n19051, n19050, n19049, n19048, 
        n19047, n19046, n5631, n19045, n19044, n19043, n19042, 
        n19041, n19040, n19039, n19038, n19037, n19036, n19035, 
        n19034, n19033, n19032, quadA_debounced, quadB_debounced, 
        n19031, n19030, n19029, n19028, n19027, n5632, n19026, 
        n19025, n19024, n19023, n19022, n19021, n19020, n19019, 
        quadA_debounced_adj_4922, quadB_debounced_adj_4923, n35924, n19018, 
        n19017, n19016, n19015, n19014, n19013, n18671, n19012, 
        n36787, n19011, n19010, n5131, n19009, n19008, rw;
    wire [7:0]state_adj_5104;   // verilog/eeprom.v(23[11:16])
    
    wire n19007, n19006, n19005, n19004, n19003, n19002, n19001, 
        n10_adj_4926, n19000, n2134, n4_adj_4927, n18999, n18998, 
        n18997, n32403, n18996, n18995, n18994, n18993, n18992, 
        n18991, n18990, n18989, n18988, n18987, n18986, n18985, 
        n18984, n18983, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n28201, n18982, n18981, n18980, n18979, n18978, n18977, 
        n18976, n18975, n18974, n18973, n18972, n18971, n18970, 
        n18969, n18968, n18670, n18967;
    wire [2:0]r_SM_Main_2__N_3379;
    
    wire n18966, n18965, n18964, n18669, n18963, n15_adj_4928, n18962, 
        n18961, n18960, n18959, n18958, n18957, n18956, n18955, 
        n18954, n18953, n18952, n18951, n18950, n18949, n18948;
    wire [2:0]r_SM_Main_adj_5111;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5113;   // verilog/uart_tx.v(33[16:27])
    
    wire n28056, n28055, n18947;
    wire [2:0]r_SM_Main_2__N_3450;
    
    wire n18946, n18945, n28200, n18944, n18943, n18942, n18941, 
        n28199, n18940, n18939, n18938, n18937, n18936, n18935, 
        n28198, n28054, n28197, n28196, n28195, n27651, n18934, 
        n18933, n18932, n18931, n18930, n18929, n18928, n18927, 
        n18926, n18925, n18924, n18923, n18922, n16906;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n18921, n5300, n18920, n18919;
    wire [1:0]reg_B_adj_5120;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n18918, n18917, n18916, n28053, n18915, n18914;
    wire [7:0]state_adj_5132;   // verilog/i2c_controller.v(33[12:17])
    
    wire n28052;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n18913, n18912, enable_slow_N_3964, n18911, n15_adj_4936, 
        n18910, n28194, n18909, n18908;
    wire [7:0]state_7__N_3861;
    
    wire n18907, n18906, n18668, n4867, n18905, n28051, n28050, 
        n18904;
    wire [7:0]state_7__N_3877;
    
    wire n18903, n17027, n18902, n18901, n18900, n18899, n18898, 
        n18897, n18896, n28193, n28192, n28191, n28049, n28048, 
        n18895, n18667, n18666, n18665, n18664, n18663, n18660, 
        n18894, n18893, n18892, n18891, n18890, n18889, n18888, 
        n18887, n18886, n18885, n18884, n18883, n18882, n18881, 
        n18880, n18879, n18878, n18877, n18876, n18875, n18874, 
        n18866, n18865, n18864, n18863, n18862, n18861, n18860, 
        n18859, n3_adj_4937, n5_adj_4938, n6_adj_4939, n7_adj_4940, 
        n8_adj_4941, n9_adj_4942, n10_adj_4943, n11_adj_4944, n12_adj_4945, 
        n13_adj_4946, n14_adj_4947, n15_adj_4948, n16_adj_4949, n17_adj_4950, 
        n18_adj_4951, n19_adj_4952, n20_adj_4953, n21_adj_4954, n22_adj_4955, 
        n23_adj_4956, n24_adj_4957, n25_adj_4958, n18850, n28190, 
        n28189, n509, n510, n511, n513, n515, n516, n517, n518, 
        n519, n521, n523, n598_adj_4959, n619_adj_4960, n18849, 
        n18848, n18847, n674, n675, n676, n677, n678, n679, 
        n700, n18846, n728, n729, n730, n731, n732, n733, n752, 
        n753, n754, n755, n756, n757, n758, n18845, n763, n765, 
        n767, n768, n769, n770, n771, n772, n773, n774, n775, 
        n778, n18844, n806, n807, n808, n809, n810, n811, n812, 
        n830, n831, n832, n833, n834, n835, n836, n837, n856, 
        n883, n884, n885, n886, n887, n888, n889, n890, n891, 
        n18843, n28188, n908, n909, n910, n911, n912, n913, 
        n914, n915, n916, n934, n961, n962, n963, n964, n965, 
        n966, n967, n968, n969, n970, n986, n987, n988, n989, 
        n990, n991, n992, n993, n994, n995, n28047, n33837, 
        n28187, n1012, n1039, n1040, n1041, n1042, n1043, n1044, 
        n1045, n1046, n1047, n1048, n1049, n1064, n1065, n1066, 
        n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
        n1090, n30832, n1117, n1118, n1119, n1120, n1121, n1122, 
        n1123, n1124, n1125, n1126, n1127, n1128, n1142, n1143, 
        n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, 
        n1152, n1153, n1168, n18336, n1195, n1196, n1197, n1198, 
        n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
        n1207, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
        n1227, n1228, n1229, n1230, n1231, n1232, n1246, n1273, 
        n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, 
        n1282, n1283, n1284, n1285, n1286, n1298, n1299, n1300, 
        n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
        n1309, n1310, n1311, n1324, n1351, n1352, n1353, n1354, 
        n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
        n1363, n1364, n1365, n1376, n1377, n1378, n1379, n1380, 
        n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
        n1389, n1390, n1402, n1429, n1430, n1431, n1432, n1433, 
        n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
        n1442, n1443, n1444, n1454, n1455, n1456, n1457, n1458, 
        n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
        n1467, n1468, n1469, n1480, n1507, n1508, n1509, n1510, 
        n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
        n1519, n1520, n1521, n1522, n1523, n1532, n1533, n1534, 
        n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
        n1543, n1544, n1545, n1546, n1547, n1548, n1558, n1585, 
        n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, 
        n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, 
        n1602, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
        n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, 
        n1625, n1626, n1627, n1636, n1663, n1664, n1665, n1666, 
        n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, 
        n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1688, 
        n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
        n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
        n1705, n1706, n1714, n1741, n1742, n1743, n1744, n1745, 
        n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, 
        n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1766, 
        n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
        n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
        n1783, n1784, n1785, n1792, n32394, n1819, n1820, n1821, 
        n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
        n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, 
        n1838, n1839, n1844, n1845, n1846, n1847, n1848, n1849, 
        n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, 
        n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1870, 
        n28186, n32166, n1897, n1898, n1899, n1900, n1901, n1902, 
        n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, 
        n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
        n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
        n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, 
        n1938, n1939, n1940, n1941, n1942, n1943, n1948, n1975, 
        n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, 
        n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, 
        n1992, n1993, n1994, n1995, n1996, n1997, n2000, n2001, 
        n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
        n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
        n2018, n2019, n2020, n2021, n2022, n2026, n4_adj_4961, 
        n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
        n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, 
        n2069, n2070, n2071, n2073, n2076, n4_adj_4962, n37245, 
        n24710, n35900, n28185, n5826, n5825, n5824, n5823, n5822, 
        n5821, n5820, n5819, n5818, n5817, n5816, n5815, n5814, 
        n5813, n5812, n5811, n5810, n5809, n5808, n5806, n5805, 
        n18489, n26_adj_4963, n32_adj_4964, n56, n16908, n36290, 
        n18223, n18590, n18834, n18833, n18832, n18831, n18830, 
        n18163, n63, n28184, n1_adj_4965, n18652, n10_adj_4966, 
        n28046, n36544, n4_adj_4967, n6_adj_4968, n7_adj_4969, n8_adj_4970, 
        n9_adj_4971, n10_adj_4972, n11_adj_4973, n12_adj_4974, n13_adj_4975, 
        n15_adj_4976, n17_adj_4977, n19_adj_4978, n21_adj_4979, n36621, 
        n23_adj_4980, n25_adj_4981, n27_adj_4982, n36619, n29_adj_4983, 
        n30_adj_4984, n31_adj_4985, n33_adj_4986, n35, n32397, n28183, 
        n28182, n28045, n28181, n28180, n28179, n28044, n35881, 
        n35879, n28178, n28043, n14_adj_4987, n36713, n9_adj_4988, 
        n18829, n18828, n18827, n32413, n8_adj_4989, n7_adj_4990, 
        n36945, n18651, n18650, n18649, n18648, n18647, n18646, 
        n18645, n18644, n18643, n18802, n18801, n18641, n18640, 
        n18639, n18637, n18636, n18635, n18800, n18799, n18798, 
        n18797, n18796, n18795, n34304, n18786, n18785, n18784, 
        n18783, n18782, n18781, n18780, n18779, n18770, n18769, 
        n18768, n18767, n18766, n18765, n18764, n18763, n24_adj_4991, 
        n34934, n21_adj_4992, n20_adj_4993, n17_adj_4994, n32404, 
        n28177, n28042, n28176, n28041, n2_adj_4995, n3_adj_4996, 
        n4_adj_4997, n5_adj_4998, n6_adj_4999, n7_adj_5000, n8_adj_5001, 
        n9_adj_5002, n10_adj_5003, n11_adj_5004, n12_adj_5005, n13_adj_5006, 
        n14_adj_5007, n15_adj_5008, n16_adj_5009, n17_adj_5010, n18_adj_5011, 
        n19_adj_5012, n20_adj_5013, n21_adj_5014, n22_adj_5015, n23_adj_5016, 
        n24_adj_5017, n25_adj_5018, n28040, n24630, n28175, n28039, 
        n28038, n34140, n28037, n28036, n28174, n28035, n28173, 
        n28172, n28171, n33211, n28170, n28169, n28168, n28034, 
        n28167, n28033, n28166, n28032, n28031, n28165, n28164, 
        n28163, n27638, n27650, n28162, n27637, n28161, n27649, 
        n28160, n28021, n28159, n28158, n13_adj_5019, n28157, n23_adj_5020, 
        n27_adj_5021, n29_adj_5022, n28156, n37_adj_5023, n27648, 
        n39, n28155, n43, n45, n49, n28020, n33126, n32402, 
        n33118, n32410, n32409, n33134, n30_adj_5024, n29_adj_5025, 
        n28_adj_5026, n27_adj_5027, n18_adj_5028, n12_adj_5029, n34993, 
        n27636, n32064, n8_adj_5030, n4_adj_5031, n34_adj_5032, n31_adj_5033, 
        n30_adj_5034, n28_adj_5035, n28019, n22_adj_5036, n21_adj_5037, 
        n28018, n24462, n28154, n18634, n18633, n18632, n28017, 
        n28016, n28153, n28152, n18625, n14_adj_5038, n9_adj_5039, 
        n17079, n20_adj_5040, n19_adj_5041, n18_adj_5042, n28151, 
        n17053, n34334, n33924, n28150, n28149, n28315, n33407, 
        n28148, n36013, n36007, n36005, n36001, n35999, n28621, 
        n28620, n28619, n28618, n28617, n28616, n28615, n28614, 
        n28613, n28612, n37310, n28611, n28610, n28609, n28608, 
        n36622, n33787, n7_adj_5043, n28_adj_5044, n27_adj_5045, n26_adj_5046, 
        n25_adj_5047, n28607, n28606, n28605, n28604, n28603, n28602, 
        n6_adj_5048, n34883, n28601, n28600, n28599, n28598, n28147, 
        n6_adj_5049, n5_adj_5050, n28314, n14_adj_5051, n10_adj_5052, 
        n32359, n31970, n28313, n28146, n28145, n4_adj_5053, n28312, 
        n27647, n28144, n28311, n32068, n33160, n28310, n28309, 
        n28143, n27635, n28142, n28141, n28140, n28139, n28308, 
        n28307, n28306, n28138, n28137, n28305, n28136, n27646, 
        n27645, n28304, n28303, n28135, n17084, n24620, n28134, 
        n27749, n28302, n27644, n28133, n27665, n28132, n17058, 
        n32920, n27998, n27664, n27997, n10_adj_5054, n28131, n27748, 
        n27643, n6_adj_5055, n29929, n27663, n28301, n32699, n28300, 
        n27996, n27995, n32722, n14410, n28299, n28130, n27905, 
        n32831, n18626, n28129, n28298, n28297, n28128, n28127, 
        n27994, n27662, n28_adj_5056, n32400, n26_adj_5057, n31374, 
        n24_adj_5058, n28126, n23726, n27993, n32385, n27661, n33450, 
        n19_adj_5059, n16_adj_5060, n28125, n27747, n27660, n28296, 
        n33905, n34465, n27992, n24702, n28124, n28295, n28294, 
        n28123, n28293, n28292, n28291, n12_adj_5061, n28290, n28122, 
        n28289, n28121, n27659, n28120, n28288, n28287, n26_adj_5062, 
        n24_adj_5063, n22_adj_5064, n33114, n28286, n18_adj_5065, 
        n27904, n32658, n28119, n34405, n32412, n27991, n28285;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .data_o({quadA_debounced, quadB_debounced}), 
            .GND_net(GND_net), .n34934(n34934), .reg_B({reg_B}), .VCC_net(VCC_net), 
            .ENCODER0_B_c_0(ENCODER0_B_c_0), .n18641(n18641), .n19175(n19175), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(185[15] 190[4])
    SB_LUT4 i14294_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n34304), 
            .I3(GND_net), .O(n19083));   // verilog/coms.v(127[12] 300[6])
    defparam i14294_3_lut.LUT_INIT = 16'hacac;
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_49 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i30548_1_lut (.I0(n778), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n36945));
    defparam i30548_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_58[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF read_56 (.Q(read), .C(CLK_c), .D(\ID_READOUT_FSM.state_2__N_207 ));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_3877[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i14295_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n34304), 
            .I3(GND_net), .O(n19084));   // verilog/coms.v(127[12] 300[6])
    defparam i14295_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4937));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h2_48 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4868));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    neopixel nx (.GND_net(GND_net), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), .clk32MHz(clk32MHz), 
            .VCC_net(VCC_net), .n6(n6_adj_4918), .n33407(n33407), .\state[0] (state[0]), 
            .\state[1] (state[1]), .start(start), .n5(n5_adj_4919), .n2134(n2134), 
            .timer({timer}), .n4(n4_adj_4961), .n26386(n26386), .LED_c(LED_c), 
            .neopxl_color({neopxl_color}), .n31374(n31374), .n19149(n19149), 
            .n19148(n19148), .n19147(n19147), .n19146(n19146), .n19145(n19145), 
            .n19144(n19144), .n19143(n19143), .n19142(n19142), .n19141(n19141), 
            .n19140(n19140), .n19139(n19139), .n19138(n19138), .n19137(n19137), 
            .n19136(n19136), .n19135(n19135), .n19134(n19134), .n19133(n19133), 
            .n19132(n19132), .n19131(n19131), .n19130(n19130), .n19129(n19129), 
            .n19128(n19128), .n19127(n19127), .n19126(n19126), .n19125(n19125), 
            .n19124(n19124), .n19123(n19123), .n19122(n19122), .n19121(n19121), 
            .n19120(n19120), .n19119(n19119), .NEOPXL_c(NEOPXL_c), .n18625(n18625)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[10] 49[2])
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14296_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n34304), 
            .I3(GND_net), .O(n19085));   // verilog/coms.v(127[12] 300[6])
    defparam i14296_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14297_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n34304), 
            .I3(GND_net), .O(n19086));   // verilog/coms.v(127[12] 300[6])
    defparam i14297_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_9_lut (.I0(n36945), .I1(n752), 
            .I2(VCC_net), .I3(n28037), .O(n830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14298_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n34304), 
            .I3(GND_net), .O(n19087));   // verilog/coms.v(127[12] 300[6])
    defparam i14298_3_lut.LUT_INIT = 16'hacac;
    SB_DFF dir_53 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_23__I_0_add_513_8_lut (.I0(GND_net), .I1(n753), 
            .I2(VCC_net), .I3(n28036), .O(n806)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_8 (.CI(n28036), .I0(n753), 
            .I1(VCC_net), .CO(n28037));
    SB_LUT4 i14299_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19088));   // verilog/coms.v(127[12] 300[6])
    defparam i14299_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_513_7_lut (.I0(GND_net), .I1(n754), 
            .I2(GND_net), .I3(n28035), .O(n807)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_7 (.CI(n28035), .I0(n754), 
            .I1(GND_net), .CO(n28036));
    SB_LUT4 i2_2_lut (.I0(pwm_counter[27]), .I1(pwm_counter[28]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_5052));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14300_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19089));   // verilog/coms.v(127[12] 300[6])
    defparam i14300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14301_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19090));   // verilog/coms.v(127[12] 300[6])
    defparam i14301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[23]), .I1(pwm_counter[29]), .I2(pwm_counter[25]), 
            .I3(pwm_counter[26]), .O(n14_adj_5051));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14302_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19091));   // verilog/coms.v(127[12] 300[6])
    defparam i14302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut (.I0(pwm_counter[30]), .I1(n14_adj_5051), .I2(n10_adj_5052), 
            .I3(pwm_counter[24]), .O(n16906));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14303_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19092));   // verilog/coms.v(127[12] 300[6])
    defparam i14303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14304_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19093));   // verilog/coms.v(127[12] 300[6])
    defparam i14304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14305_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19094));   // verilog/coms.v(127[12] 300[6])
    defparam i14305_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14306_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19095));   // verilog/coms.v(127[12] 300[6])
    defparam i14306_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14307_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19096));   // verilog/coms.v(127[12] 300[6])
    defparam i14307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14308_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19097));   // verilog/coms.v(127[12] 300[6])
    defparam i14308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13896_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n34304), .I3(GND_net), .O(n18685));   // verilog/coms.v(127[12] 300[6])
    defparam i13896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14309_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19098));   // verilog/coms.v(127[12] 300[6])
    defparam i14309_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14310_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19099));   // verilog/coms.v(127[12] 300[6])
    defparam i14310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13897_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n34304), .I3(GND_net), .O(n18686));   // verilog/coms.v(127[12] 300[6])
    defparam i13897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14311_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19100));   // verilog/coms.v(127[12] 300[6])
    defparam i14311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14312_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19101));   // verilog/coms.v(127[12] 300[6])
    defparam i14312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14313_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19102));   // verilog/coms.v(127[12] 300[6])
    defparam i14313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5018));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14314_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19103));   // verilog/coms.v(127[12] 300[6])
    defparam i14314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5017));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5016));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14315_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19104));   // verilog/coms.v(127[12] 300[6])
    defparam i14315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14316_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19105));   // verilog/coms.v(127[12] 300[6])
    defparam i14316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14317_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19106));   // verilog/coms.v(127[12] 300[6])
    defparam i14317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14318_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19107));   // verilog/coms.v(127[12] 300[6])
    defparam i14318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14319_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19108));   // verilog/coms.v(127[12] 300[6])
    defparam i14319_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1322_3_lut (.I0(n1934), .I1(n1987), 
            .I2(n1948), .I3(GND_net), .O(n2012));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14320_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19109));   // verilog/coms.v(127[12] 300[6])
    defparam i14320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14321_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19110));   // verilog/coms.v(127[12] 300[6])
    defparam i14321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1315_3_lut (.I0(n1927), .I1(n1980), 
            .I2(n1948), .I3(GND_net), .O(n2005));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1327_3_lut (.I0(n1939), .I1(n1992), 
            .I2(n1948), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14322_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19111));   // verilog/coms.v(127[12] 300[6])
    defparam i14322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1324_3_lut (.I0(n1936), .I1(n1989), 
            .I2(n1948), .I3(GND_net), .O(n2014));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1325_3_lut (.I0(n1937), .I1(n1990), 
            .I2(n1948), .I3(GND_net), .O(n2015));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1313_3_lut (.I0(n1925), .I1(n1978), 
            .I2(n1948), .I3(GND_net), .O(n2003));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1332_3_lut (.I0(n774), .I1(n1997), 
            .I2(n1948), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1331_3_lut (.I0(n1943), .I1(n1996), 
            .I2(n1948), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4895), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n775));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1317_3_lut (.I0(n1929), .I1(n1982), 
            .I2(n1948), .I3(GND_net), .O(n2007));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1323_3_lut (.I0(n1935), .I1(n1988), 
            .I2(n1948), .I3(GND_net), .O(n2013));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14323_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19112));   // verilog/coms.v(127[12] 300[6])
    defparam i14323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14324_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19113));   // verilog/coms.v(127[12] 300[6])
    defparam i14324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14325_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19114));   // verilog/coms.v(127[12] 300[6])
    defparam i14325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14326_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19115));   // verilog/coms.v(127[12] 300[6])
    defparam i14326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14327_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19116));   // verilog/coms.v(127[12] 300[6])
    defparam i14327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14328_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19117));   // verilog/coms.v(127[12] 300[6])
    defparam i14328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14329_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19118));   // verilog/coms.v(127[12] 300[6])
    defparam i14329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14330_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n2134), .I3(GND_net), .O(n19119));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14331_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n2134), .I3(GND_net), .O(n19120));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1314_3_lut (.I0(n1926), .I1(n1979), 
            .I2(n1948), .I3(GND_net), .O(n2004));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1319_3_lut (.I0(n1931), .I1(n1984), 
            .I2(n1948), .I3(GND_net), .O(n2009));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1316_3_lut (.I0(n1928), .I1(n1981), 
            .I2(n1948), .I3(GND_net), .O(n2006));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1320_3_lut (.I0(n1932), .I1(n1985), 
            .I2(n1948), .I3(GND_net), .O(n2010));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14332_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n2134), .I3(GND_net), .O(n19121));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1326_3_lut (.I0(n1938), .I1(n1991), 
            .I2(n1948), .I3(GND_net), .O(n2016));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1326_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14333_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n2134), .I3(GND_net), .O(n19122));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1310_3_lut (.I0(n1922), .I1(n1975), 
            .I2(n1948), .I3(GND_net), .O(n2000));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1330_3_lut (.I0(n1942), .I1(n1995), 
            .I2(n1948), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1328_3_lut (.I0(n1940), .I1(n1993), 
            .I2(n1948), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14334_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n2134), .I3(GND_net), .O(n19123));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14335_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n2134), .I3(GND_net), .O(n19124));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14336_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n2134), .I3(GND_net), .O(n19125));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1329_3_lut (.I0(n1941), .I1(n1994), 
            .I2(n1948), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1311_3_lut (.I0(n1923), .I1(n1976), 
            .I2(n1948), .I3(GND_net), .O(n2001));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1318_3_lut (.I0(n1930), .I1(n1983), 
            .I2(n1948), .I3(GND_net), .O(n2008));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14337_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n2134), .I3(GND_net), .O(n19126));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1321_3_lut (.I0(n1933), .I1(n1986), 
            .I2(n1948), .I3(GND_net), .O(n2011));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1312_3_lut (.I0(n1924), .I1(n1977), 
            .I2(n1948), .I3(GND_net), .O(n2002));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14338_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n2134), .I3(GND_net), .O(n19127));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut (.I0(n2002), .I1(n2011), .I2(n2008), .I3(n2001), 
            .O(n30_adj_4879));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14339_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n2134), .I3(GND_net), .O(n19128));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19788_3_lut (.I0(n775), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n24570));
    defparam i19788_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut (.I0(n2019), .I1(n2018), .I2(n24570), .I3(n2020), 
            .O(n33723));
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i14340_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n2134), .I3(GND_net), .O(n19129));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15_4_lut (.I0(n2003), .I1(n30_adj_4879), .I2(n2015), .I3(n2014), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2000), .I1(n2016), .I2(n2010), .I3(n2006), 
            .O(n32));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14341_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n2134), .I3(GND_net), .O(n19130));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14342_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n2134), .I3(GND_net), .O(n19131));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14343_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n2134), .I3(GND_net), .O(n19132));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14_4_lut (.I0(n2009), .I1(n2004), .I2(n2013), .I3(n2007), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2017), .I1(n2005), .I2(n2012), .I3(n33723), 
            .O(n31));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14344_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n2134), .I3(GND_net), .O(n19133));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30843_4_lut (.I0(n31), .I1(n33), .I2(n32), .I3(n34), .O(n2026));
    defparam i30843_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14345_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n2134), .I3(GND_net), .O(n19134));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1494_3_lut (.I0(n2026), .I1(n5825), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1494_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1274_3_lut (.I0(n1861), .I1(n1914), 
            .I2(n1870), .I3(GND_net), .O(n1939));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14346_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n2134), .I3(GND_net), .O(n19135));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1269_3_lut (.I0(n1856), .I1(n1909), 
            .I2(n1870), .I3(GND_net), .O(n1934));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1275_3_lut (.I0(n1862), .I1(n1915), 
            .I2(n1870), .I3(GND_net), .O(n1940));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14347_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n2134), .I3(GND_net), .O(n19136));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14348_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n2134), .I3(GND_net), .O(n19137));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1278_3_lut (.I0(n773), .I1(n1918), 
            .I2(n1870), .I3(GND_net), .O(n1943));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1277_3_lut (.I0(n1864), .I1(n1917), 
            .I2(n1870), .I3(GND_net), .O(n1942));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1276_3_lut (.I0(n1863), .I1(n1916), 
            .I2(n1870), .I3(GND_net), .O(n1941));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14349_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n2134), .I3(GND_net), .O(n19138));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3291_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4896), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n774));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14350_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n2134), .I3(GND_net), .O(n19139));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14351_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n2134), .I3(GND_net), .O(n19140));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1259_3_lut (.I0(n1846), .I1(n1899), 
            .I2(n1870), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1264_3_lut (.I0(n1851), .I1(n1904), 
            .I2(n1870), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14352_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n2134), .I3(GND_net), .O(n19141));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1268_3_lut (.I0(n1855), .I1(n1908), 
            .I2(n1870), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14353_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n2134), .I3(GND_net), .O(n19142));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14354_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n2134), .I3(GND_net), .O(n19143));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1261_3_lut (.I0(n1848), .I1(n1901), 
            .I2(n1870), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14355_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n2134), .I3(GND_net), .O(n19144));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14356_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n2134), .I3(GND_net), .O(n19145));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1258_3_lut (.I0(n1845), .I1(n1898), 
            .I2(n1870), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1262_3_lut (.I0(n1849), .I1(n1902), 
            .I2(n1870), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14357_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n2134), .I3(GND_net), .O(n19146));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1271_3_lut (.I0(n1858), .I1(n1911), 
            .I2(n1870), .I3(GND_net), .O(n1936));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14358_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n2134), .I3(GND_net), .O(n19147));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14359_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n2134), .I3(GND_net), .O(n19148));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14360_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n2134), .I3(GND_net), .O(n19149));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1257_3_lut (.I0(n1844), .I1(n1897), 
            .I2(n1870), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13907_3_lut (.I0(n33251), .I1(r_Bit_Index[0]), .I2(n33211), 
            .I3(GND_net), .O(n18696));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13907_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 encoder0_position_23__I_0_i1265_3_lut (.I0(n1852), .I1(n1905), 
            .I2(n1870), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1266_3_lut (.I0(n1853), .I1(n1906), 
            .I2(n1870), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14362_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n34304), .I3(GND_net), .O(n19151));   // verilog/coms.v(127[12] 300[6])
    defparam i14362_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1270_3_lut (.I0(n1857), .I1(n1910), 
            .I2(n1870), .I3(GND_net), .O(n1935));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1263_3_lut (.I0(n1850), .I1(n1903), 
            .I2(n1870), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1267_3_lut (.I0(n1854), .I1(n1907), 
            .I2(n1870), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14363_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n34304), .I3(GND_net), .O(n19152));   // verilog/coms.v(127[12] 300[6])
    defparam i14363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1272_3_lut (.I0(n1859), .I1(n1912), 
            .I2(n1870), .I3(GND_net), .O(n1937));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1273_3_lut (.I0(n1860), .I1(n1913), 
            .I2(n1870), .I3(GND_net), .O(n1938));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1260_3_lut (.I0(n1847), .I1(n1900), 
            .I2(n1870), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_4_lut (.I0(n1925), .I1(n1938), .I2(n1937), .I3(n1932), 
            .O(n28_adj_5035));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1643 (.I0(n1926), .I1(n1933), .I2(n1929), .I3(n1924), 
            .O(n31_adj_5033));
    defparam i13_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i14364_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n34304), .I3(GND_net), .O(n19153));   // verilog/coms.v(127[12] 300[6])
    defparam i14364_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n18163), 
            .D(n617), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n18163), 
            .D(n616), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n18163), 
            .D(n615), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n18163), 
            .D(n614), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n18163), 
            .D(n613), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n18163), 
            .D(n612), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i19906_4_lut (.I0(n774), .I1(n1941), .I2(n1942), .I3(n1943), 
            .O(n24688));
    defparam i19906_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_2_lut (.I0(n1928), .I1(n1935), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_5036));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESR delay_counter_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n18163), 
            .D(n611), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i14365_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n34304), .I3(GND_net), .O(n19154));   // verilog/coms.v(127[12] 300[6])
    defparam i14365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1644 (.I0(n1931), .I1(n1930), .I2(n1922), .I3(n1936), 
            .O(n30_adj_5034));
    defparam i12_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n31_adj_5033), .I1(n1927), .I2(n28_adj_5035), 
            .I3(n1923), .O(n34_adj_5032));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut (.I0(n1940), .I1(n1934), .I2(n1939), .I3(n24688), 
            .O(n21_adj_5037));
    defparam i3_4_lut.LUT_INIT = 16'heccc;
    SB_DFFESR delay_counter_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n18163), 
            .D(n610), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i6_4_lut_adj_1645 (.I0(n32831), .I1(n30832), .I2(n32658), 
            .I3(\data_out_frame[23] [0]), .O(n14_adj_5038));
    defparam i6_4_lut_adj_1645.LUT_INIT = 16'h6996;
    SB_LUT4 i14366_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n34304), .I3(GND_net), .O(n19155));   // verilog/coms.v(127[12] 300[6])
    defparam i14366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n32920), .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[24] [7]), 
            .I3(n32722), .O(n9_adj_5039));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_DFFESR delay_counter_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n18163), 
            .D(n609), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n18163), 
            .D(n608), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n18163), 
            .D(n607), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n18163), 
            .D(n606), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i7_4_lut_adj_1646 (.I0(n9_adj_5039), .I1(n14_adj_5038), .I2(n32699), 
            .I3(n30803), .O(n29929));
    defparam i7_4_lut_adj_1646.LUT_INIT = 16'h6996;
    SB_LUT4 i14367_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n34304), .I3(GND_net), .O(n19156));   // verilog/coms.v(127[12] 300[6])
    defparam i14367_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n18163), 
            .D(n605), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n18163), 
            .D(n604), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i30818_4_lut (.I0(n21_adj_5037), .I1(n34_adj_5032), .I2(n30_adj_5034), 
            .I3(n22_adj_5036), .O(n1948));
    defparam i30818_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1493_3_lut (.I0(n1948), .I1(n5824), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1493_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1217_3_lut (.I0(n1779), .I1(n1832), 
            .I2(n1792), .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1215_3_lut (.I0(n1777), .I1(n1830), 
            .I2(n1792), .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1218_3_lut (.I0(n1780), .I1(n1833), 
            .I2(n1792), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1218_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n18163), 
            .D(n603), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder0_position_23__I_0_i1214_3_lut (.I0(n1776), .I1(n1829), 
            .I2(n1792), .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1214_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n18163), 
            .D(n602), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i14368_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n34304), .I3(GND_net), .O(n19157));   // verilog/coms.v(127[12] 300[6])
    defparam i14368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1207_3_lut (.I0(n1769), .I1(n1822), 
            .I2(n1792), .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1207_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n18163), 
            .D(n601), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder0_position_23__I_0_i1219_3_lut (.I0(n1781), .I1(n1834), 
            .I2(n1792), .I3(GND_net), .O(n1859));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_6_lut (.I0(GND_net), .I1(n755), 
            .I2(GND_net), .I3(n28034), .O(n808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n18163), 
            .D(n600), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n18163), 
            .D(n599), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n18163), 
            .D(n598), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n18163), 
            .D(n597), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder0_position_23__I_0_i1204_3_lut (.I0(n1766), .I1(n1819), 
            .I2(n1792), .I3(GND_net), .O(n1844));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14369_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n34304), .I3(GND_net), .O(n19158));   // verilog/coms.v(127[12] 300[6])
    defparam i14369_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n18163), 
            .D(n596), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFFESR delay_counter_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n18163), 
            .D(n595), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i14370_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n34304), .I3(GND_net), .O(n19159));   // verilog/coms.v(127[12] 300[6])
    defparam i14370_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1224_3_lut (.I0(n772), .I1(n1839), 
            .I2(n1792), .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1224_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1223_3_lut (.I0(n1785), .I1(n1838), 
            .I2(n1792), .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14371_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n34304), .I3(GND_net), .O(n19160));   // verilog/coms.v(127[12] 300[6])
    defparam i14371_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14372_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n34304), .I3(GND_net), .O(n19161));   // verilog/coms.v(127[12] 300[6])
    defparam i14372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4897), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n773));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_513_6 (.CI(n28034), .I0(n755), 
            .I1(GND_net), .CO(n28035));
    SB_LUT4 encoder0_position_23__I_0_i1213_3_lut (.I0(n1775), .I1(n1828), 
            .I2(n1792), .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14373_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n34304), .I3(GND_net), .O(n19162));   // verilog/coms.v(127[12] 300[6])
    defparam i14373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1206_3_lut (.I0(n1768), .I1(n1821), 
            .I2(n1792), .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1209_3_lut (.I0(n1771), .I1(n1824), 
            .I2(n1792), .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1216_3_lut (.I0(n1778), .I1(n1831), 
            .I2(n1792), .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1210_3_lut (.I0(n1772), .I1(n1825), 
            .I2(n1792), .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1205_3_lut (.I0(n1767), .I1(n1820), 
            .I2(n1792), .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14374_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n34304), .I3(GND_net), .O(n19163));   // verilog/coms.v(127[12] 300[6])
    defparam i14374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1212_3_lut (.I0(n1774), .I1(n1827), 
            .I2(n1792), .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1222_3_lut (.I0(n1784), .I1(n1837), 
            .I2(n1792), .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1220_3_lut (.I0(n1782), .I1(n1835), 
            .I2(n1792), .I3(GND_net), .O(n1860));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1221_3_lut (.I0(n1783), .I1(n1836), 
            .I2(n1792), .I3(GND_net), .O(n1861));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5015));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1208_3_lut (.I0(n1770), .I1(n1823), 
            .I2(n1792), .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1211_3_lut (.I0(n1773), .I1(n1826), 
            .I2(n1792), .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14375_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n34304), .I3(GND_net), .O(n19164));   // verilog/coms.v(127[12] 300[6])
    defparam i14375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut (.I0(n1851), .I1(n1848), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5028));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19814_3_lut (.I0(n773), .I1(n1863), .I2(n1864), .I3(GND_net), 
            .O(n24596));
    defparam i19814_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1647 (.I0(n1861), .I1(n1860), .I2(n24596), .I3(n1862), 
            .O(n33837));
    defparam i2_4_lut_adj_1647.LUT_INIT = 16'h8880;
    SB_LUT4 i14376_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n34304), .I3(GND_net), .O(n19165));   // verilog/coms.v(127[12] 300[6])
    defparam i14376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_4_lut_adj_1648 (.I0(n1844), .I1(n1859), .I2(n1847), .I3(n18_adj_5028), 
            .O(n30_adj_5024));
    defparam i13_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1649 (.I0(n1852), .I1(n33837), .I2(n1845), .I3(n1850), 
            .O(n28_adj_5026));
    defparam i11_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1650 (.I0(n1856), .I1(n1849), .I2(n1846), .I3(n1853), 
            .O(n29_adj_5025));
    defparam i12_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1651 (.I0(n1854), .I1(n1858), .I2(n1855), .I3(n1857), 
            .O(n27_adj_5027));
    defparam i10_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i30791_4_lut (.I0(n27_adj_5027), .I1(n29_adj_5025), .I2(n28_adj_5026), 
            .I3(n30_adj_5024), .O(n1870));
    defparam i30791_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14377_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n34304), .I3(GND_net), .O(n19166));   // verilog/coms.v(127[12] 300[6])
    defparam i14377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14378_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n34304), .I3(GND_net), .O(n19167));   // verilog/coms.v(127[12] 300[6])
    defparam i14378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1492_3_lut (.I0(n1870), .I1(n5823), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1492_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i14379_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n34304), .I3(GND_net), .O(n19168));   // verilog/coms.v(127[12] 300[6])
    defparam i14379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1165_3_lut (.I0(n1702), .I1(n1755), 
            .I2(n1714), .I3(GND_net), .O(n1780));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1165_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1154_3_lut (.I0(n1691), .I1(n1744), 
            .I2(n1714), .I3(GND_net), .O(n1769));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14380_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n34304), .I3(GND_net), .O(n19169));   // verilog/coms.v(127[12] 300[6])
    defparam i14380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_5_lut (.I0(GND_net), .I1(n756), 
            .I2(VCC_net), .I3(n28033), .O(n809)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14381_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n34304), .I3(GND_net), .O(n19170));   // verilog/coms.v(127[12] 300[6])
    defparam i14381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1161_3_lut (.I0(n1698), .I1(n1751), 
            .I2(n1714), .I3(GND_net), .O(n1776));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1153_3_lut (.I0(n1690), .I1(n1743), 
            .I2(n1714), .I3(GND_net), .O(n1768));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1159_3_lut (.I0(n1696), .I1(n1749), 
            .I2(n1714), .I3(GND_net), .O(n1774));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14382_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n34304), .I3(GND_net), .O(n19171));   // verilog/coms.v(127[12] 300[6])
    defparam i14382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1162_3_lut (.I0(n1699), .I1(n1752), 
            .I2(n1714), .I3(GND_net), .O(n1777));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1162_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_513_5 (.CI(n28033), .I0(n756), 
            .I1(VCC_net), .CO(n28034));
    SB_LUT4 encoder0_position_23__I_0_i1163_3_lut (.I0(n1700), .I1(n1753), 
            .I2(n1714), .I3(GND_net), .O(n1778));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1163_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1170_3_lut (.I0(n771), .I1(n1760), 
            .I2(n1714), .I3(GND_net), .O(n1785));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1169_3_lut (.I0(n1706), .I1(n1759), 
            .I2(n1714), .I3(GND_net), .O(n1784));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4898), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n772));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1156_3_lut (.I0(n1693), .I1(n1746), 
            .I2(n1714), .I3(GND_net), .O(n1771));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14383_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n34304), .I3(GND_net), .O(n19172));   // verilog/coms.v(127[12] 300[6])
    defparam i14383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1151_3_lut (.I0(n1688), .I1(n1741), 
            .I2(n1714), .I3(GND_net), .O(n1766));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1158_3_lut (.I0(n1695), .I1(n1748), 
            .I2(n1714), .I3(GND_net), .O(n1773));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1155_3_lut (.I0(n1692), .I1(n1745), 
            .I2(n1714), .I3(GND_net), .O(n1770));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1164_3_lut (.I0(n1701), .I1(n1754), 
            .I2(n1714), .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14384_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n34304), .I3(GND_net), .O(n19173));   // verilog/coms.v(127[12] 300[6])
    defparam i14384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1160_3_lut (.I0(n1697), .I1(n1750), 
            .I2(n1714), .I3(GND_net), .O(n1775));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1160_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1152_3_lut (.I0(n1689), .I1(n1742), 
            .I2(n1714), .I3(GND_net), .O(n1767));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1157_3_lut (.I0(n1694), .I1(n1747), 
            .I2(n1714), .I3(GND_net), .O(n1772));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14385_4_lut (.I0(state_7__N_3877[3]), .I1(data[1]), .I2(n10_adj_4966), 
            .I3(n17058), .O(n19174));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i14385_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14386_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n34934), 
            .I3(GND_net), .O(n19175));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1168_3_lut (.I0(n1705), .I1(n1758), 
            .I2(n1714), .I3(GND_net), .O(n1783));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1166_3_lut (.I0(n1703), .I1(n1756), 
            .I2(n1714), .I3(GND_net), .O(n1781));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1167_3_lut (.I0(n1704), .I1(n1757), 
            .I2(n1714), .I3(GND_net), .O(n1782));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19816_3_lut (.I0(n772), .I1(n1784), .I2(n1785), .I3(GND_net), 
            .O(n24598));
    defparam i19816_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i29790_4_lut (.I0(n33407), .I1(n5_adj_4919), .I2(n6_adj_4918), 
            .I3(state[0]), .O(n35881));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29790_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i2_4_lut_adj_1652 (.I0(n1782), .I1(n1781), .I2(n24598), .I3(n1783), 
            .O(n33450));
    defparam i2_4_lut_adj_1652.LUT_INIT = 16'h8880;
    SB_LUT4 i18_4_lut (.I0(n35881), .I1(n35879), .I2(state[1]), .I3(n4_adj_4961), 
            .O(n31374));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i12_4_lut_adj_1653 (.I0(n1772), .I1(n1767), .I2(n1775), .I3(n1779), 
            .O(n28_adj_5044));
    defparam i12_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i14396_3_lut (.I0(quadA_debounced_adj_4922), .I1(reg_B_adj_5120[1]), 
            .I2(n34883), .I3(GND_net), .O(n19185));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13871_3_lut (.I0(n18590), .I1(r_Bit_Index_adj_5113[0]), .I2(n18336), 
            .I3(GND_net), .O(n18660));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13871_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i10_4_lut_adj_1654 (.I0(n1770), .I1(n1773), .I2(n1766), .I3(n1771), 
            .O(n26_adj_5046));
    defparam i10_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1655 (.I0(n1778), .I1(n1777), .I2(n1774), .I3(n1768), 
            .O(n27_adj_5045));
    defparam i11_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n33450), .I1(n1776), .I2(n1769), .I3(n1780), 
            .O(n25_adj_5047));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30765_4_lut (.I0(n25_adj_5047), .I1(n27_adj_5045), .I2(n26_adj_5046), 
            .I3(n28_adj_5044), .O(n1792));
    defparam i30765_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1491_3_lut (.I0(n1792), .I1(n5822), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1491_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1109_3_lut (.I0(n1621), .I1(n1674), 
            .I2(n1636), .I3(GND_net), .O(n1699));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1099_3_lut (.I0(n1611), .I1(n1664), 
            .I2(n1636), .I3(GND_net), .O(n1689));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1099_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1101_3_lut (.I0(n1613), .I1(n1666), 
            .I2(n1636), .I3(GND_net), .O(n1691));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1104_3_lut (.I0(n1616), .I1(n1669), 
            .I2(n1636), .I3(GND_net), .O(n1694));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1107_3_lut (.I0(n1619), .I1(n1672), 
            .I2(n1636), .I3(GND_net), .O(n1697));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14399_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n33905), .I3(GND_net), 
            .O(n19188));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i14399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1112_3_lut (.I0(n1624), .I1(n1677), 
            .I2(n1636), .I3(GND_net), .O(n1702));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14400_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n33905), .I3(GND_net), 
            .O(n19189));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i14400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14401_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n33905), .I3(GND_net), 
            .O(n19190));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i14401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5014));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1113_3_lut (.I0(n1625), .I1(n1678), 
            .I2(n1636), .I3(GND_net), .O(n1703));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1110_3_lut (.I0(n1622), .I1(n1675), 
            .I2(n1636), .I3(GND_net), .O(n1700));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1116_3_lut (.I0(n770), .I1(n1681), 
            .I2(n1636), .I3(GND_net), .O(n1706));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1115_3_lut (.I0(n1627), .I1(n1680), 
            .I2(n1636), .I3(GND_net), .O(n1705));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5013));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5012));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1114_3_lut (.I0(n1626), .I1(n1679), 
            .I2(n1636), .I3(GND_net), .O(n1704));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4899), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n771));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1106_3_lut (.I0(n1618), .I1(n1671), 
            .I2(n1636), .I3(GND_net), .O(n1696));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14402_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n33905), .I3(GND_net), 
            .O(n19191));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i14402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1100_3_lut (.I0(n1612), .I1(n1665), 
            .I2(n1636), .I3(GND_net), .O(n1690));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1103_3_lut (.I0(n1615), .I1(n1668), 
            .I2(n1636), .I3(GND_net), .O(n1693));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1108_3_lut (.I0(n1620), .I1(n1673), 
            .I2(n1636), .I3(GND_net), .O(n1698));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14403_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n33905), .I3(GND_net), 
            .O(n19192));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i14403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1111_3_lut (.I0(n1623), .I1(n1676), 
            .I2(n1636), .I3(GND_net), .O(n1701));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14404_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n33905), .I3(GND_net), 
            .O(n19193));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i14404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1102_3_lut (.I0(n1614), .I1(n1667), 
            .I2(n1636), .I3(GND_net), .O(n1692));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1105_3_lut (.I0(n1617), .I1(n1670), 
            .I2(n1636), .I3(GND_net), .O(n1695));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1098_3_lut (.I0(n1610), .I1(n1663), 
            .I2(n1636), .I3(GND_net), .O(n1688));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19920_4_lut (.I0(n771), .I1(n1704), .I2(n1705), .I3(n1706), 
            .O(n24702));
    defparam i19920_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i14405_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n33905), .I3(GND_net), 
            .O(n19194));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i14405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i11_4_lut_adj_1656 (.I0(n1688), .I1(n1695), .I2(n1692), .I3(n1701), 
            .O(n26_adj_5057));
    defparam i11_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(n1700), .I1(n1703), .I2(n1702), .I3(n24702), 
            .O(n19_adj_5059));
    defparam i4_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i259_2_lut (.I0(n619), .I1(n15_adj_4867), .I2(GND_net), .I3(GND_net), 
            .O(n1172));   // verilog/TinyFPGA_B.v(252[9] 258[12])
    defparam i259_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1657 (.I0(n1698), .I1(n1693), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_5060));
    defparam i1_2_lut_adj_1657.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1658 (.I0(n1697), .I1(n1694), .I2(n1691), .I3(n1689), 
            .O(n24_adj_5058));
    defparam i9_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1659 (.I0(n19_adj_5059), .I1(n26_adj_5057), .I2(n1690), 
            .I3(n1696), .O(n28_adj_5056));
    defparam i13_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i30740_4_lut (.I0(n1699), .I1(n28_adj_5056), .I2(n24_adj_5058), 
            .I3(n16_adj_5060), .O(n1714));
    defparam i30740_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1490_3_lut (.I0(n1714), .I1(n5821), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1490_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1054_3_lut (.I0(n1541), .I1(n1594), 
            .I2(n1558), .I3(GND_net), .O(n1619));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1660 (.I0(n23704), .I1(n32413), .I2(state_adj_5104[0]), 
            .I3(read), .O(n32064));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1660.LUT_INIT = 16'h8280;
    SB_LUT4 encoder0_position_23__I_0_i1056_3_lut (.I0(n1543), .I1(n1596), 
            .I2(n1558), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1055_3_lut (.I0(n1542), .I1(n1595), 
            .I2(n1558), .I3(GND_net), .O(n1620));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1057_3_lut (.I0(n1544), .I1(n1597), 
            .I2(n1558), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1045_3_lut (.I0(n1532), .I1(n1585), 
            .I2(n1558), .I3(GND_net), .O(n1610));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14408_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n23776), 
            .I3(n17084), .O(n19197));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14408_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_23__I_0_i1053_3_lut (.I0(n1540), .I1(n1593), 
            .I2(n1558), .I3(GND_net), .O(n1618));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1046_3_lut (.I0(n1533), .I1(n1586), 
            .I2(n1558), .I3(GND_net), .O(n1611));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1062_3_lut (.I0(n769), .I1(n1602), 
            .I2(n1558), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5011));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5010));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1061_3_lut (.I0(n1548), .I1(n1601), 
            .I2(n1558), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14409_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n23776), 
            .I3(n17079), .O(n19198));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14409_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 mux_3291_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4900), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n770));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1048_3_lut (.I0(n1535), .I1(n1588), 
            .I2(n1558), .I3(GND_net), .O(n1613));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1051_3_lut (.I0(n1538), .I1(n1591), 
            .I2(n1558), .I3(GND_net), .O(n1616));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1050_3_lut (.I0(n1537), .I1(n1590), 
            .I2(n1558), .I3(GND_net), .O(n1615));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5009));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1052_3_lut (.I0(n1539), .I1(n1592), 
            .I2(n1558), .I3(GND_net), .O(n1617));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1047_3_lut (.I0(n1534), .I1(n1587), 
            .I2(n1558), .I3(GND_net), .O(n1612));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5008));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14410_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4921), 
            .I3(n17084), .O(n19199));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14410_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i1049_3_lut (.I0(n1536), .I1(n1589), 
            .I2(n1558), .I3(GND_net), .O(n1614));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1060_3_lut (.I0(n1547), .I1(n1600), 
            .I2(n1558), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1058_3_lut (.I0(n1545), .I1(n1598), 
            .I2(n1558), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1059_3_lut (.I0(n1546), .I1(n1599), 
            .I2(n1558), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19824_3_lut (.I0(n770), .I1(n1626), .I2(n1627), .I3(GND_net), 
            .O(n24606));
    defparam i19824_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1661 (.I0(n1624), .I1(n1623), .I2(n24606), .I3(n1625), 
            .O(n34140));
    defparam i2_4_lut_adj_1661.LUT_INIT = 16'h8880;
    SB_LUT4 i4_2_lut_adj_1662 (.I0(n1611), .I1(n1618), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5065));
    defparam i4_2_lut_adj_1662.LUT_INIT = 16'heeee;
    SB_LUT4 i14411_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4921), 
            .I3(n17079), .O(n19200));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14411_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i10_4_lut_adj_1663 (.I0(n1614), .I1(n1612), .I2(n1617), .I3(n1615), 
            .O(n24_adj_5063));
    defparam i10_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i14412_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4), .I3(n17084), 
            .O(n19201));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14412_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8_4_lut (.I0(n1610), .I1(n1622), .I2(n1620), .I3(n34140), 
            .O(n22_adj_5064));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14413_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4), .I3(n17079), 
            .O(n19202));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14413_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12_4_lut_adj_1664 (.I0(n1616), .I1(n24_adj_5063), .I2(n18_adj_5065), 
            .I3(n1613), .O(n26_adj_5062));
    defparam i12_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i30716_4_lut (.I0(n1621), .I1(n26_adj_5062), .I2(n22_adj_5064), 
            .I3(n1619), .O(n1636));
    defparam i30716_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5007));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5006));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5005));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5004));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5003));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30848_1_lut (.I0(n700), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37245));
    defparam i30848_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5002));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5001));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1489_3_lut (.I0(n1636), .I1(n5820), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1489_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1001_3_lut (.I0(n1463), .I1(n1516), 
            .I2(n1480), .I3(GND_net), .O(n1541));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i995_3_lut (.I0(n1457), .I1(n1510), 
            .I2(n1480), .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5000));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1003_3_lut (.I0(n1465), .I1(n1518), 
            .I2(n1480), .I3(GND_net), .O(n1543));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i996_3_lut (.I0(n1458), .I1(n1511), 
            .I2(n1480), .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i999_3_lut (.I0(n1461), .I1(n1514), 
            .I2(n1480), .I3(GND_net), .O(n1539));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1000_3_lut (.I0(n1462), .I1(n1515), 
            .I2(n1480), .I3(GND_net), .O(n1540));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26776_4_lut (.I0(n7_adj_5043), .I1(state_adj_5104[0]), .I2(n6_adj_5055), 
            .I3(state_adj_5132[0]), .O(n33160));
    defparam i26776_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 encoder0_position_23__I_0_i998_3_lut (.I0(n1460), .I1(n1513), 
            .I2(n1480), .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1002_3_lut (.I0(n1464), .I1(n1517), 
            .I2(n1480), .I3(GND_net), .O(n1542));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i993_3_lut (.I0(n1455), .I1(n1508), 
            .I2(n1480), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1008_3_lut (.I0(n768), .I1(n1523), 
            .I2(n1480), .I3(GND_net), .O(n1548));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1007_3_lut (.I0(n1469), .I1(n1522), 
            .I2(n1480), .I3(GND_net), .O(n1547));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1006_3_lut (.I0(n1468), .I1(n1521), 
            .I2(n1480), .I3(GND_net), .O(n1546));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1006_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_4901), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n769));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i992_3_lut (.I0(n1454), .I1(n1507), 
            .I2(n1480), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut (.I0(state_adj_5104[1]), .I1(read), .I2(n32413), 
            .I3(GND_net), .O(n12_adj_5029));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 encoder0_position_23__I_0_i997_3_lut (.I0(n1459), .I1(n1512), 
            .I2(n1480), .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4999));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1004_3_lut (.I0(n1466), .I1(n1519), 
            .I2(n1480), .I3(GND_net), .O(n1544));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4998));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1665 (.I0(n23704), .I1(n12_adj_5029), .I2(state_adj_5104[0]), 
            .I3(n32413), .O(n32068));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1665.LUT_INIT = 16'h88a8;
    SB_LUT4 encoder0_position_23__I_0_i994_3_lut (.I0(n1456), .I1(n1509), 
            .I2(n1480), .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1005_3_lut (.I0(n1467), .I1(n1520), 
            .I2(n1480), .I3(GND_net), .O(n1545));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19927_4_lut (.I0(n769), .I1(n1546), .I2(n1547), .I3(n1548), 
            .O(n24710));
    defparam i19927_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4997));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4996));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4995));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_4_lut_adj_1666 (.I0(n1545), .I1(n1534), .I2(n1544), .I3(n24710), 
            .O(n17_adj_4994));
    defparam i4_4_lut_adj_1666.LUT_INIT = 16'heccc;
    SB_LUT4 i8_4_lut_adj_1667 (.I0(n1533), .I1(n1542), .I2(n1538), .I3(n1540), 
            .O(n21_adj_4992));
    defparam i8_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i14415_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4893), 
            .I3(n17084), .O(n19204));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14415_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i7_3_lut (.I0(n1539), .I1(n1536), .I2(n1543), .I3(GND_net), 
            .O(n20_adj_4993));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1668 (.I0(n21_adj_4992), .I1(n17_adj_4994), .I2(n1537), 
            .I3(n1532), .O(n24_adj_4991));
    defparam i11_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i13852_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n34934), 
            .I3(GND_net), .O(n18641));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1669 (.I0(enable_slow_N_3964), .I1(data_ready), 
            .I2(state_adj_5104[1]), .I3(state_adj_5104[0]), .O(n32166));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1669.LUT_INIT = 16'hccd0;
    SB_LUT4 mux_72_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[0]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i30693_4_lut (.I0(n1535), .I1(n24_adj_4991), .I2(n20_adj_4993), 
            .I3(n1541), .O(n1558));
    defparam i30693_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_70_i1_3_lut (.I0(encoder0_position_scaled[0]), .I1(motor_state_23__N_82[0]), 
            .I2(n15), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13854_4_lut (.I0(rw), .I1(state_adj_5104[0]), .I2(state_adj_5104[1]), 
            .I3(n3568), .O(n18643));   // verilog/eeprom.v(26[8] 58[4])
    defparam i13854_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 mux_72_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[1]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i2_3_lut (.I0(encoder0_position_scaled[1]), .I1(motor_state_23__N_82[1]), 
            .I2(n15), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_23__I_0_i1488_3_lut (.I0(n1558), .I1(n5819), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1488_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 mux_72_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[2]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_i940_3_lut (.I0(n1377), .I1(n1430), 
            .I2(n1402), .I3(GND_net), .O(n1455));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i947_3_lut (.I0(n1384), .I1(n1437), 
            .I2(n1402), .I3(GND_net), .O(n1462));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i3_3_lut (.I0(encoder0_position_scaled[2]), .I1(motor_state_23__N_82[2]), 
            .I2(n15), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_23__I_0_i944_3_lut (.I0(n1381), .I1(n1434), 
            .I2(n1402), .I3(GND_net), .O(n1459));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13855_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5111[1]), .I2(n10125), 
            .I3(n4_adj_5053), .O(n18644));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13855_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 encoder0_position_23__I_0_i946_3_lut (.I0(n1383), .I1(n1436), 
            .I2(n1402), .I3(GND_net), .O(n1461));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i950_3_lut (.I0(n1387), .I1(n1440), 
            .I2(n1402), .I3(GND_net), .O(n1465));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i950_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13856_3_lut (.I0(quadB_debounced_adj_4923), .I1(reg_B_adj_5120[0]), 
            .I2(n34883), .I3(GND_net), .O(n18645));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13856_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i951_3_lut (.I0(n1388), .I1(n1441), 
            .I2(n1402), .I3(GND_net), .O(n1466));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i951_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i942_3_lut (.I0(n1379), .I1(n1432), 
            .I2(n1402), .I3(GND_net), .O(n1457));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i954_3_lut (.I0(n767), .I1(n1444), 
            .I2(n1402), .I3(GND_net), .O(n1469));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13857_4_lut (.I0(state_7__N_3877[3]), .I1(data[5]), .I2(n4_adj_4927), 
            .I3(n17058), .O(n18646));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13857_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i953_3_lut (.I0(n1390), .I1(n1443), 
            .I2(n1402), .I3(GND_net), .O(n1468));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i952_3_lut (.I0(n1389), .I1(n1442), 
            .I2(n1402), .I3(GND_net), .O(n1467));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4902), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n768));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i939_3_lut (.I0(n1376), .I1(n1429), 
            .I2(n1402), .I3(GND_net), .O(n1454));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i945_3_lut (.I0(n1382), .I1(n1435), 
            .I2(n1402), .I3(GND_net), .O(n1460));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i941_3_lut (.I0(n1378), .I1(n1431), 
            .I2(n1402), .I3(GND_net), .O(n1456));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i948_3_lut (.I0(n1385), .I1(n1438), 
            .I2(n1402), .I3(GND_net), .O(n1463));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i948_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i943_3_lut (.I0(n1380), .I1(n1433), 
            .I2(n1402), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_72_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[3]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_i949_3_lut (.I0(n1386), .I1(n1439), 
            .I2(n1402), .I3(GND_net), .O(n1464));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i4_3_lut (.I0(encoder0_position_scaled[3]), .I1(motor_state_23__N_82[3]), 
            .I2(n15), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_72_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[4]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i19929_4_lut (.I0(n768), .I1(n1467), .I2(n1468), .I3(n1469), 
            .O(n24712));
    defparam i19929_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i8_4_lut_adj_1670 (.I0(n1464), .I1(n1458), .I2(n1463), .I3(n1456), 
            .O(n20_adj_4888));
    defparam i8_4_lut_adj_1670.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1671 (.I0(n1457), .I1(n1466), .I2(n1465), .I3(n24712), 
            .O(n13_adj_4890));
    defparam i1_4_lut_adj_1671.LUT_INIT = 16'heaaa;
    SB_LUT4 i6_2_lut (.I0(n1461), .I1(n1459), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4889));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_70_i5_3_lut (.I0(encoder0_position_scaled[4]), .I1(motor_state_23__N_82[4]), 
            .I2(n15), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i10_4_lut_adj_1672 (.I0(n13_adj_4890), .I1(n20_adj_4888), .I2(n1460), 
            .I3(n1454), .O(n22_adj_4887));
    defparam i10_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i30609_4_lut (.I0(n1462), .I1(n22_adj_4887), .I2(n18_adj_4889), 
            .I3(n1455), .O(n1480));
    defparam i30609_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1487_3_lut (.I0(n1480), .I1(n5818), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1487_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i892_3_lut (.I0(n1304), .I1(n1357), 
            .I2(n1324), .I3(GND_net), .O(n1382));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i886_3_lut (.I0(n1298), .I1(n1351), 
            .I2(n1324), .I3(GND_net), .O(n1376));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i891_3_lut (.I0(n1303), .I1(n1356), 
            .I2(n1324), .I3(GND_net), .O(n1381));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i895_3_lut (.I0(n1307), .I1(n1360), 
            .I2(n1324), .I3(GND_net), .O(n1385));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i898_3_lut (.I0(n1310), .I1(n1363), 
            .I2(n1324), .I3(GND_net), .O(n1388));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i898_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i896_3_lut (.I0(n1308), .I1(n1361), 
            .I2(n1324), .I3(GND_net), .O(n1386));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i897_3_lut (.I0(n1309), .I1(n1362), 
            .I2(n1324), .I3(GND_net), .O(n1387));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i900_3_lut (.I0(n523), .I1(n1365), 
            .I2(n1324), .I3(GND_net), .O(n1390));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i899_3_lut (.I0(n1311), .I1(n1364), 
            .I2(n1324), .I3(GND_net), .O(n1389));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4903), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n767));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i888_3_lut (.I0(n1300), .I1(n1353), 
            .I2(n1324), .I3(GND_net), .O(n1378));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i894_3_lut (.I0(n1306), .I1(n1359), 
            .I2(n1324), .I3(GND_net), .O(n1384));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i894_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i889_3_lut (.I0(n1301), .I1(n1354), 
            .I2(n1324), .I3(GND_net), .O(n1379));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13858_4_lut (.I0(state_7__N_3877[3]), .I1(data[4]), .I2(n4_adj_4927), 
            .I3(n17053), .O(n18647));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13858_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i887_3_lut (.I0(n1299), .I1(n1352), 
            .I2(n1324), .I3(GND_net), .O(n1377));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i890_3_lut (.I0(n1302), .I1(n1355), 
            .I2(n1324), .I3(GND_net), .O(n1380));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i890_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i893_3_lut (.I0(n1305), .I1(n1358), 
            .I2(n1324), .I3(GND_net), .O(n1383));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19834_3_lut (.I0(n767), .I1(n1389), .I2(n1390), .I3(GND_net), 
            .O(n24616));
    defparam i19834_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1673 (.I0(n1387), .I1(n1386), .I2(n24616), .I3(n1388), 
            .O(n34465));
    defparam i2_4_lut_adj_1673.LUT_INIT = 16'h8880;
    SB_LUT4 i7_4_lut_adj_1674 (.I0(n1383), .I1(n1380), .I2(n1377), .I3(n34465), 
            .O(n18));
    defparam i7_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1385), .I1(n1381), .I2(GND_net), .I3(GND_net), 
            .O(n16));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_add_513_4_lut (.I0(GND_net), .I1(n757), 
            .I2(GND_net), .I3(n28032), .O(n810)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1675 (.I0(n1379), .I1(n18), .I2(n1384), .I3(n1378), 
            .O(n20));
    defparam i9_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 i30545_4_lut (.I0(n1376), .I1(n20), .I2(n16), .I3(n1382), 
            .O(n1402));
    defparam i30545_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1486_3_lut (.I0(n1402), .I1(n5817), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1486_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i834_3_lut (.I0(n1221), .I1(n1274), 
            .I2(n1246), .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i836_3_lut (.I0(n1223), .I1(n1276), 
            .I2(n1246), .I3(GND_net), .O(n1301));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i839_3_lut (.I0(n1226), .I1(n1279), 
            .I2(n1246), .I3(GND_net), .O(n1304));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i841_3_lut (.I0(n1228), .I1(n1281), 
            .I2(n1246), .I3(GND_net), .O(n1306));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i835_3_lut (.I0(n1222), .I1(n1275), 
            .I2(n1246), .I3(GND_net), .O(n1300));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i846_3_lut (.I0(n765), .I1(n1286), 
            .I2(n1246), .I3(GND_net), .O(n1311));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i845_3_lut (.I0(n1232), .I1(n1285), 
            .I2(n1246), .I3(GND_net), .O(n1310));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4904), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i840_3_lut (.I0(n1227), .I1(n1280), 
            .I2(n1246), .I3(GND_net), .O(n1305));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i833_3_lut (.I0(n1220), .I1(n1273), 
            .I2(n1246), .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i833_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i837_3_lut (.I0(n1224), .I1(n1277), 
            .I2(n1246), .I3(GND_net), .O(n1302));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i838_3_lut (.I0(n1225), .I1(n1278), 
            .I2(n1246), .I3(GND_net), .O(n1303));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i844_3_lut (.I0(n1231), .I1(n1284), 
            .I2(n1246), .I3(GND_net), .O(n1309));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13859_4_lut (.I0(state_7__N_3877[3]), .I1(data[3]), .I2(n4_adj_4865), 
            .I3(n17058), .O(n18648));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13859_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i842_3_lut (.I0(n1229), .I1(n1282), 
            .I2(n1246), .I3(GND_net), .O(n1307));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i843_3_lut (.I0(n1230), .I1(n1283), 
            .I2(n1246), .I3(GND_net), .O(n1308));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13860_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_3861[0]), 
            .I3(enable_slow_N_3964), .O(n18649));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13860_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 i19838_3_lut (.I0(n523), .I1(n1310), .I2(n1311), .I3(GND_net), 
            .O(n24620));
    defparam i19838_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1676 (.I0(n1308), .I1(n1307), .I2(n24620), .I3(n1309), 
            .O(n34334));
    defparam i2_4_lut_adj_1676.LUT_INIT = 16'h8880;
    SB_LUT4 i6_4_lut_adj_1677 (.I0(n1300), .I1(n34334), .I2(n1306), .I3(n1304), 
            .O(n16_adj_4882));
    defparam i6_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1678 (.I0(n1303), .I1(n1302), .I2(n1298), .I3(n1305), 
            .O(n17_adj_4881));
    defparam i7_4_lut_adj_1678.LUT_INIT = 16'hfffe;
    SB_LUT4 i13861_4_lut (.I0(state_7__N_3877[3]), .I1(data[2]), .I2(n4_adj_4865), 
            .I3(n17053), .O(n18650));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13861_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30517_4_lut (.I0(n17_adj_4881), .I1(n1301), .I2(n16_adj_4882), 
            .I3(n1299), .O(n1324));
    defparam i30517_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i2_3_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), .I2(\ID_READOUT_FSM.state [1]), 
            .I3(GND_net), .O(n33905));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 encoder0_position_23__I_0_i1485_3_lut (.I0(n1324), .I1(n5816), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1485_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i780_3_lut (.I0(n1142), .I1(n1195), 
            .I2(n1168), .I3(GND_net), .O(n1220));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i786_3_lut (.I0(n1148), .I1(n1201), 
            .I2(n1168), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i788_3_lut (.I0(n1150), .I1(n1203), 
            .I2(n1168), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13862_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n33905), .I3(GND_net), 
            .O(n18651));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i13862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i782_3_lut (.I0(n1144), .I1(n1197), 
            .I2(n1168), .I3(GND_net), .O(n1222));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i789_3_lut (.I0(n1151), .I1(n1204), 
            .I2(n1168), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13863_4_lut (.I0(state_7__N_3877[3]), .I1(data[0]), .I2(n10_adj_4966), 
            .I3(n17053), .O(n18652));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13863_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_i781_3_lut (.I0(n1143), .I1(n1196), 
            .I2(n1168), .I3(GND_net), .O(n1221));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i787_3_lut (.I0(n1149), .I1(n1202), 
            .I2(n1168), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i785_3_lut (.I0(n1147), .I1(n1200), 
            .I2(n1168), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i784_3_lut (.I0(n1146), .I1(n1199), 
            .I2(n1168), .I3(GND_net), .O(n1224));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i783_3_lut (.I0(n1145), .I1(n1198), 
            .I2(n1168), .I3(GND_net), .O(n1223));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i792_3_lut (.I0(n521), .I1(n1207), 
            .I2(n1168), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i791_3_lut (.I0(n1153), .I1(n1206), 
            .I2(n1168), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i790_3_lut (.I0(n1152), .I1(n1205), 
            .I2(n1168), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4905), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n765));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19840_4_lut (.I0(n765), .I1(n1230), .I2(n1231), .I3(n1232), 
            .O(n24622));
    defparam i19840_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1679 (.I0(n1223), .I1(n1224), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4885));
    defparam i1_2_lut_adj_1679.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_1680 (.I0(n1229), .I1(n1222), .I2(n1228), .I3(n24622), 
            .O(n12_adj_4884));
    defparam i3_4_lut_adj_1680.LUT_INIT = 16'heccc;
    SB_LUT4 i7_4_lut_adj_1681 (.I0(n1225), .I1(n1227), .I2(n1221), .I3(n10_adj_4885), 
            .O(n16_adj_4883));
    defparam i7_4_lut_adj_1681.LUT_INIT = 16'hfffe;
    SB_LUT4 i30877_4_lut (.I0(n1226), .I1(n16_adj_4883), .I2(n12_adj_4884), 
            .I3(n1220), .O(n1246));
    defparam i30877_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1484_3_lut (.I0(n1246), .I1(n5815), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1484_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i2_2_lut_adj_1682 (.I0(ID[1]), .I1(ID[2]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4892));   // verilog/TinyFPGA_B.v(252[12:17])
    defparam i2_2_lut_adj_1682.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_i728_3_lut (.I0(n1065), .I1(n1118), 
            .I2(n1090), .I3(GND_net), .O(n1143));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i727_3_lut (.I0(n1064), .I1(n1117), 
            .I2(n1090), .I3(GND_net), .O(n1142));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i738_3_lut (.I0(n763), .I1(n1128), 
            .I2(n1090), .I3(GND_net), .O(n1153));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i737_3_lut (.I0(n1074), .I1(n1127), 
            .I2(n1090), .I3(GND_net), .O(n1152));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i736_3_lut (.I0(n1073), .I1(n1126), 
            .I2(n1090), .I3(GND_net), .O(n1151));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i736_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4906), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i734_3_lut (.I0(n1071), .I1(n1124), 
            .I2(n1090), .I3(GND_net), .O(n1149));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i734_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_513_4 (.CI(n28032), .I0(n757), 
            .I1(GND_net), .CO(n28033));
    SB_LUT4 encoder0_position_23__I_0_i730_3_lut (.I0(n1067), .I1(n1120), 
            .I2(n1090), .I3(GND_net), .O(n1145));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i730_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i735_3_lut (.I0(n1072), .I1(n1125), 
            .I2(n1090), .I3(GND_net), .O(n1150));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i732_3_lut (.I0(n1069), .I1(n1122), 
            .I2(n1090), .I3(GND_net), .O(n1147));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i732_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i729_3_lut (.I0(n1066), .I1(n1119), 
            .I2(n1090), .I3(GND_net), .O(n1144));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i733_3_lut (.I0(n1070), .I1(n1123), 
            .I2(n1090), .I3(GND_net), .O(n1148));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i733_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1683 (.I0(\FRAME_MATCHER.i_31__N_2461 ), .I1(n63), 
            .I2(n3303), .I3(n123), .O(n4_adj_4866));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1683.LUT_INIT = 16'haaa2;
    SB_LUT4 encoder0_position_23__I_0_i731_3_lut (.I0(n1068), .I1(n1121), 
            .I2(n1090), .I3(GND_net), .O(n1146));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19842_4_lut (.I0(n521), .I1(n1151), .I2(n1152), .I3(n1153), 
            .O(n24624));
    defparam i19842_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n123), .I1(n1), .I2(n63), .I3(n32404), 
            .O(n7));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'haf8c;
    SB_LUT4 i6_4_lut_adj_1685 (.I0(n1146), .I1(n1148), .I2(n1144), .I3(n1147), 
            .O(n14_adj_4987));
    defparam i6_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1686 (.I0(n34405), .I1(n7), .I2(n1_adj_4965), 
            .I3(n4_adj_4866), .O(n37934));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1686.LUT_INIT = 16'hfffd;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n1150), .I1(n1145), .I2(n1149), .I3(n24624), 
            .O(n9_adj_4988));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'heccc;
    SB_LUT4 i30671_4_lut (.I0(n9_adj_4988), .I1(n14_adj_4987), .I2(n1142), 
            .I3(n1143), .O(n1168));
    defparam i30671_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1483_3_lut (.I0(n1168), .I1(n5814), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1483_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i679_3_lut (.I0(n991), .I1(n1044), 
            .I2(n1012), .I3(GND_net), .O(n1069));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i679_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i676_3_lut (.I0(n988), .I1(n1041), 
            .I2(n1012), .I3(GND_net), .O(n1066));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i677_3_lut (.I0(n989), .I1(n1042), 
            .I2(n1012), .I3(GND_net), .O(n1067));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i677_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n18163), 
            .D(n594), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder0_position_23__I_0_i682_3_lut (.I0(n994), .I1(n1047), 
            .I2(n1012), .I3(GND_net), .O(n1072));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i682_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13874_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n34304), .I3(GND_net), .O(n18663));   // verilog/coms.v(127[12] 300[6])
    defparam i13874_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13875_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n34304), .I3(GND_net), .O(n18664));   // verilog/coms.v(127[12] 300[6])
    defparam i13875_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i680_3_lut (.I0(n992), .I1(n1045), 
            .I2(n1012), .I3(GND_net), .O(n1070));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i680_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i681_3_lut (.I0(n993), .I1(n1046), 
            .I2(n1012), .I3(GND_net), .O(n1071));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13876_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n34304), .I3(GND_net), .O(n18665));   // verilog/coms.v(127[12] 300[6])
    defparam i13876_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13877_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n34304), .I3(GND_net), .O(n18666));   // verilog/coms.v(127[12] 300[6])
    defparam i13877_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i678_3_lut (.I0(n990), .I1(n1043), 
            .I2(n1012), .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i674_3_lut (.I0(n986), .I1(n1039), 
            .I2(n1012), .I3(GND_net), .O(n1064));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i675_3_lut (.I0(n987), .I1(n1040), 
            .I2(n1012), .I3(GND_net), .O(n1065));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13878_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n34304), .I3(GND_net), .O(n18667));   // verilog/coms.v(127[12] 300[6])
    defparam i13878_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i684_3_lut (.I0(n519), .I1(n1049), 
            .I2(n1012), .I3(GND_net), .O(n1074));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i684_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_513_3_lut (.I0(GND_net), .I1(n758), 
            .I2(VCC_net), .I3(n28031), .O(n811)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i683_3_lut (.I0(n995), .I1(n1048), 
            .I2(n1012), .I3(GND_net), .O(n1073));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4907), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n763));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19683_3_lut (.I0(n763), .I1(n1073), .I2(n1074), .I3(GND_net), 
            .O(n24462));
    defparam i19683_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13879_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n34304), .I3(GND_net), .O(n18668));   // verilog/coms.v(127[12] 300[6])
    defparam i13879_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13880_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n34304), .I3(GND_net), .O(n18669));   // verilog/coms.v(127[12] 300[6])
    defparam i13880_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13881_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n34304), .I3(GND_net), .O(n18670));   // verilog/coms.v(127[12] 300[6])
    defparam i13881_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1688 (.I0(n1071), .I1(n1070), .I2(n24462), .I3(n1072), 
            .O(n33924));
    defparam i2_4_lut_adj_1688.LUT_INIT = 16'h8880;
    SB_LUT4 i13882_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n34304), .I3(GND_net), .O(n18671));   // verilog/coms.v(127[12] 300[6])
    defparam i13882_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i5_4_lut (.I0(n1065), .I1(n1064), .I2(n33924), .I3(n1068), 
            .O(n12_adj_5061));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30654_4_lut (.I0(n1067), .I1(n12_adj_5061), .I2(n1066), .I3(n1069), 
            .O(n1090));
    defparam i30654_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_23__I_0_add_513_3 (.CI(n28031), .I0(n758), 
            .I1(VCC_net), .CO(n28032));
    SB_LUT4 encoder0_position_23__I_0_add_513_2_lut (.I0(GND_net), .I1(n516), 
            .I2(GND_net), .I3(VCC_net), .O(n812)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1482_3_lut (.I0(n1090), .I1(n5813), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1482_3_lut.LUT_INIT = 16'hc5c5;
    SB_CARRY encoder0_position_23__I_0_add_513_2 (.CI(VCC_net), .I0(n516), 
            .I1(GND_net), .CO(n28031));
    SB_LUT4 encoder0_position_23__I_0_i621_3_lut (.I0(n908), .I1(n961), 
            .I2(n934), .I3(GND_net), .O(n986));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13883_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n34304), .I3(GND_net), .O(n18672));   // verilog/coms.v(127[12] 300[6])
    defparam i13883_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13884_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n34304), .I3(GND_net), .O(n18673));   // verilog/coms.v(127[12] 300[6])
    defparam i13884_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i622_3_lut (.I0(n909), .I1(n962), 
            .I2(n934), .I3(GND_net), .O(n987));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i622_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13885_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n34304), .I3(GND_net), .O(n18674));   // verilog/coms.v(127[12] 300[6])
    defparam i13885_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13886_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n34304), .I3(GND_net), .O(n18675));   // verilog/coms.v(127[12] 300[6])
    defparam i13886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i630_3_lut (.I0(n518), .I1(n970), 
            .I2(n934), .I3(GND_net), .O(n995));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i630_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i629_3_lut (.I0(n916), .I1(n969), 
            .I2(n934), .I3(GND_net), .O(n994));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i629_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i628_3_lut (.I0(n915), .I1(n968), 
            .I2(n934), .I3(GND_net), .O(n993));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i628_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4908), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13887_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n34304), .I3(GND_net), .O(n18676));   // verilog/coms.v(127[12] 300[6])
    defparam i13887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i626_3_lut (.I0(n913), .I1(n966), 
            .I2(n934), .I3(GND_net), .O(n991));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i626_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13888_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n34304), .I3(GND_net), .O(n18677));   // verilog/coms.v(127[12] 300[6])
    defparam i13888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i627_3_lut (.I0(n914), .I1(n967), 
            .I2(n934), .I3(GND_net), .O(n992));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i627_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i625_3_lut (.I0(n912), .I1(n965), 
            .I2(n934), .I3(GND_net), .O(n990));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i623_3_lut (.I0(n910), .I1(n963), 
            .I2(n934), .I3(GND_net), .O(n988));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i623_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_72_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[5]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_i624_3_lut (.I0(n911), .I1(n964), 
            .I2(n934), .I3(GND_net), .O(n989));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i624_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19848_4_lut (.I0(n519), .I1(n993), .I2(n994), .I3(n995), 
            .O(n24630));
    defparam i19848_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_2_lut_adj_1689 (.I0(n989), .I1(n988), .I2(GND_net), .I3(GND_net), 
            .O(n8_adj_4989));
    defparam i2_2_lut_adj_1689.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n990), .I1(n992), .I2(n991), .I3(n24630), 
            .O(n7_adj_4990));
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'heaaa;
    SB_LUT4 i30638_4_lut (.I0(n987), .I1(n7_adj_4990), .I2(n986), .I3(n8_adj_4989), 
            .O(n1012));
    defparam i30638_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_70_i6_3_lut (.I0(encoder0_position_scaled[5]), .I1(motor_state_23__N_82[5]), 
            .I2(n15), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_23__I_0_i1481_3_lut (.I0(n1012), .I1(n5812), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1481_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i570_3_lut (.I0(n832), .I1(n885), 
            .I2(n856), .I3(GND_net), .O(n910));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i569_3_lut (.I0(n831), .I1(n884), 
            .I2(n856), .I3(GND_net), .O(n909));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i571_3_lut (.I0(n833), .I1(n886), 
            .I2(n856), .I3(GND_net), .O(n911));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i571_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i576_3_lut (.I0(n517), .I1(n891), 
            .I2(n856), .I3(GND_net), .O(n916));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i575_3_lut (.I0(n837), .I1(n890), 
            .I2(n856), .I3(GND_net), .O(n915));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i575_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n18163), 
            .D(n593), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder0_position_23__I_0_i574_3_lut (.I0(n836), .I1(n889), 
            .I2(n856), .I3(GND_net), .O(n914));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13889_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n34304), .I3(GND_net), .O(n18678));   // verilog/coms.v(127[12] 300[6])
    defparam i13889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_1691 (.I0(ID[7]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_4891));   // verilog/TinyFPGA_B.v(252[12:17])
    defparam i6_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_3291_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4909), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i572_3_lut (.I0(n834), .I1(n887), 
            .I2(n856), .I3(GND_net), .O(n912));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i572_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[0]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFFESR delay_counter_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n18163), 
            .D(n592), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder0_position_23__I_0_i568_3_lut (.I0(n830), .I1(n883), 
            .I2(n856), .I3(GND_net), .O(n908));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i568_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n18163), 
            .D(n591), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i7_4_lut_adj_1692 (.I0(ID[0]), .I1(n14_adj_4891), .I2(n10_adj_4892), 
            .I3(ID[3]), .O(n15_adj_4867));   // verilog/TinyFPGA_B.v(252[12:17])
    defparam i7_4_lut_adj_1692.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i573_3_lut (.I0(n835), .I1(n888), 
            .I2(n856), .I3(GND_net), .O(n913));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19852_4_lut (.I0(n518), .I1(n914), .I2(n915), .I3(n916), 
            .O(n24634));
    defparam i19852_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1693 (.I0(n913), .I1(n908), .I2(n912), .I3(n24634), 
            .O(n7_adj_4880));
    defparam i2_4_lut_adj_1693.LUT_INIT = 16'heccc;
    SB_DFFESR delay_counter_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n18163), 
            .D(n590), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 i30623_4_lut (.I0(n7_adj_4880), .I1(n911), .I2(n909), .I3(n910), 
            .O(n934));
    defparam i30623_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1480_3_lut (.I0(n934), .I1(n5811), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1480_3_lut.LUT_INIT = 16'hc5c5;
    SB_DFFESR delay_counter_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n18163), 
            .D(n589), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[6]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i7_3_lut (.I0(encoder0_position_scaled[6]), .I1(motor_state_23__N_82[6]), 
            .I2(n15), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i7_4_lut_adj_1694 (.I0(delay_counter[3]), .I1(delay_counter[9]), 
            .I2(delay_counter[8]), .I3(delay_counter[5]), .O(n18_adj_5042));
    defparam i7_4_lut_adj_1694.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1695 (.I0(delay_counter[1]), .I1(n18_adj_5042), 
            .I2(delay_counter[2]), .I3(delay_counter[6]), .O(n20_adj_5040));
    defparam i9_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1696 (.I0(delay_counter[10]), .I1(delay_counter[0]), 
            .I2(delay_counter[7]), .I3(delay_counter[4]), .O(n19_adj_5041));
    defparam i8_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i1891_4_lut (.I0(n19_adj_5041), .I1(delay_counter[12]), .I2(delay_counter[11]), 
            .I3(n20_adj_5040), .O(n26_adj_4963));
    defparam i1891_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[7]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1894_4_lut (.I0(n26_adj_4963), .I1(delay_counter[15]), .I2(delay_counter[14]), 
            .I3(delay_counter[13]), .O(n32_adj_4964));
    defparam i1894_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 mux_70_i8_3_lut (.I0(encoder0_position_scaled[7]), .I1(motor_state_23__N_82[7]), 
            .I2(n15), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i8_3_lut.LUT_INIT = 16'h3535;
    SB_DFF h1_47 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_23__I_0_i516_3_lut (.I0(n753), .I1(n806), 
            .I2(n778), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i517_3_lut (.I0(n754), .I1(n807), 
            .I2(n778), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13890_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n34304), .I3(GND_net), .O(n18679));   // verilog/coms.v(127[12] 300[6])
    defparam i13890_3_lut.LUT_INIT = 16'hacac;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFFESR delay_counter_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n18163), 
            .D(n588), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder0_position_23__I_0_i520_3_lut (.I0(n757), .I1(n810), 
            .I2(n778), .I3(GND_net), .O(n835));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i518_3_lut (.I0(n755), .I1(n808), 
            .I2(n778), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i519_3_lut (.I0(n756), .I1(n809), 
            .I2(n778), .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i522_3_lut (.I0(n516), .I1(n812), 
            .I2(n778), .I3(GND_net), .O(n837));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1697 (.I0(n32_adj_4964), .I1(delay_counter[18]), 
            .I2(delay_counter[16]), .I3(delay_counter[17]), .O(n33396));
    defparam i2_4_lut_adj_1697.LUT_INIT = 16'hffec;
    SB_LUT4 i2_2_lut_adj_1698 (.I0(delay_counter[20]), .I1(delay_counter[21]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5049));
    defparam i2_2_lut_adj_1698.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_i521_3_lut (.I0(n758), .I1(n811), 
            .I2(n778), .I3(GND_net), .O(n836));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3291_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4910), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n517));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19691_3_lut (.I0(n517), .I1(n836), .I2(n837), .I3(GND_net), 
            .O(n24470));
    defparam i19691_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1699 (.I0(n834), .I1(n833), .I2(n24470), .I3(n835), 
            .O(n33787));
    defparam i2_4_lut_adj_1699.LUT_INIT = 16'h8880;
    SB_LUT4 i30572_4_lut (.I0(n33787), .I1(n830), .I2(n832), .I3(n831), 
            .O(n856));
    defparam i30572_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1479_3_lut (.I0(n856), .I1(n5810), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1479_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1478_3_lut (.I0(n778), .I1(n5809), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1478_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1477_3_lut (.I0(n700), .I1(n5808), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1477_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 add_28_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n27637), .O(n615)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n18163), 
            .D(n587), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 mux_72_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[8]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i9_3_lut (.I0(encoder0_position_scaled[8]), .I1(motor_state_23__N_82[8]), 
            .I2(n15), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13898_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n34304), .I3(GND_net), .O(n18687));   // verilog/coms.v(127[12] 300[6])
    defparam i13898_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13899_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n34304), .I3(GND_net), .O(n18688));   // verilog/coms.v(127[12] 300[6])
    defparam i13899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13900_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n34304), .I3(GND_net), .O(n18689));   // verilog/coms.v(127[12] 300[6])
    defparam i13900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13901_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n34304), .I3(GND_net), .O(n18690));   // verilog/coms.v(127[12] 300[6])
    defparam i13901_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13902_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n34304), .I3(GND_net), .O(n18691));   // verilog/coms.v(127[12] 300[6])
    defparam i13902_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13903_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n34304), .I3(GND_net), .O(n18692));   // verilog/coms.v(127[12] 300[6])
    defparam i13903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1700 (.I0(n33396), .I1(delay_counter[22]), .I2(delay_counter[19]), 
            .I3(GND_net), .O(n5_adj_5050));
    defparam i1_3_lut_adj_1700.LUT_INIT = 16'hecec;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_4995), .I3(n28621), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_4996), .I3(n28620), .O(n3_adj_4917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_25 (.CI(n28620), 
            .I0(GND_net), .I1(n3_adj_4996), .CO(n28621));
    SB_LUT4 mux_72_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[9]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i10_3_lut (.I0(encoder0_position_scaled[9]), .I1(motor_state_23__N_82[9]), 
            .I2(n15), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_4997), .I3(n28619), .O(n4_adj_4916)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_24 (.CI(n28619), 
            .I0(GND_net), .I1(n4_adj_4997), .CO(n28620));
    SB_LUT4 i13891_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n34304), .I3(GND_net), .O(n18680));   // verilog/coms.v(127[12] 300[6])
    defparam i13891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_4998), .I3(n28618), .O(n5_adj_4915)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_23 (.CI(n28618), 
            .I0(GND_net), .I1(n5_adj_4998), .CO(n28619));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_4999), .I3(n28617), .O(n6_adj_4914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_22 (.CI(n28617), 
            .I0(GND_net), .I1(n6_adj_4999), .CO(n28618));
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4869));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13892_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n34304), .I3(GND_net), .O(n18681));   // verilog/coms.v(127[12] 300[6])
    defparam i13892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13893_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n34304), .I3(GND_net), .O(n18682));   // verilog/coms.v(127[12] 300[6])
    defparam i13893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13904_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n32403), .I3(GND_net), .O(n18693));   // verilog/coms.v(127[12] 300[6])
    defparam i13904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13908_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n32403), .I3(GND_net), .O(n18697));   // verilog/coms.v(127[12] 300[6])
    defparam i13908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_5000), .I3(n28616), .O(n7_adj_4913)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13909_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n32403), .I3(GND_net), .O(n18698));   // verilog/coms.v(127[12] 300[6])
    defparam i13909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13910_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n32403), .I3(GND_net), .O(n18699));   // verilog/coms.v(127[12] 300[6])
    defparam i13910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13911_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n32403), .I3(GND_net), .O(n18700));   // verilog/coms.v(127[12] 300[6])
    defparam i13911_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_21 (.CI(n28616), 
            .I0(GND_net), .I1(n7_adj_5000), .CO(n28617));
    SB_LUT4 i13912_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n32403), .I3(GND_net), .O(n18701));   // verilog/coms.v(127[12] 300[6])
    defparam i13912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13894_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n34304), .I3(GND_net), .O(n18683));   // verilog/coms.v(127[12] 300[6])
    defparam i13894_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_5001), .I3(n28615), .O(n8_adj_4912)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13913_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n32403), .I3(GND_net), .O(n18702));   // verilog/coms.v(127[12] 300[6])
    defparam i13913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13914_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n32403), .I3(GND_net), .O(n18703));   // verilog/coms.v(127[12] 300[6])
    defparam i13914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_28_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n27645), .O(n607)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_20 (.CI(n28615), 
            .I0(GND_net), .I1(n8_adj_5001), .CO(n28616));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_5002), .I3(n28614), .O(n9_adj_4911)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_19 (.CI(n28614), 
            .I0(GND_net), .I1(n9_adj_5002), .CO(n28615));
    SB_LUT4 encoder0_position_23__I_0_add_460_8_lut (.I0(n37245), .I1(n674), 
            .I2(VCC_net), .I3(n28021), .O(n752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_5003), .I3(n28613), .O(n10_adj_4910)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_18 (.CI(n28613), 
            .I0(GND_net), .I1(n10_adj_5003), .CO(n28614));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5004), .I3(n28612), .O(n11_adj_4909)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_13 (.CI(n27645), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n27646));
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_28_5 (.CI(n27637), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n27638));
    SB_LUT4 encoder0_position_23__I_0_add_460_7_lut (.I0(GND_net), .I1(n675), 
            .I2(GND_net), .I3(n28020), .O(n728)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_17 (.CI(n28612), 
            .I0(GND_net), .I1(n11_adj_5004), .CO(n28613));
    SB_CARRY encoder0_position_23__I_0_add_460_7 (.CI(n28020), .I0(n675), 
            .I1(GND_net), .CO(n28021));
    SB_LUT4 i13923_3_lut (.I0(\data_in_frame[19] [7]), .I1(rx_data[7]), 
            .I2(n32402), .I3(GND_net), .O(n18712));   // verilog/coms.v(127[12] 300[6])
    defparam i13923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13924_3_lut (.I0(\data_in_frame[19] [6]), .I1(rx_data[6]), 
            .I2(n32402), .I3(GND_net), .O(n18713));   // verilog/coms.v(127[12] 300[6])
    defparam i13924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5005), .I3(n28611), .O(n12_adj_4908)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_16 (.CI(n28611), 
            .I0(GND_net), .I1(n12_adj_5005), .CO(n28612));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5006), .I3(n28610), .O(n13_adj_4907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_15 (.CI(n28610), 
            .I0(GND_net), .I1(n13_adj_5006), .CO(n28611));
    SB_LUT4 i13925_3_lut (.I0(\data_in_frame[19] [5]), .I1(rx_data[5]), 
            .I2(n32402), .I3(GND_net), .O(n18714));   // verilog/coms.v(127[12] 300[6])
    defparam i13925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_4_lut_adj_1701 (.I0(n5_adj_5050), .I1(delay_counter[24]), 
            .I2(n6_adj_5049), .I3(delay_counter[23]), .O(n33948));
    defparam i2_4_lut_adj_1701.LUT_INIT = 16'hc800;
    SB_LUT4 encoder0_position_23__I_0_add_460_6_lut (.I0(GND_net), .I1(n676), 
            .I2(GND_net), .I3(n28019), .O(n729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_6 (.CI(n28019), .I0(n676), 
            .I1(GND_net), .CO(n28020));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5007), .I3(n28609), .O(n14_adj_4906)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_14 (.CI(n28609), 
            .I0(GND_net), .I1(n14_adj_5007), .CO(n28610));
    SB_LUT4 i13926_3_lut (.I0(\data_in_frame[19] [4]), .I1(rx_data[4]), 
            .I2(n32402), .I3(GND_net), .O(n18715));   // verilog/coms.v(127[12] 300[6])
    defparam i13926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13927_3_lut (.I0(\data_in_frame[19] [3]), .I1(rx_data[3]), 
            .I2(n32402), .I3(GND_net), .O(n18716));   // verilog/coms.v(127[12] 300[6])
    defparam i13927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13928_3_lut (.I0(\data_in_frame[19] [2]), .I1(rx_data[2]), 
            .I2(n32402), .I3(GND_net), .O(n18717));   // verilog/coms.v(127[12] 300[6])
    defparam i13928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5008), .I3(n28608), .O(n15_adj_4905)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_460_5_lut (.I0(GND_net), .I1(n677), 
            .I2(VCC_net), .I3(n28018), .O(n730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_13 (.CI(n28608), 
            .I0(GND_net), .I1(n15_adj_5008), .CO(n28609));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5009), .I3(n28607), .O(n16_adj_4904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13929_3_lut (.I0(\data_in_frame[19] [1]), .I1(rx_data[1]), 
            .I2(n32402), .I3(GND_net), .O(n18718));   // verilog/coms.v(127[12] 300[6])
    defparam i13929_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_460_5 (.CI(n28018), .I0(n677), 
            .I1(VCC_net), .CO(n28019));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_12 (.CI(n28607), 
            .I0(GND_net), .I1(n16_adj_5009), .CO(n28608));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5010), .I3(n28606), .O(n17_adj_4903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_11 (.CI(n28606), 
            .I0(GND_net), .I1(n17_adj_5010), .CO(n28607));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5011), .I3(n28605), .O(n18_adj_4902)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_10 (.CI(n28605), 
            .I0(GND_net), .I1(n18_adj_5011), .CO(n28606));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5012), .I3(n28604), .O(n19_adj_4901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_9 (.CI(n28604), 
            .I0(GND_net), .I1(n19_adj_5012), .CO(n28605));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5013), .I3(n28603), .O(n20_adj_4900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_460_4_lut (.I0(GND_net), .I1(n678), 
            .I2(GND_net), .I3(n28017), .O(n731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13930_3_lut (.I0(\data_in_frame[19] [0]), .I1(rx_data[0]), 
            .I2(n32402), .I3(GND_net), .O(n18719));   // verilog/coms.v(127[12] 300[6])
    defparam i13930_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_8 (.CI(n28603), 
            .I0(GND_net), .I1(n20_adj_5013), .CO(n28604));
    SB_CARRY encoder0_position_23__I_0_add_460_4 (.CI(n28017), .I0(n678), 
            .I1(GND_net), .CO(n28018));
    SB_LUT4 i13931_3_lut (.I0(\data_in_frame[18] [7]), .I1(rx_data[7]), 
            .I2(n32385), .I3(GND_net), .O(n18720));   // verilog/coms.v(127[12] 300[6])
    defparam i13931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5014), .I3(n28602), .O(n21_adj_4899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13932_3_lut (.I0(\data_in_frame[18] [6]), .I1(rx_data[6]), 
            .I2(n32385), .I3(GND_net), .O(n18721));   // verilog/coms.v(127[12] 300[6])
    defparam i13932_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_7 (.CI(n28602), 
            .I0(GND_net), .I1(n21_adj_5014), .CO(n28603));
    SB_LUT4 i13933_3_lut (.I0(\data_in_frame[18] [5]), .I1(rx_data[5]), 
            .I2(n32385), .I3(GND_net), .O(n18722));   // verilog/coms.v(127[12] 300[6])
    defparam i13933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13934_3_lut (.I0(\data_in_frame[18] [4]), .I1(rx_data[4]), 
            .I2(n32385), .I3(GND_net), .O(n18723));   // verilog/coms.v(127[12] 300[6])
    defparam i13934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13935_3_lut (.I0(\data_in_frame[18] [3]), .I1(rx_data[3]), 
            .I2(n32385), .I3(GND_net), .O(n18724));   // verilog/coms.v(127[12] 300[6])
    defparam i13935_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13936_3_lut (.I0(\data_in_frame[18] [2]), .I1(rx_data[2]), 
            .I2(n32385), .I3(GND_net), .O(n18725));   // verilog/coms.v(127[12] 300[6])
    defparam i13936_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_460_3_lut (.I0(GND_net), .I1(n679), 
            .I2(VCC_net), .I3(n28016), .O(n732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5015), .I3(n28601), .O(n22_adj_4898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_6 (.CI(n28601), 
            .I0(GND_net), .I1(n22_adj_5015), .CO(n28602));
    SB_LUT4 i13937_3_lut (.I0(\data_in_frame[18] [1]), .I1(rx_data[1]), 
            .I2(n32385), .I3(GND_net), .O(n18726));   // verilog/coms.v(127[12] 300[6])
    defparam i13937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13938_3_lut (.I0(\data_in_frame[18] [0]), .I1(rx_data[0]), 
            .I2(n32385), .I3(GND_net), .O(n18727));   // verilog/coms.v(127[12] 300[6])
    defparam i13938_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13939_3_lut (.I0(\data_in_frame[17] [7]), .I1(rx_data[7]), 
            .I2(n32400), .I3(GND_net), .O(n18728));   // verilog/coms.v(127[12] 300[6])
    defparam i13939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13940_3_lut (.I0(\data_in_frame[17] [6]), .I1(rx_data[6]), 
            .I2(n32400), .I3(GND_net), .O(n18729));   // verilog/coms.v(127[12] 300[6])
    defparam i13940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13941_3_lut (.I0(\data_in_frame[17] [5]), .I1(rx_data[5]), 
            .I2(n32400), .I3(GND_net), .O(n18730));   // verilog/coms.v(127[12] 300[6])
    defparam i13941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13942_3_lut (.I0(\data_in_frame[17] [4]), .I1(rx_data[4]), 
            .I2(n32400), .I3(GND_net), .O(n18731));   // verilog/coms.v(127[12] 300[6])
    defparam i13942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_72_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[10]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i11_3_lut (.I0(encoder0_position_scaled[10]), .I1(motor_state_23__N_82[10]), 
            .I2(n15), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13943_3_lut (.I0(\data_in_frame[17] [3]), .I1(rx_data[3]), 
            .I2(n32400), .I3(GND_net), .O(n18732));   // verilog/coms.v(127[12] 300[6])
    defparam i13943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13944_3_lut (.I0(\data_in_frame[17] [2]), .I1(rx_data[2]), 
            .I2(n32400), .I3(GND_net), .O(n18733));   // verilog/coms.v(127[12] 300[6])
    defparam i13944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13945_3_lut (.I0(\data_in_frame[17] [1]), .I1(rx_data[1]), 
            .I2(n32400), .I3(GND_net), .O(n18734));   // verilog/coms.v(127[12] 300[6])
    defparam i13945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13946_3_lut (.I0(\data_in_frame[17] [0]), .I1(rx_data[0]), 
            .I2(n32400), .I3(GND_net), .O(n18735));   // verilog/coms.v(127[12] 300[6])
    defparam i13946_3_lut.LUT_INIT = 16'hacac;
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_732_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4971));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i9_2_lut.LUT_INIT = 16'h6666;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 LessThan_732_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4973));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4977));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4982));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1702 (.I0(delay_counter[28]), .I1(delay_counter[29]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_5048));
    defparam i2_2_lut_adj_1702.LUT_INIT = 16'heeee;
    SB_LUT4 LessThan_732_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4976));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4975));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4969));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4979));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4980));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4978));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4983));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4985));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4986));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_732_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4981));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3330_4_lut (.I0(n33948), .I1(delay_counter[27]), .I2(delay_counter[26]), 
            .I3(delay_counter[25]), .O(n56));
    defparam i3330_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 LessThan_732_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5016), .I3(n28600), .O(n23_adj_4897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_5 (.CI(n28600), 
            .I0(GND_net), .I1(n23_adj_5016), .CO(n28601));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5017), .I3(n28599), .O(n24_adj_4896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_4 (.CI(n28599), 
            .I0(GND_net), .I1(n24_adj_5017), .CO(n28600));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5018), .I3(n28598), .O(n25_adj_4895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_3 (.CI(n28598), 
            .I0(GND_net), .I1(n25_adj_5018), .CO(n28599));
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n28598));
    SB_CARRY encoder0_position_23__I_0_add_460_3 (.CI(n28016), .I0(n679), 
            .I1(VCC_net), .CO(n28017));
    SB_LUT4 i19011_4_lut (.I0(n56), .I1(delay_counter[31]), .I2(n6_adj_5048), 
            .I3(delay_counter[30]), .O(n619));   // verilog/TinyFPGA_B.v(254[14:40])
    defparam i19011_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i13729_2_lut (.I0(n18163), .I1(n619), .I2(GND_net), .I3(GND_net), 
            .O(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i13729_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_23__I_0_add_460_2_lut (.I0(GND_net), .I1(n515), 
            .I2(GND_net), .I3(VCC_net), .O(n733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_72_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[11]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i12_3_lut (.I0(encoder0_position_scaled[11]), .I1(motor_state_23__N_82[11]), 
            .I2(n15), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i12_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_23__I_0_add_460_2 (.CI(VCC_net), .I0(n515), 
            .I1(GND_net), .CO(n28016));
    SB_LUT4 i13974_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n32412), .I3(GND_net), .O(n18763));   // verilog/coms.v(127[12] 300[6])
    defparam i13974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13975_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n32412), .I3(GND_net), .O(n18764));   // verilog/coms.v(127[12] 300[6])
    defparam i13975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_72_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[12]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_660_24_lut (.I0(duty[22]), .I1(n37310), .I2(n3), .I3(n27749), 
            .O(pwm_setpoint_22__N_11[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13976_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n32412), .I3(GND_net), .O(n18765));   // verilog/coms.v(127[12] 300[6])
    defparam i13976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_660_23_lut (.I0(duty[21]), .I1(n37310), .I2(n4_adj_4868), 
            .I3(n27748), .O(pwm_setpoint_22__N_11[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_70_i13_3_lut (.I0(encoder0_position_scaled[12]), .I1(motor_state_23__N_82[12]), 
            .I2(n15), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i13_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY add_660_23 (.CI(n27748), .I0(n37310), .I1(n4_adj_4868), .CO(n27749));
    SB_LUT4 i13836_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n2134), .I3(GND_net), .O(n18625));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13836_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13977_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n32412), .I3(GND_net), .O(n18766));   // verilog/coms.v(127[12] 300[6])
    defparam i13977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13978_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n32412), .I3(GND_net), .O(n18767));   // verilog/coms.v(127[12] 300[6])
    defparam i13978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_660_22_lut (.I0(duty[20]), .I1(n37310), .I2(n5), .I3(n27747), 
            .O(pwm_setpoint_22__N_11[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_i1495_3_lut (.I0(n24674), .I1(n5826), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1495_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i13979_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n32412), .I3(GND_net), .O(n18768));   // verilog/coms.v(127[12] 300[6])
    defparam i13979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13980_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n32412), .I3(GND_net), .O(n18769));   // verilog/coms.v(127[12] 300[6])
    defparam i13980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13981_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n32412), .I3(GND_net), .O(n18770));   // verilog/coms.v(127[12] 300[6])
    defparam i13981_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_58[23]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_CARRY add_660_22 (.CI(n27747), .I0(n37310), .I1(n5), .CO(n27748));
    SB_LUT4 add_660_21_lut (.I0(duty[19]), .I1(n37310), .I2(n6), .I3(n27746), 
            .O(pwm_setpoint_22__N_11[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_21 (.CI(n27746), .I0(n37310), .I1(n6), .CO(n27747));
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_58[22]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_58[21]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_58[20]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_58[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_58[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_58[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_58[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_58[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_58[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_58[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_58[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_58[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_58[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_58[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_58[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_58[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_58[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_58[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_58[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_58[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_58[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_58[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 mux_72_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[13]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i14_3_lut (.I0(encoder0_position_scaled[13]), .I1(motor_state_23__N_82[13]), 
            .I2(n15), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i14_3_lut.LUT_INIT = 16'h3535;
    SB_DFFSR encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
            .C(clk32MHz), .D(n5805), .R(n2_adj_4995));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 add_660_20_lut (.I0(duty[18]), .I1(n37310), .I2(n7_adj_4869), 
            .I3(n27745), .O(pwm_setpoint_22__N_11[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_72_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[14]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i15_3_lut (.I0(encoder0_position_scaled[14]), .I1(motor_state_23__N_82[14]), 
            .I2(n15), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i15_3_lut.LUT_INIT = 16'h3535;
    SB_DFFSR encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
            .C(clk32MHz), .D(n5806), .R(n2_adj_4995));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i13990_3_lut (.I0(\data_in_frame[11] [7]), .I1(rx_data[7]), 
            .I2(n32410), .I3(GND_net), .O(n18779));   // verilog/coms.v(127[12] 300[6])
    defparam i13990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13895_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n34304), .I3(GND_net), .O(n18684));   // verilog/coms.v(127[12] 300[6])
    defparam i13895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_72_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[15]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i16_3_lut (.I0(encoder0_position_scaled[15]), .I1(motor_state_23__N_82[15]), 
            .I2(n15), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_72_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[16]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i17_3_lut (.I0(encoder0_position_scaled[16]), .I1(motor_state_23__N_82[16]), 
            .I2(n15), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13991_3_lut (.I0(\data_in_frame[11] [6]), .I1(rx_data[6]), 
            .I2(n32410), .I3(GND_net), .O(n18780));   // verilog/coms.v(127[12] 300[6])
    defparam i13991_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[17]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i18_3_lut (.I0(encoder0_position_scaled[17]), .I1(motor_state_23__N_82[17]), 
            .I2(n15), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13992_3_lut (.I0(\data_in_frame[11] [5]), .I1(rx_data[5]), 
            .I2(n32410), .I3(GND_net), .O(n18781));   // verilog/coms.v(127[12] 300[6])
    defparam i13992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13993_3_lut (.I0(\data_in_frame[11] [4]), .I1(rx_data[4]), 
            .I2(n32410), .I3(GND_net), .O(n18782));   // verilog/coms.v(127[12] 300[6])
    defparam i13993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4958));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[18]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i19_3_lut (.I0(encoder0_position_scaled[18]), .I1(motor_state_23__N_82[18]), 
            .I2(n15), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 add_28_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n27644), .O(n608)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4957));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13994_3_lut (.I0(\data_in_frame[11] [3]), .I1(rx_data[3]), 
            .I2(n32410), .I3(GND_net), .O(n18783));   // verilog/coms.v(127[12] 300[6])
    defparam i13994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13995_3_lut (.I0(\data_in_frame[11] [2]), .I1(rx_data[2]), 
            .I2(n32410), .I3(GND_net), .O(n18784));   // verilog/coms.v(127[12] 300[6])
    defparam i13995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13996_3_lut (.I0(\data_in_frame[11] [1]), .I1(rx_data[1]), 
            .I2(n32410), .I3(GND_net), .O(n18785));   // verilog/coms.v(127[12] 300[6])
    defparam i13996_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_660_20 (.CI(n27745), .I0(n37310), .I1(n7_adj_4869), .CO(n27746));
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(143[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i13997_3_lut (.I0(\data_in_frame[11] [0]), .I1(rx_data[0]), 
            .I2(n32410), .I3(GND_net), .O(n18786));   // verilog/coms.v(127[12] 300[6])
    defparam i13997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_660_19_lut (.I0(duty[17]), .I1(n37310), .I2(n8), .I3(n27744), 
            .O(pwm_setpoint_22__N_11[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_19 (.CI(n27744), .I0(n37310), .I1(n8), .CO(n27745));
    SB_LUT4 i3360_3_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n619), .I3(n15_adj_4867), .O(n5131));   // verilog/TinyFPGA_B.v(251[7:11])
    defparam i3360_3_lut_3_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 add_660_18_lut (.I0(duty[16]), .I1(n37310), .I2(n9), .I3(n27743), 
            .O(pwm_setpoint_22__N_11[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_18 (.CI(n27743), .I0(n37310), .I1(n9), .CO(n27744));
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[22]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[21]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[20]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[19]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[18]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[17]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[16]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[15]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[14]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[13]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[12]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[11]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[10]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[9]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[8]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[7]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[6]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[5]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[4]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[3]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[2]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[1]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 LessThan_732_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4968));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_732_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4972));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_660_17_lut (.I0(duty[15]), .I1(n37310), .I2(n10), .I3(n27742), 
            .O(pwm_setpoint_22__N_11[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n3_adj_4937), .I3(n27998), .O(displacement_23__N_58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29603_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n35999));
    defparam i29603_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_732_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4974));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_732_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4970));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4937), .I3(n27997), .O(displacement_23__N_58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29617_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n36013));
    defparam i29617_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n27997), .I0(encoder1_position[22]), 
            .I1(n3_adj_4937), .CO(n27998));
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n3_adj_4937), .I3(n27996), .O(displacement_23__N_58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14006_3_lut (.I0(\data_in_frame[9] [7]), .I1(rx_data[7]), .I2(n32409), 
            .I3(GND_net), .O(n18795));   // verilog/coms.v(127[12] 300[6])
    defparam i14006_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_660_17 (.CI(n27742), .I0(n37310), .I1(n10), .CO(n27743));
    SB_LUT4 i14007_3_lut (.I0(\data_in_frame[9] [6]), .I1(rx_data[6]), .I2(n32409), 
            .I3(GND_net), .O(n18796));   // verilog/coms.v(127[12] 300[6])
    defparam i14007_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n27996), .I0(encoder1_position[21]), 
            .I1(n3_adj_4937), .CO(n27997));
    SB_LUT4 i14008_3_lut (.I0(\data_in_frame[9] [5]), .I1(rx_data[5]), .I2(n32409), 
            .I3(GND_net), .O(n18797));   // verilog/coms.v(127[12] 300[6])
    defparam i14008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4938), .I3(n27995), .O(displacement_23__N_58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n27995), .I0(encoder1_position[20]), 
            .I1(n5_adj_4938), .CO(n27996));
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4939), .I3(n27994), .O(displacement_23__N_58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n27994), .I0(encoder1_position[19]), 
            .I1(n6_adj_4939), .CO(n27995));
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4940), .I3(n27993), .O(displacement_23__N_58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14009_3_lut (.I0(\data_in_frame[9] [4]), .I1(rx_data[4]), .I2(n32409), 
            .I3(GND_net), .O(n18798));   // verilog/coms.v(127[12] 300[6])
    defparam i14009_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_660_16_lut (.I0(duty[14]), .I1(n37310), .I2(n11), .I3(n27741), 
            .O(pwm_setpoint_22__N_11[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_16 (.CI(n27741), .I0(n37310), .I1(n11), .CO(n27742));
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n27993), .I0(encoder1_position[18]), 
            .I1(n7_adj_4940), .CO(n27994));
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4941), .I3(n27992), .O(displacement_23__N_58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n27992), .I0(encoder1_position[17]), 
            .I1(n8_adj_4941), .CO(n27993));
    SB_LUT4 add_660_15_lut (.I0(duty[13]), .I1(n37310), .I2(n12), .I3(n27740), 
            .O(pwm_setpoint_22__N_11[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14010_3_lut (.I0(\data_in_frame[9] [3]), .I1(rx_data[3]), .I2(n32409), 
            .I3(GND_net), .O(n18799));   // verilog/coms.v(127[12] 300[6])
    defparam i14010_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_660_15 (.CI(n27740), .I0(n37310), .I1(n12), .CO(n27741));
    SB_LUT4 i14011_3_lut (.I0(\data_in_frame[9] [2]), .I1(rx_data[2]), .I2(n32409), 
            .I3(GND_net), .O(n18800));   // verilog/coms.v(127[12] 300[6])
    defparam i14011_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14012_3_lut (.I0(\data_in_frame[9] [1]), .I1(rx_data[1]), .I2(n32409), 
            .I3(GND_net), .O(n18801));   // verilog/coms.v(127[12] 300[6])
    defparam i14012_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14013_3_lut (.I0(\data_in_frame[9] [0]), .I1(rx_data[0]), .I2(n32409), 
            .I3(GND_net), .O(n18802));   // verilog/coms.v(127[12] 300[6])
    defparam i14013_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_660_14_lut (.I0(duty[12]), .I1(n37310), .I2(n13), .I3(n27739), 
            .O(pwm_setpoint_22__N_11[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_14 (.CI(n27739), .I0(n37310), .I1(n13), .CO(n27740));
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4942), .I3(n27991), .O(displacement_23__N_58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n27991), .I0(encoder1_position[16]), 
            .I1(n9_adj_4942), .CO(n27992));
    SB_LUT4 add_660_13_lut (.I0(duty[11]), .I1(n37310), .I2(n14), .I3(n27738), 
            .O(pwm_setpoint_22__N_11[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_13 (.CI(n27738), .I0(n37310), .I1(n14), .CO(n27739));
    SB_LUT4 add_660_12_lut (.I0(duty[10]), .I1(n37310), .I2(n15_adj_4870), 
            .I3(n27737), .O(pwm_setpoint_22__N_11[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_12 (.CI(n27737), .I0(n37310), .I1(n15_adj_4870), 
            .CO(n27738));
    SB_LUT4 add_660_11_lut (.I0(duty[9]), .I1(n37310), .I2(n16_adj_4871), 
            .I3(n27736), .O(pwm_setpoint_22__N_11[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_660_11 (.CI(n27736), .I0(n37310), .I1(n16_adj_4871), 
            .CO(n27737));
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4943), .I3(n27990), .O(displacement_23__N_58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n27990), .I0(encoder1_position[15]), 
            .I1(n10_adj_4943), .CO(n27991));
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4944), .I3(n27989), .O(displacement_23__N_58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_660_10_lut (.I0(duty[8]), .I1(n37310), .I2(n17), .I3(n27735), 
            .O(pwm_setpoint_22__N_11[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n27989), .I0(encoder1_position[14]), 
            .I1(n11_adj_4944), .CO(n27990));
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4945), .I3(n27988), .O(displacement_23__N_58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n27988), .I0(encoder1_position[13]), 
            .I1(n12_adj_4945), .CO(n27989));
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4946), .I3(n27987), .O(displacement_23__N_58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_26_lut (.I0(GND_net), .I1(n2000), 
            .I2(VCC_net), .I3(n28315), .O(n2053)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_25_lut (.I0(GND_net), .I1(n2001), 
            .I2(VCC_net), .I3(n28314), .O(n2054)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_25 (.CI(n28314), .I0(n2001), 
            .I1(VCC_net), .CO(n28315));
    SB_LUT4 encoder0_position_23__I_0_add_1361_24_lut (.I0(GND_net), .I1(n2002), 
            .I2(VCC_net), .I3(n28313), .O(n2055)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_24 (.CI(n28313), .I0(n2002), 
            .I1(VCC_net), .CO(n28314));
    SB_CARRY add_660_10 (.CI(n27735), .I0(n37310), .I1(n17), .CO(n27736));
    SB_LUT4 encoder0_position_23__I_0_add_1361_23_lut (.I0(GND_net), .I1(n2003), 
            .I2(VCC_net), .I3(n28312), .O(n2056)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_23 (.CI(n28312), .I0(n2003), 
            .I1(VCC_net), .CO(n28313));
    SB_LUT4 encoder0_position_23__I_0_add_1361_22_lut (.I0(GND_net), .I1(n2004), 
            .I2(VCC_net), .I3(n28311), .O(n2057)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_22 (.CI(n28311), .I0(n2004), 
            .I1(VCC_net), .CO(n28312));
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n17027), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_4936));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1703 (.I0(control_mode[0]), .I1(n17027), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i1_2_lut_3_lut_adj_1703.LUT_INIT = 16'hfefe;
    SB_CARRY add_28_12 (.CI(n27644), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n27645));
    SB_LUT4 encoder0_position_23__I_0_add_1361_21_lut (.I0(GND_net), .I1(n2005), 
            .I2(VCC_net), .I3(n28310), .O(n2058)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_21 (.CI(n28310), .I0(n2005), 
            .I1(VCC_net), .CO(n28311));
    SB_LUT4 encoder0_position_23__I_0_add_1361_20_lut (.I0(GND_net), .I1(n2006), 
            .I2(VCC_net), .I3(n28309), .O(n2059)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_20 (.CI(n28309), .I0(n2006), 
            .I1(VCC_net), .CO(n28310));
    SB_LUT4 encoder0_position_23__I_0_add_1361_19_lut (.I0(GND_net), .I1(n2007), 
            .I2(VCC_net), .I3(n28308), .O(n2060)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_19 (.CI(n28308), .I0(n2007), 
            .I1(VCC_net), .CO(n28309));
    SB_LUT4 encoder0_position_23__I_0_add_1361_18_lut (.I0(GND_net), .I1(n2008), 
            .I2(VCC_net), .I3(n28307), .O(n2061)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_18 (.CI(n28307), .I0(n2008), 
            .I1(VCC_net), .CO(n28308));
    SB_LUT4 encoder0_position_23__I_0_add_1361_17_lut (.I0(GND_net), .I1(n2009), 
            .I2(VCC_net), .I3(n28306), .O(n2062)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_17 (.CI(n28306), .I0(n2009), 
            .I1(VCC_net), .CO(n28307));
    SB_LUT4 encoder0_position_23__I_0_add_1361_16_lut (.I0(GND_net), .I1(n2010), 
            .I2(VCC_net), .I3(n28305), .O(n2063)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_16 (.CI(n28305), .I0(n2010), 
            .I1(VCC_net), .CO(n28306));
    SB_LUT4 i19647_2_lut_3_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n619), .I3(n15_adj_4867), .O(n24425));   // verilog/TinyFPGA_B.v(251[7:11])
    defparam i19647_2_lut_3_lut_4_lut.LUT_INIT = 16'hffbf;
    SB_LUT4 encoder0_position_23__I_0_add_1361_15_lut (.I0(GND_net), .I1(n2011), 
            .I2(VCC_net), .I3(n28304), .O(n2064)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_15 (.CI(n28304), .I0(n2011), 
            .I1(VCC_net), .CO(n28305));
    SB_LUT4 encoder0_position_23__I_0_add_1361_14_lut (.I0(GND_net), .I1(n2012), 
            .I2(VCC_net), .I3(n28303), .O(n2065)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_14 (.CI(n28303), .I0(n2012), 
            .I1(VCC_net), .CO(n28304));
    SB_LUT4 encoder0_position_23__I_0_add_1361_13_lut (.I0(GND_net), .I1(n2013), 
            .I2(VCC_net), .I3(n28302), .O(n2066)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_13 (.CI(n28302), .I0(n2013), 
            .I1(VCC_net), .CO(n28303));
    SB_LUT4 encoder0_position_23__I_0_add_1361_12_lut (.I0(GND_net), .I1(n2014), 
            .I2(VCC_net), .I3(n28301), .O(n2067)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_12 (.CI(n28301), .I0(n2014), 
            .I1(VCC_net), .CO(n28302));
    SB_LUT4 encoder0_position_23__I_0_add_1361_11_lut (.I0(GND_net), .I1(n2015), 
            .I2(VCC_net), .I3(n28300), .O(n2068)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_11 (.CI(n28300), .I0(n2015), 
            .I1(VCC_net), .CO(n28301));
    SB_LUT4 encoder0_position_23__I_0_add_1361_10_lut (.I0(GND_net), .I1(n2016), 
            .I2(VCC_net), .I3(n28299), .O(n2069)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_10 (.CI(n28299), .I0(n2016), 
            .I1(VCC_net), .CO(n28300));
    SB_LUT4 encoder0_position_23__I_0_add_1361_9_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n28298), .O(n2070)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_9 (.CI(n28298), .I0(n2017), 
            .I1(VCC_net), .CO(n28299));
    SB_LUT4 encoder0_position_23__I_0_add_1361_8_lut (.I0(GND_net), .I1(n2018), 
            .I2(GND_net), .I3(n28297), .O(n2071)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_8 (.CI(n28297), .I0(n2018), 
            .I1(GND_net), .CO(n28298));
    SB_LUT4 encoder0_position_23__I_0_add_1361_7_lut (.I0(n2073), .I1(n2019), 
            .I2(GND_net), .I3(n28296), .O(n35924)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_23__I_0_add_1361_7 (.CI(n28296), .I0(n2019), 
            .I1(GND_net), .CO(n28297));
    SB_LUT4 i14038_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n32397), 
            .I3(GND_net), .O(n18827));   // verilog/coms.v(127[12] 300[6])
    defparam i14038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14039_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n32397), 
            .I3(GND_net), .O(n18828));   // verilog/coms.v(127[12] 300[6])
    defparam i14039_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_6_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n28295), .O(n2073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_6 (.CI(n28295), .I0(n2020), 
            .I1(VCC_net), .CO(n28296));
    SB_LUT4 i14040_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n32397), 
            .I3(GND_net), .O(n18829));   // verilog/coms.v(127[12] 300[6])
    defparam i14040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_5_lut (.I0(n6_adj_4920), .I1(n2021), 
            .I2(GND_net), .I3(n28294), .O(n35957)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder0_position_23__I_0_add_1361_5 (.CI(n28294), .I0(n2021), 
            .I1(GND_net), .CO(n28295));
    SB_LUT4 i14041_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n32397), 
            .I3(GND_net), .O(n18830));   // verilog/coms.v(127[12] 300[6])
    defparam i14041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14042_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n32397), 
            .I3(GND_net), .O(n18831));   // verilog/coms.v(127[12] 300[6])
    defparam i14042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14043_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n32397), 
            .I3(GND_net), .O(n18832));   // verilog/coms.v(127[12] 300[6])
    defparam i14043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i463_3_lut (.I0(n675), .I1(n728), 
            .I2(n700), .I3(GND_net), .O(n753));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14044_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n32397), 
            .I3(GND_net), .O(n18833));   // verilog/coms.v(127[12] 300[6])
    defparam i14044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i465_3_lut (.I0(n677), .I1(n730), 
            .I2(n700), .I3(GND_net), .O(n755));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14045_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n32397), 
            .I3(GND_net), .O(n18834));   // verilog/coms.v(127[12] 300[6])
    defparam i14045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_4_lut (.I0(n2076), .I1(n2022), 
            .I2(VCC_net), .I3(n28293), .O(n6_adj_4920)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_23__I_0_add_1361_4 (.CI(n28293), .I0(n2022), 
            .I1(VCC_net), .CO(n28294));
    SB_LUT4 encoder0_position_23__I_0_i467_3_lut (.I0(n679), .I1(n732), 
            .I2(n700), .I3(GND_net), .O(n757));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i466_3_lut (.I0(n678), .I1(n731), 
            .I2(n700), .I3(GND_net), .O(n756));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i464_3_lut (.I0(n676), .I1(n729), 
            .I2(n700), .I3(GND_net), .O(n754));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1361_3_lut (.I0(GND_net), .I1(n775), 
            .I2(GND_net), .I3(n28292), .O(n2076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_660_9_lut (.I0(duty[7]), .I1(n37310), .I2(n18_adj_4872), 
            .I3(n27734), .O(pwm_setpoint_22__N_11[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_1361_3 (.CI(n28292), .I0(n775), 
            .I1(GND_net), .CO(n28293));
    SB_LUT4 i30893_2_lut_3_lut (.I0(n3_adj_4917), .I1(n4_adj_4962), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n619_adj_4960));
    defparam i30893_2_lut_3_lut.LUT_INIT = 16'h7f7f;
    SB_CARRY add_660_9 (.CI(n27734), .I0(n37310), .I1(n18_adj_4872), .CO(n27735));
    SB_CARRY encoder0_position_23__I_0_add_1361_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n28292));
    SB_LUT4 add_1877_23_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n28291), .O(n5805)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n27665), .O(n587)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3933_2_lut (.I0(n2), .I1(encoder0_position[23]), .I2(GND_net), 
            .I3(GND_net), .O(n509));
    defparam i3933_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26735_4_lut (.I0(encoder0_position[22]), .I1(n35954), .I2(encoder0_position[23]), 
            .I3(n3_adj_4917), .O(n675));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26735_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 add_1877_22_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n28290), .O(n5806)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26752_3_lut (.I0(encoder0_position[21]), .I1(n33134), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n676));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14054_3_lut (.I0(\data_in_frame[3] [7]), .I1(rx_data[7]), .I2(n32394), 
            .I3(GND_net), .O(n18843));   // verilog/coms.v(127[12] 300[6])
    defparam i14054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26751_3_lut_4_lut (.I0(n3_adj_4917), .I1(n4_adj_4962), .I2(n5629), 
            .I3(n4_adj_4916), .O(n33134));
    defparam i26751_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 add_28_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n27664), .O(n588)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3291_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4913), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n598_adj_4959));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14055_3_lut (.I0(\data_in_frame[3] [6]), .I1(rx_data[6]), .I2(n32394), 
            .I3(GND_net), .O(n18844));   // verilog/coms.v(127[12] 300[6])
    defparam i14055_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1877_22 (.CI(n28290), .I0(GND_net), .I1(VCC_net), .CO(n28291));
    SB_LUT4 i26743_3_lut_4_lut (.I0(n3_adj_4917), .I1(n4_adj_4962), .I2(n5632), 
            .I3(n7_adj_4913), .O(n33126));
    defparam i26743_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 add_1877_21_lut (.I0(encoder0_position[23]), .I1(GND_net), .I2(n619_adj_4960), 
            .I3(n28289), .O(encoder0_position_scaled_23__N_34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1877_21 (.CI(n28289), .I0(GND_net), .I1(n619_adj_4960), 
            .CO(n28290));
    SB_LUT4 add_660_8_lut (.I0(duty[6]), .I1(n37310), .I2(n19), .I3(n27733), 
            .O(pwm_setpoint_22__N_11[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i26736_3_lut_4_lut (.I0(n3_adj_4917), .I1(n4_adj_4962), .I2(n5631), 
            .I3(n6_adj_4914), .O(n33118));
    defparam i26736_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY add_28_32 (.CI(n27664), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n27665));
    SB_CARRY add_660_8 (.CI(n27733), .I0(n37310), .I1(n19), .CO(n27734));
    SB_LUT4 add_660_7_lut (.I0(duty[5]), .I1(n37310), .I2(n20_adj_4873), 
            .I3(n27732), .O(pwm_setpoint_22__N_11[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14056_3_lut (.I0(\data_in_frame[3] [5]), .I1(rx_data[5]), .I2(n32394), 
            .I3(GND_net), .O(n18845));   // verilog/coms.v(127[12] 300[6])
    defparam i14056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26732_3_lut_4_lut (.I0(n3_adj_4917), .I1(n4_adj_4962), .I2(n5630), 
            .I3(n5_adj_4915), .O(n33114));
    defparam i26732_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_adj_1704 (.I0(n598_adj_4959), .I1(n6_adj_4914), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4894));
    defparam i1_2_lut_adj_1704.LUT_INIT = 16'heeee;
    SB_LUT4 add_1877_20_lut (.I0(GND_net), .I1(GND_net), .I2(n700), .I3(n28288), 
            .O(n5808)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14057_3_lut (.I0(\data_in_frame[3] [4]), .I1(rx_data[4]), .I2(n32394), 
            .I3(GND_net), .O(n18846));   // verilog/coms.v(127[12] 300[6])
    defparam i14057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1831_7_lut (.I0(GND_net), .I1(n509), .I2(GND_net), .I3(n27905), 
            .O(n5627)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1831_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1831_6_lut (.I0(n34993), .I1(n510), .I2(GND_net), .I3(n27904), 
            .O(n35954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1831_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_660_7 (.CI(n27732), .I0(n37310), .I1(n20_adj_4873), .CO(n27733));
    SB_CARRY add_1877_20 (.CI(n28288), .I0(GND_net), .I1(n700), .CO(n28289));
    SB_LUT4 add_660_6_lut (.I0(duty[4]), .I1(n37310), .I2(n21), .I3(n27731), 
            .O(pwm_setpoint_22__N_11[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1877_19_lut (.I0(GND_net), .I1(GND_net), .I2(n778), .I3(n28287), 
            .O(n5809)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_19 (.CI(n28287), .I0(GND_net), .I1(n778), .CO(n28288));
    SB_LUT4 add_28_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n27663), .O(n589)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_660_6 (.CI(n27731), .I0(n37310), .I1(n21), .CO(n27732));
    SB_LUT4 add_1877_18_lut (.I0(GND_net), .I1(GND_net), .I2(n856), .I3(n28286), 
            .O(n5810)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_18 (.CI(n28286), .I0(GND_net), .I1(n856), .CO(n28287));
    SB_LUT4 i14058_3_lut (.I0(\data_in_frame[3] [3]), .I1(rx_data[3]), .I2(n32394), 
            .I3(GND_net), .O(n18847));   // verilog/coms.v(127[12] 300[6])
    defparam i14058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1877_17_lut (.I0(GND_net), .I1(GND_net), .I2(n934), .I3(n28285), 
            .O(n5811)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14059_3_lut (.I0(\data_in_frame[3] [2]), .I1(rx_data[2]), .I2(n32394), 
            .I3(GND_net), .O(n18848));   // verilog/coms.v(127[12] 300[6])
    defparam i14059_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_28_31 (.CI(n27663), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n27664));
    SB_CARRY add_1877_17 (.CI(n28285), .I0(GND_net), .I1(n934), .CO(n28286));
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n4_adj_4916), .I1(n2), .I2(n5_adj_4915), 
            .I3(n7_adj_4894), .O(n4_adj_4962));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'hc888;
    SB_LUT4 add_1877_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1012), .I3(n28284), 
            .O(n5812)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_16 (.CI(n28284), .I0(GND_net), .I1(n1012), .CO(n28285));
    SB_LUT4 add_1877_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1090), .I3(n28283), 
            .O(n5813)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14060_3_lut (.I0(\data_in_frame[3] [1]), .I1(rx_data[1]), .I2(n32394), 
            .I3(GND_net), .O(n18849));   // verilog/coms.v(127[12] 300[6])
    defparam i14060_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1877_15 (.CI(n28283), .I0(GND_net), .I1(n1090), .CO(n28284));
    SB_CARRY add_1831_6 (.CI(n27904), .I0(n510), .I1(GND_net), .CO(n27905));
    SB_LUT4 add_1877_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1168), .I3(n28282), 
            .O(n5814)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n27643), .O(n609)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_14 (.CI(n28282), .I0(GND_net), .I1(n1168), .CO(n28283));
    SB_LUT4 add_1831_5_lut (.I0(GND_net), .I1(n511), .I2(VCC_net), .I3(n27903), 
            .O(n5629)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1831_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1877_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1246), .I3(n28281), 
            .O(n5815)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_13 (.CI(n28281), .I0(GND_net), .I1(n1246), .CO(n28282));
    SB_LUT4 add_660_5_lut (.I0(duty[3]), .I1(n37310), .I2(n22), .I3(n27730), 
            .O(pwm_setpoint_22__N_11[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1877_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1324), .I3(n28280), 
            .O(n5816)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_12 (.CI(n28280), .I0(GND_net), .I1(n1324), .CO(n28281));
    SB_LUT4 add_1877_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1402), .I3(n28279), 
            .O(n5817)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n27987), .I0(encoder1_position[12]), 
            .I1(n13_adj_4946), .CO(n27988));
    SB_CARRY add_1877_11 (.CI(n28279), .I0(GND_net), .I1(n1402), .CO(n28280));
    SB_LUT4 add_1877_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1480), .I3(n28278), 
            .O(n5818)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_10 (.CI(n28278), .I0(GND_net), .I1(n1480), .CO(n28279));
    SB_LUT4 add_1877_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1558), .I3(n28277), 
            .O(n5819)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_9 (.CI(n28277), .I0(GND_net), .I1(n1558), .CO(n28278));
    SB_CARRY add_1831_5 (.CI(n27903), .I0(n511), .I1(VCC_net), .CO(n27904));
    SB_LUT4 add_1877_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1636), .I3(n28276), 
            .O(n5820)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n27636), .O(n616)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1831_4_lut (.I0(GND_net), .I1(n425), .I2(GND_net), .I3(n27902), 
            .O(n5630)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1831_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_8 (.CI(n28276), .I0(GND_net), .I1(n1636), .CO(n28277));
    SB_CARRY add_1831_4 (.CI(n27902), .I0(n425), .I1(GND_net), .CO(n27903));
    SB_LUT4 add_1877_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1714), .I3(n28275), 
            .O(n5821)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_7 (.CI(n28275), .I0(GND_net), .I1(n1714), .CO(n28276));
    SB_LUT4 add_1877_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1792), .I3(n28274), 
            .O(n5822)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4947), .I3(n27986), .O(displacement_23__N_58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_6 (.CI(n28274), .I0(GND_net), .I1(n1792), .CO(n28275));
    SB_LUT4 add_1877_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1870), .I3(n28273), 
            .O(n5823)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_5 (.CI(n28273), .I0(GND_net), .I1(n1870), .CO(n28274));
    SB_LUT4 add_1877_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1948), .I3(n28272), 
            .O(n5824)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_4 (.CI(n28272), .I0(GND_net), .I1(n1948), .CO(n28273));
    SB_CARRY add_660_5 (.CI(n27730), .I0(n37310), .I1(n22), .CO(n27731));
    SB_LUT4 add_1877_3_lut (.I0(GND_net), .I1(GND_net), .I2(n2026), .I3(n28271), 
            .O(n5825)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1831_3_lut (.I0(GND_net), .I1(n513), .I2(VCC_net), .I3(n27901), 
            .O(n5631)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1831_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n27662), .O(n590)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n27986), .I0(encoder1_position[11]), 
            .I1(n14_adj_4947), .CO(n27987));
    SB_CARRY add_1877_3 (.CI(n28271), .I0(GND_net), .I1(n2026), .CO(n28272));
    SB_LUT4 add_660_4_lut (.I0(duty[2]), .I1(n37310), .I2(n23), .I3(n27729), 
            .O(pwm_setpoint_22__N_11[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4948), .I3(n27985), .O(displacement_23__N_58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n27985), .I0(encoder1_position[10]), 
            .I1(n15_adj_4948), .CO(n27986));
    SB_LUT4 add_1877_2_lut (.I0(GND_net), .I1(GND_net), .I2(n24674), .I3(VCC_net), 
            .O(n5826)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1877_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1877_2 (.CI(VCC_net), .I0(GND_net), .I1(n24674), .CO(n28271));
    SB_LUT4 encoder0_position_23__I_0_add_1308_24_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n28270), .O(n1975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1308_23_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n28269), .O(n1976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4949), .I3(n27984), .O(displacement_23__N_58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_23 (.CI(n28269), .I0(n1923), 
            .I1(VCC_net), .CO(n28270));
    SB_CARRY add_1831_3 (.CI(n27901), .I0(n513), .I1(VCC_net), .CO(n27902));
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n27984), .I0(encoder1_position[9]), 
            .I1(n16_adj_4949), .CO(n27985));
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4950), .I3(n27983), .O(displacement_23__N_58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n27983), .I0(encoder1_position[8]), 
            .I1(n17_adj_4950), .CO(n27984));
    SB_LUT4 encoder0_position_23__I_0_add_1308_22_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n28268), .O(n1977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_660_4 (.CI(n27729), .I0(n37310), .I1(n23), .CO(n27730));
    SB_CARRY encoder0_position_23__I_0_add_1308_22 (.CI(n28268), .I0(n1924), 
            .I1(VCC_net), .CO(n28269));
    SB_LUT4 add_1831_2_lut (.I0(GND_net), .I1(n598_adj_4959), .I2(GND_net), 
            .I3(VCC_net), .O(n5632)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1831_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1831_2 (.CI(VCC_net), .I0(n598_adj_4959), .I1(GND_net), 
            .CO(n27901));
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4951), .I3(n27982), .O(displacement_23__N_58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_11 (.CI(n27643), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n27644));
    SB_LUT4 encoder0_position_23__I_0_add_1308_21_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n28267), .O(n1978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_21 (.CI(n28267), .I0(n1925), 
            .I1(VCC_net), .CO(n28268));
    SB_LUT4 encoder0_position_23__I_0_add_1308_20_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n28266), .O(n1979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_20 (.CI(n28266), .I0(n1926), 
            .I1(VCC_net), .CO(n28267));
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n27982), .I0(encoder1_position[7]), 
            .I1(n18_adj_4951), .CO(n27983));
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4952), .I3(n27981), .O(displacement_23__N_58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_30 (.CI(n27662), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n27663));
    SB_LUT4 encoder0_position_23__I_0_add_1308_19_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n28265), .O(n1980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_19 (.CI(n28265), .I0(n1927), 
            .I1(VCC_net), .CO(n28266));
    SB_LUT4 add_660_3_lut (.I0(duty[1]), .I1(n37310), .I2(n24), .I3(n27728), 
            .O(pwm_setpoint_22__N_11[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_1308_18_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n28264), .O(n1981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_18 (.CI(n28264), .I0(n1928), 
            .I1(VCC_net), .CO(n28265));
    SB_LUT4 i14061_3_lut (.I0(\data_in_frame[3] [0]), .I1(rx_data[0]), .I2(n32394), 
            .I3(GND_net), .O(n18850));   // verilog/coms.v(127[12] 300[6])
    defparam i14061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_17_lut (.I0(GND_net), .I1(n1929), 
            .I2(VCC_net), .I3(n28263), .O(n1982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n27981), .I0(encoder1_position[6]), 
            .I1(n19_adj_4952), .CO(n27982));
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4953), .I3(n27980), .O(displacement_23__N_58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n27980), .I0(encoder1_position[5]), 
            .I1(n20_adj_4953), .CO(n27981));
    SB_CARRY encoder0_position_23__I_0_add_1308_17 (.CI(n28263), .I0(n1929), 
            .I1(VCC_net), .CO(n28264));
    SB_LUT4 encoder0_position_23__I_0_i409_3_lut_4_lut (.I0(n2), .I1(encoder0_position[23]), 
            .I2(n619_adj_4960), .I3(n5627), .O(n674));
    defparam encoder0_position_23__I_0_i409_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_LUT4 encoder0_position_23__I_0_add_1308_16_lut (.I0(GND_net), .I1(n1930), 
            .I2(VCC_net), .I3(n28262), .O(n1983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_16 (.CI(n28262), .I0(n1930), 
            .I1(VCC_net), .CO(n28263));
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4954), .I3(n27979), .O(displacement_23__N_58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1706 (.I0(n4452), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n66), .I3(GND_net), .O(n1));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1706.LUT_INIT = 16'h0404;
    SB_LUT4 encoder0_position_23__I_0_add_1308_15_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n28261), .O(n1984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_15 (.CI(n28261), .I0(n1931), 
            .I1(VCC_net), .CO(n28262));
    SB_LUT4 encoder0_position_23__I_0_add_1308_14_lut (.I0(GND_net), .I1(n1932), 
            .I2(VCC_net), .I3(n28260), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n27979), .I0(encoder1_position[4]), 
            .I1(n21_adj_4954), .CO(n27980));
    SB_CARRY encoder0_position_23__I_0_add_1308_14 (.CI(n28260), .I0(n1932), 
            .I1(VCC_net), .CO(n28261));
    SB_LUT4 encoder0_position_23__I_0_add_1308_13_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n28259), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_13 (.CI(n28259), .I0(n1933), 
            .I1(VCC_net), .CO(n28260));
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4955), .I3(n27978), .O(displacement_23__N_58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n27978), .I0(encoder1_position[3]), 
            .I1(n22_adj_4955), .CO(n27979));
    SB_LUT4 encoder0_position_23__I_0_add_1308_12_lut (.I0(GND_net), .I1(n1934), 
            .I2(VCC_net), .I3(n28258), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_12 (.CI(n28258), .I0(n1934), 
            .I1(VCC_net), .CO(n28259));
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4956), .I3(n27977), .O(displacement_23__N_58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n27977), .I0(encoder1_position[2]), 
            .I1(n23_adj_4956), .CO(n27978));
    SB_LUT4 encoder0_position_23__I_0_add_1308_11_lut (.I0(GND_net), .I1(n1935), 
            .I2(VCC_net), .I3(n28257), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_660_3 (.CI(n27728), .I0(n37310), .I1(n24), .CO(n27729));
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4957), .I3(n27976), .O(displacement_23__N_58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_11 (.CI(n28257), .I0(n1935), 
            .I1(VCC_net), .CO(n28258));
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n27976), .I0(encoder1_position[1]), 
            .I1(n24_adj_4957), .CO(n27977));
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4958), .I3(VCC_net), .O(displacement_23__N_58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_4 (.CI(n27636), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n27637));
    SB_LUT4 add_660_2_lut (.I0(duty[0]), .I1(n37310), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_11[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_660_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4958), .CO(n27976));
    SB_LUT4 add_28_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n27642), .O(n610)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1308_10_lut (.I0(GND_net), .I1(n1936), 
            .I2(VCC_net), .I3(n28256), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_10 (.CI(n28256), .I0(n1936), 
            .I1(VCC_net), .CO(n28257));
    SB_CARRY add_660_2 (.CI(VCC_net), .I0(n37310), .I1(n25), .CO(n27728));
    SB_LUT4 add_28_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n27661), .O(n591)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_10 (.CI(n27642), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n27643));
    SB_CARRY add_28_29 (.CI(n27661), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n27662));
    SB_LUT4 add_28_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n27660), .O(n592)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1308_9_lut (.I0(GND_net), .I1(n1937), 
            .I2(VCC_net), .I3(n28255), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_28 (.CI(n27660), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n27661));
    SB_CARRY encoder0_position_23__I_0_add_1308_9 (.CI(n28255), .I0(n1937), 
            .I1(VCC_net), .CO(n28256));
    SB_LUT4 encoder0_position_23__I_0_add_1308_8_lut (.I0(GND_net), .I1(n1938), 
            .I2(VCC_net), .I3(n28254), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_8 (.CI(n28254), .I0(n1938), 
            .I1(VCC_net), .CO(n28255));
    SB_LUT4 encoder0_position_23__I_0_add_1308_7_lut (.I0(GND_net), .I1(n1939), 
            .I2(GND_net), .I3(n28253), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_7 (.CI(n28253), .I0(n1939), 
            .I1(GND_net), .CO(n28254));
    SB_LUT4 encoder0_position_23__I_0_add_1308_6_lut (.I0(GND_net), .I1(n1940), 
            .I2(GND_net), .I3(n28252), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n27659), .O(n593)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_6 (.CI(n28252), .I0(n1940), 
            .I1(GND_net), .CO(n28253));
    SB_LUT4 encoder0_position_23__I_0_add_1308_5_lut (.I0(GND_net), .I1(n1941), 
            .I2(VCC_net), .I3(n28251), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_5 (.CI(n28251), .I0(n1941), 
            .I1(VCC_net), .CO(n28252));
    SB_LUT4 encoder0_position_23__I_0_add_1308_4_lut (.I0(GND_net), .I1(n1942), 
            .I2(GND_net), .I3(n28250), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_4 (.CI(n28250), .I0(n1942), 
            .I1(GND_net), .CO(n28251));
    SB_LUT4 encoder0_position_23__I_0_add_1308_3_lut (.I0(GND_net), .I1(n1943), 
            .I2(VCC_net), .I3(n28249), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5132[0]), .I1(n35900), .I2(n4867), 
            .I3(n10_adj_4926), .O(n8_adj_5030));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_CARRY encoder0_position_23__I_0_add_1308_3 (.CI(n28249), .I0(n1943), 
            .I1(VCC_net), .CO(n28250));
    SB_CARRY add_28_27 (.CI(n27659), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n27660));
    SB_LUT4 encoder0_position_23__I_0_add_1308_2_lut (.I0(GND_net), .I1(n774), 
            .I2(GND_net), .I3(VCC_net), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_2 (.CI(VCC_net), .I0(n774), 
            .I1(GND_net), .CO(n28249));
    SB_LUT4 encoder0_position_23__I_0_add_1255_23_lut (.I0(GND_net), .I1(n1844), 
            .I2(VCC_net), .I3(n28248), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_22_lut (.I0(GND_net), .I1(n1845), 
            .I2(VCC_net), .I3(n28247), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_22 (.CI(n28247), .I0(n1845), 
            .I1(VCC_net), .CO(n28248));
    SB_LUT4 encoder0_position_23__I_0_add_1255_21_lut (.I0(GND_net), .I1(n1846), 
            .I2(VCC_net), .I3(n28246), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_21 (.CI(n28246), .I0(n1846), 
            .I1(VCC_net), .CO(n28247));
    SB_LUT4 add_28_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n27658), .O(n594)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_20_lut (.I0(GND_net), .I1(n1847), 
            .I2(VCC_net), .I3(n28245), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_20 (.CI(n28245), .I0(n1847), 
            .I1(VCC_net), .CO(n28246));
    SB_CARRY add_28_26 (.CI(n27658), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n27659));
    SB_LUT4 encoder0_position_23__I_0_add_1255_19_lut (.I0(GND_net), .I1(n1848), 
            .I2(VCC_net), .I3(n28244), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_19 (.CI(n28244), .I0(n1848), 
            .I1(VCC_net), .CO(n28245));
    SB_LUT4 encoder0_position_23__I_0_add_1255_18_lut (.I0(GND_net), .I1(n1849), 
            .I2(VCC_net), .I3(n28243), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_18 (.CI(n28243), .I0(n1849), 
            .I1(VCC_net), .CO(n28244));
    SB_LUT4 encoder0_position_23__I_0_add_1255_17_lut (.I0(GND_net), .I1(n1850), 
            .I2(VCC_net), .I3(n28242), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_17 (.CI(n28242), .I0(n1850), 
            .I1(VCC_net), .CO(n28243));
    SB_LUT4 encoder0_position_23__I_0_add_1255_16_lut (.I0(GND_net), .I1(n1851), 
            .I2(VCC_net), .I3(n28241), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_16 (.CI(n28241), .I0(n1851), 
            .I1(VCC_net), .CO(n28242));
    SB_LUT4 encoder0_position_23__I_0_add_1255_15_lut (.I0(GND_net), .I1(n1852), 
            .I2(VCC_net), .I3(n28240), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n27657), .O(n595)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14070_3_lut (.I0(\data_in_frame[1] [7]), .I1(rx_data[7]), .I2(n32395), 
            .I3(GND_net), .O(n18859));   // verilog/coms.v(127[12] 300[6])
    defparam i14070_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14071_3_lut (.I0(\data_in_frame[1] [6]), .I1(rx_data[6]), .I2(n32395), 
            .I3(GND_net), .O(n18860));   // verilog/coms.v(127[12] 300[6])
    defparam i14071_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14072_3_lut (.I0(\data_in_frame[1] [5]), .I1(rx_data[5]), .I2(n32395), 
            .I3(GND_net), .O(n18861));   // verilog/coms.v(127[12] 300[6])
    defparam i14072_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1255_15 (.CI(n28240), .I0(n1852), 
            .I1(VCC_net), .CO(n28241));
    SB_LUT4 encoder0_position_23__I_0_add_1255_14_lut (.I0(GND_net), .I1(n1853), 
            .I2(VCC_net), .I3(n28239), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_14 (.CI(n28239), .I0(n1853), 
            .I1(VCC_net), .CO(n28240));
    SB_LUT4 encoder0_position_23__I_0_add_1255_13_lut (.I0(GND_net), .I1(n1854), 
            .I2(VCC_net), .I3(n28238), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_13 (.CI(n28238), .I0(n1854), 
            .I1(VCC_net), .CO(n28239));
    SB_LUT4 encoder0_position_23__I_0_add_1255_12_lut (.I0(GND_net), .I1(n1855), 
            .I2(VCC_net), .I3(n28237), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_12 (.CI(n28237), .I0(n1855), 
            .I1(VCC_net), .CO(n28238));
    SB_LUT4 encoder0_position_23__I_0_add_1255_11_lut (.I0(GND_net), .I1(n1856), 
            .I2(VCC_net), .I3(n28236), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_11 (.CI(n28236), .I0(n1856), 
            .I1(VCC_net), .CO(n28237));
    SB_LUT4 encoder0_position_23__I_0_add_1255_10_lut (.I0(GND_net), .I1(n1857), 
            .I2(VCC_net), .I3(n28235), .O(n1910)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_10 (.CI(n28235), .I0(n1857), 
            .I1(VCC_net), .CO(n28236));
    SB_LUT4 encoder0_position_23__I_0_add_1255_9_lut (.I0(GND_net), .I1(n1858), 
            .I2(VCC_net), .I3(n28234), .O(n1911)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n27635), .O(n617)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_9 (.CI(n28234), .I0(n1858), 
            .I1(VCC_net), .CO(n28235));
    SB_LUT4 encoder0_position_23__I_0_add_1255_8_lut (.I0(GND_net), .I1(n1859), 
            .I2(VCC_net), .I3(n28233), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_8 (.CI(n28233), .I0(n1859), 
            .I1(VCC_net), .CO(n28234));
    SB_LUT4 encoder0_position_23__I_0_add_1255_7_lut (.I0(GND_net), .I1(n1860), 
            .I2(GND_net), .I3(n28232), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_7 (.CI(n28232), .I0(n1860), 
            .I1(GND_net), .CO(n28233));
    SB_LUT4 encoder0_position_23__I_0_add_1255_6_lut (.I0(GND_net), .I1(n1861), 
            .I2(GND_net), .I3(n28231), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_25 (.CI(n27657), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n27658));
    SB_LUT4 add_28_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n27641), .O(n611)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_6 (.CI(n28231), .I0(n1861), 
            .I1(GND_net), .CO(n28232));
    SB_LUT4 encoder0_position_23__I_0_add_1255_5_lut (.I0(GND_net), .I1(n1862), 
            .I2(VCC_net), .I3(n28230), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_5 (.CI(n28230), .I0(n1862), 
            .I1(VCC_net), .CO(n28231));
    SB_CARRY add_28_9 (.CI(n27641), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n27642));
    SB_LUT4 encoder0_position_23__I_0_add_1255_4_lut (.I0(GND_net), .I1(n1863), 
            .I2(GND_net), .I3(n28229), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_4 (.CI(n28229), .I0(n1863), 
            .I1(GND_net), .CO(n28230));
    SB_LUT4 add_28_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n27656), .O(n596)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_3_lut (.I0(GND_net), .I1(n1864), 
            .I2(VCC_net), .I3(n28228), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_24 (.CI(n27656), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n27657));
    SB_CARRY encoder0_position_23__I_0_add_1255_3 (.CI(n28228), .I0(n1864), 
            .I1(VCC_net), .CO(n28229));
    SB_LUT4 add_28_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n27655), .O(n597)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_23 (.CI(n27655), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n27656));
    SB_LUT4 encoder0_position_23__I_0_add_1255_2_lut (.I0(GND_net), .I1(n773), 
            .I2(GND_net), .I3(VCC_net), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14073_3_lut (.I0(\data_in_frame[1] [4]), .I1(rx_data[4]), .I2(n32395), 
            .I3(GND_net), .O(n18862));   // verilog/coms.v(127[12] 300[6])
    defparam i14073_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14074_3_lut (.I0(\data_in_frame[1] [3]), .I1(rx_data[3]), .I2(n32395), 
            .I3(GND_net), .O(n18863));   // verilog/coms.v(127[12] 300[6])
    defparam i14074_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14075_3_lut (.I0(\data_in_frame[1] [2]), .I1(rx_data[2]), .I2(n32395), 
            .I3(GND_net), .O(n18864));   // verilog/coms.v(127[12] 300[6])
    defparam i14075_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14076_3_lut (.I0(\data_in_frame[1] [1]), .I1(rx_data[1]), .I2(n32395), 
            .I3(GND_net), .O(n18865));   // verilog/coms.v(127[12] 300[6])
    defparam i14076_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14077_3_lut (.I0(\data_in_frame[1] [0]), .I1(rx_data[0]), .I2(n32395), 
            .I3(GND_net), .O(n18866));   // verilog/coms.v(127[12] 300[6])
    defparam i14077_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_72_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[19]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i20_3_lut (.I0(encoder0_position_scaled[19]), .I1(motor_state_23__N_82[19]), 
            .I2(n15), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i14085_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n34118), .I3(GND_net), .O(n18874));   // verilog/coms.v(127[12] 300[6])
    defparam i14085_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4956));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14086_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n34118), .I3(GND_net), .O(n18875));   // verilog/coms.v(127[12] 300[6])
    defparam i14086_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4955));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14087_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n34118), .I3(GND_net), .O(n18876));   // verilog/coms.v(127[12] 300[6])
    defparam i14087_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4954));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_28_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n27654), .O(n598)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_2 (.CI(VCC_net), .I0(n773), 
            .I1(GND_net), .CO(n28228));
    SB_LUT4 encoder0_position_23__I_0_add_1202_22_lut (.I0(GND_net), .I1(n1766), 
            .I2(VCC_net), .I3(n28227), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_72_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[20]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_add_1202_21_lut (.I0(GND_net), .I1(n1767), 
            .I2(VCC_net), .I3(n28226), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_21 (.CI(n28226), .I0(n1767), 
            .I1(VCC_net), .CO(n28227));
    SB_LUT4 mux_70_i21_3_lut (.I0(encoder0_position_scaled[20]), .I1(motor_state_23__N_82[20]), 
            .I2(n15), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 encoder0_position_23__I_0_add_1202_20_lut (.I0(GND_net), .I1(n1768), 
            .I2(VCC_net), .I3(n28225), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_20 (.CI(n28225), .I0(n1768), 
            .I1(VCC_net), .CO(n28226));
    SB_LUT4 encoder0_position_23__I_0_add_1202_19_lut (.I0(GND_net), .I1(n1769), 
            .I2(VCC_net), .I3(n28224), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_19_lut.LUT_INIT = 16'hC33C;
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n18651));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4953));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14088_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n34118), .I3(GND_net), .O(n18877));   // verilog/coms.v(127[12] 300[6])
    defparam i14088_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_72_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[21]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14089_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n34118), .I3(GND_net), .O(n18878));   // verilog/coms.v(127[12] 300[6])
    defparam i14089_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i22_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_82[21]), 
            .I2(n15), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i22_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_23__I_0_add_1202_19 (.CI(n28224), .I0(n1769), 
            .I1(VCC_net), .CO(n28225));
    SB_LUT4 encoder0_position_23__I_0_add_1202_18_lut (.I0(GND_net), .I1(n1770), 
            .I2(VCC_net), .I3(n28223), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_18 (.CI(n28223), .I0(n1770), 
            .I1(VCC_net), .CO(n28224));
    SB_LUT4 encoder0_position_23__I_0_add_1202_17_lut (.I0(GND_net), .I1(n1771), 
            .I2(VCC_net), .I3(n28222), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_17 (.CI(n28222), .I0(n1771), 
            .I1(VCC_net), .CO(n28223));
    SB_LUT4 encoder0_position_23__I_0_add_1202_16_lut (.I0(GND_net), .I1(n1772), 
            .I2(VCC_net), .I3(n28221), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_16 (.CI(n28221), .I0(n1772), 
            .I1(VCC_net), .CO(n28222));
    SB_LUT4 encoder0_position_23__I_0_add_1202_15_lut (.I0(GND_net), .I1(n1773), 
            .I2(VCC_net), .I3(n28220), .O(n1826)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_15 (.CI(n28220), .I0(n1773), 
            .I1(VCC_net), .CO(n28221));
    SB_LUT4 encoder0_position_23__I_0_add_1202_14_lut (.I0(GND_net), .I1(n1774), 
            .I2(VCC_net), .I3(n28219), .O(n1827)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_14 (.CI(n28219), .I0(n1774), 
            .I1(VCC_net), .CO(n28220));
    SB_LUT4 encoder0_position_23__I_0_add_1202_13_lut (.I0(GND_net), .I1(n1775), 
            .I2(VCC_net), .I3(n28218), .O(n1828)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_13 (.CI(n28218), .I0(n1775), 
            .I1(VCC_net), .CO(n28219));
    SB_LUT4 encoder0_position_23__I_0_add_1202_12_lut (.I0(GND_net), .I1(n1776), 
            .I2(VCC_net), .I3(n28217), .O(n1829)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_12 (.CI(n28217), .I0(n1776), 
            .I1(VCC_net), .CO(n28218));
    SB_LUT4 encoder0_position_23__I_0_add_1202_11_lut (.I0(GND_net), .I1(n1777), 
            .I2(VCC_net), .I3(n28216), .O(n1830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_11 (.CI(n28216), .I0(n1777), 
            .I1(VCC_net), .CO(n28217));
    SB_LUT4 encoder0_position_23__I_0_add_1202_10_lut (.I0(GND_net), .I1(n1778), 
            .I2(VCC_net), .I3(n28215), .O(n1831)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_10 (.CI(n28215), .I0(n1778), 
            .I1(VCC_net), .CO(n28216));
    SB_LUT4 encoder0_position_23__I_0_add_1202_9_lut (.I0(GND_net), .I1(n1779), 
            .I2(VCC_net), .I3(n28214), .O(n1832)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_9 (.CI(n28214), .I0(n1779), 
            .I1(VCC_net), .CO(n28215));
    SB_LUT4 encoder0_position_23__I_0_add_1202_8_lut (.I0(GND_net), .I1(n1780), 
            .I2(VCC_net), .I3(n28213), .O(n1833)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_8 (.CI(n28213), .I0(n1780), 
            .I1(VCC_net), .CO(n28214));
    SB_LUT4 encoder0_position_23__I_0_add_1202_7_lut (.I0(GND_net), .I1(n1781), 
            .I2(GND_net), .I3(n28212), .O(n1834)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_7 (.CI(n28212), .I0(n1781), 
            .I1(GND_net), .CO(n28213));
    SB_CARRY add_28_22 (.CI(n27654), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n27655));
    SB_LUT4 encoder0_position_23__I_0_add_1202_6_lut (.I0(GND_net), .I1(n1782), 
            .I2(GND_net), .I3(n28211), .O(n1835)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n27653), .O(n599)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_6 (.CI(n28211), .I0(n1782), 
            .I1(GND_net), .CO(n28212));
    SB_LUT4 encoder0_position_23__I_0_add_1202_5_lut (.I0(GND_net), .I1(n1783), 
            .I2(VCC_net), .I3(n28210), .O(n1836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_5 (.CI(n28210), .I0(n1783), 
            .I1(VCC_net), .CO(n28211));
    SB_LUT4 encoder0_position_23__I_0_add_1202_4_lut (.I0(GND_net), .I1(n1784), 
            .I2(GND_net), .I3(n28209), .O(n1837)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_4 (.CI(n28209), .I0(n1784), 
            .I1(GND_net), .CO(n28210));
    SB_LUT4 encoder0_position_23__I_0_add_1202_3_lut (.I0(GND_net), .I1(n1785), 
            .I2(VCC_net), .I3(n28208), .O(n1838)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_3 (.CI(n28208), .I0(n1785), 
            .I1(VCC_net), .CO(n28209));
    SB_LUT4 encoder0_position_23__I_0_add_1202_2_lut (.I0(GND_net), .I1(n772), 
            .I2(GND_net), .I3(VCC_net), .O(n1839)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_2 (.CI(VCC_net), .I0(n772), 
            .I1(GND_net), .CO(n28208));
    SB_LUT4 encoder0_position_23__I_0_add_1149_21_lut (.I0(GND_net), .I1(n1688), 
            .I2(VCC_net), .I3(n28207), .O(n1741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1149_20_lut (.I0(GND_net), .I1(n1689), 
            .I2(VCC_net), .I3(n28206), .O(n1742)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_20 (.CI(n28206), .I0(n1689), 
            .I1(VCC_net), .CO(n28207));
    SB_LUT4 encoder0_position_23__I_0_add_1149_19_lut (.I0(GND_net), .I1(n1690), 
            .I2(VCC_net), .I3(n28205), .O(n1743)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_19 (.CI(n28205), .I0(n1690), 
            .I1(VCC_net), .CO(n28206));
    SB_LUT4 encoder0_position_23__I_0_add_1149_18_lut (.I0(GND_net), .I1(n1691), 
            .I2(VCC_net), .I3(n28204), .O(n1744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_18 (.CI(n28204), .I0(n1691), 
            .I1(VCC_net), .CO(n28205));
    SB_LUT4 encoder0_position_23__I_0_add_1149_17_lut (.I0(GND_net), .I1(n1692), 
            .I2(VCC_net), .I3(n28203), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_17 (.CI(n28203), .I0(n1692), 
            .I1(VCC_net), .CO(n28204));
    SB_LUT4 encoder0_position_23__I_0_add_1149_16_lut (.I0(GND_net), .I1(n1693), 
            .I2(VCC_net), .I3(n28202), .O(n1746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_16 (.CI(n28202), .I0(n1693), 
            .I1(VCC_net), .CO(n28203));
    SB_LUT4 encoder0_position_23__I_0_add_1149_15_lut (.I0(GND_net), .I1(n1694), 
            .I2(VCC_net), .I3(n28201), .O(n1747)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_15 (.CI(n28201), .I0(n1694), 
            .I1(VCC_net), .CO(n28202));
    SB_LUT4 i14090_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n34118), .I3(GND_net), .O(n18879));   // verilog/coms.v(127[12] 300[6])
    defparam i14090_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1149_14_lut (.I0(GND_net), .I1(n1695), 
            .I2(VCC_net), .I3(n28200), .O(n1748)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_14 (.CI(n28200), .I0(n1695), 
            .I1(VCC_net), .CO(n28201));
    SB_LUT4 encoder0_position_23__I_0_add_1149_13_lut (.I0(GND_net), .I1(n1696), 
            .I2(VCC_net), .I3(n28199), .O(n1749)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_13 (.CI(n28199), .I0(n1696), 
            .I1(VCC_net), .CO(n28200));
    SB_LUT4 encoder0_position_23__I_0_add_1149_12_lut (.I0(GND_net), .I1(n1697), 
            .I2(VCC_net), .I3(n28198), .O(n1750)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_12 (.CI(n28198), .I0(n1697), 
            .I1(VCC_net), .CO(n28199));
    SB_LUT4 encoder0_position_23__I_0_add_1149_11_lut (.I0(GND_net), .I1(n1698), 
            .I2(VCC_net), .I3(n28197), .O(n1751)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_11 (.CI(n28197), .I0(n1698), 
            .I1(VCC_net), .CO(n28198));
    SB_LUT4 encoder0_position_23__I_0_add_1149_10_lut (.I0(GND_net), .I1(n1699), 
            .I2(VCC_net), .I3(n28196), .O(n1752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_10 (.CI(n28196), .I0(n1699), 
            .I1(VCC_net), .CO(n28197));
    SB_LUT4 encoder0_position_23__I_0_add_1149_9_lut (.I0(GND_net), .I1(n1700), 
            .I2(VCC_net), .I3(n28195), .O(n1753)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_9 (.CI(n28195), .I0(n1700), 
            .I1(VCC_net), .CO(n28196));
    SB_CARRY add_28_21 (.CI(n27653), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n27654));
    SB_LUT4 encoder0_position_23__I_0_add_1149_8_lut (.I0(GND_net), .I1(n1701), 
            .I2(VCC_net), .I3(n28194), .O(n1754)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_8 (.CI(n28194), .I0(n1701), 
            .I1(VCC_net), .CO(n28195));
    SB_LUT4 encoder0_position_23__I_0_add_1149_7_lut (.I0(GND_net), .I1(n1702), 
            .I2(GND_net), .I3(n28193), .O(n1755)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_7 (.CI(n28193), .I0(n1702), 
            .I1(GND_net), .CO(n28194));
    SB_LUT4 encoder0_position_23__I_0_add_1149_6_lut (.I0(GND_net), .I1(n1703), 
            .I2(GND_net), .I3(n28192), .O(n1756)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_6 (.CI(n28192), .I0(n1703), 
            .I1(GND_net), .CO(n28193));
    SB_LUT4 encoder0_position_23__I_0_add_1149_5_lut (.I0(GND_net), .I1(n1704), 
            .I2(VCC_net), .I3(n28191), .O(n1757)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_5 (.CI(n28191), .I0(n1704), 
            .I1(VCC_net), .CO(n28192));
    SB_LUT4 encoder0_position_23__I_0_add_1149_4_lut (.I0(GND_net), .I1(n1705), 
            .I2(GND_net), .I3(n28190), .O(n1758)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_4 (.CI(n28190), .I0(n1705), 
            .I1(GND_net), .CO(n28191));
    SB_LUT4 encoder0_position_23__I_0_add_1149_3_lut (.I0(GND_net), .I1(n1706), 
            .I2(VCC_net), .I3(n28189), .O(n1759)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_3 (.CI(n28189), .I0(n1706), 
            .I1(VCC_net), .CO(n28190));
    SB_LUT4 encoder0_position_23__I_0_add_1149_2_lut (.I0(GND_net), .I1(n771), 
            .I2(GND_net), .I3(VCC_net), .O(n1760)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_2 (.CI(VCC_net), .I0(n771), 
            .I1(GND_net), .CO(n28189));
    SB_LUT4 add_28_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n27652), .O(n600)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_20_lut (.I0(GND_net), .I1(n1610), 
            .I2(VCC_net), .I3(n28188), .O(n1663)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_19_lut (.I0(GND_net), .I1(n1611), 
            .I2(VCC_net), .I3(n28187), .O(n1664)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14091_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n34118), .I3(GND_net), .O(n18880));   // verilog/coms.v(127[12] 300[6])
    defparam i14091_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4952));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14092_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n34118), .I3(GND_net), .O(n18881));   // verilog/coms.v(127[12] 300[6])
    defparam i14092_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14093_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n34118), .I3(GND_net), .O(n18882));   // verilog/coms.v(127[12] 300[6])
    defparam i14093_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_4_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n5131), .I3(n24425), .O(n31590));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hc700;
    SB_LUT4 i14094_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n34118), .I3(GND_net), .O(n18883));   // verilog/coms.v(127[12] 300[6])
    defparam i14094_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_72_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[22]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i23_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_82[22]), 
            .I2(n15), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i23_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY encoder0_position_23__I_0_add_1096_19 (.CI(n28187), .I0(n1611), 
            .I1(VCC_net), .CO(n28188));
    SB_LUT4 encoder0_position_23__I_0_add_1096_18_lut (.I0(GND_net), .I1(n1612), 
            .I2(VCC_net), .I3(n28186), .O(n1665)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n18163), 
            .D(n618), .R(n18489));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_CARRY encoder0_position_23__I_0_add_1096_18 (.CI(n28186), .I0(n1612), 
            .I1(VCC_net), .CO(n28187));
    SB_LUT4 encoder0_position_23__I_0_add_1096_17_lut (.I0(GND_net), .I1(n1613), 
            .I2(VCC_net), .I3(n28185), .O(n1666)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_17 (.CI(n28185), .I0(n1613), 
            .I1(VCC_net), .CO(n28186));
    SB_LUT4 encoder0_position_23__I_0_add_1096_16_lut (.I0(GND_net), .I1(n1614), 
            .I2(VCC_net), .I3(n28184), .O(n1667)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_16 (.CI(n28184), .I0(n1614), 
            .I1(VCC_net), .CO(n28185));
    SB_LUT4 encoder0_position_23__I_0_add_1096_15_lut (.I0(GND_net), .I1(n1615), 
            .I2(VCC_net), .I3(n28183), .O(n1668)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_15 (.CI(n28183), .I0(n1615), 
            .I1(VCC_net), .CO(n28184));
    SB_LUT4 encoder0_position_23__I_0_add_1096_14_lut (.I0(GND_net), .I1(n1616), 
            .I2(VCC_net), .I3(n28182), .O(n1669)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_14 (.CI(n28182), .I0(n1616), 
            .I1(VCC_net), .CO(n28183));
    SB_LUT4 encoder0_position_23__I_0_add_1096_13_lut (.I0(GND_net), .I1(n1617), 
            .I2(VCC_net), .I3(n28181), .O(n1670)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_13 (.CI(n28181), .I0(n1617), 
            .I1(VCC_net), .CO(n28182));
    SB_LUT4 encoder0_position_23__I_0_add_1096_12_lut (.I0(GND_net), .I1(n1618), 
            .I2(VCC_net), .I3(n28180), .O(n1671)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_12 (.CI(n28180), .I0(n1618), 
            .I1(VCC_net), .CO(n28181));
    SB_LUT4 encoder0_position_23__I_0_add_1096_11_lut (.I0(GND_net), .I1(n1619), 
            .I2(VCC_net), .I3(n28179), .O(n1672)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_11 (.CI(n28179), .I0(n1619), 
            .I1(VCC_net), .CO(n28180));
    SB_LUT4 encoder0_position_23__I_0_add_1096_10_lut (.I0(GND_net), .I1(n1620), 
            .I2(VCC_net), .I3(n28178), .O(n1673)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_10 (.CI(n28178), .I0(n1620), 
            .I1(VCC_net), .CO(n28179));
    SB_LUT4 encoder0_position_23__I_0_add_1096_9_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n28177), .O(n1674)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14095_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n34118), .I3(GND_net), .O(n18884));   // verilog/coms.v(127[12] 300[6])
    defparam i14095_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4951));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1096_9 (.CI(n28177), .I0(n1621), 
            .I1(VCC_net), .CO(n28178));
    SB_LUT4 encoder0_position_23__I_0_add_1096_8_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n28176), .O(n1675)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_8 (.CI(n28176), .I0(n1622), 
            .I1(VCC_net), .CO(n28177));
    SB_LUT4 encoder0_position_23__I_0_add_1096_7_lut (.I0(GND_net), .I1(n1623), 
            .I2(GND_net), .I3(n28175), .O(n1676)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_7 (.CI(n28175), .I0(n1623), 
            .I1(GND_net), .CO(n28176));
    SB_LUT4 encoder0_position_23__I_0_add_1096_6_lut (.I0(GND_net), .I1(n1624), 
            .I2(GND_net), .I3(n28174), .O(n1677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14096_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n34118), .I3(GND_net), .O(n18885));   // verilog/coms.v(127[12] 300[6])
    defparam i14096_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1096_6 (.CI(n28174), .I0(n1624), 
            .I1(GND_net), .CO(n28175));
    SB_LUT4 encoder0_position_23__I_0_add_1096_5_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n28173), .O(n1678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_5 (.CI(n28173), .I0(n1625), 
            .I1(VCC_net), .CO(n28174));
    SB_LUT4 encoder0_position_23__I_0_add_1096_4_lut (.I0(GND_net), .I1(n1626), 
            .I2(GND_net), .I3(n28172), .O(n1679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_4 (.CI(n28172), .I0(n1626), 
            .I1(GND_net), .CO(n28173));
    SB_LUT4 encoder0_position_23__I_0_add_1096_3_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n28171), .O(n1680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_3 (.CI(n28171), .I0(n1627), 
            .I1(VCC_net), .CO(n28172));
    SB_LUT4 encoder0_position_23__I_0_add_1096_2_lut (.I0(GND_net), .I1(n770), 
            .I2(GND_net), .I3(VCC_net), .O(n1681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_2 (.CI(VCC_net), .I0(n770), 
            .I1(GND_net), .CO(n28171));
    SB_LUT4 encoder0_position_23__I_0_add_1043_19_lut (.I0(GND_net), .I1(n1532), 
            .I2(VCC_net), .I3(n28170), .O(n1585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1043_18_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n28169), .O(n1586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n31596));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n19194));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n19193));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n19192));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n19191));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n19190));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n19189));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n19188));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n31590));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    SB_CARRY encoder0_position_23__I_0_add_1043_18 (.CI(n28169), .I0(n1533), 
            .I1(VCC_net), .CO(n28170));
    SB_LUT4 i14097_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n34118), .I3(GND_net), .O(n18886));   // verilog/coms.v(127[12] 300[6])
    defparam i14097_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1707 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5054));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i4_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_5054), .I2(control_mode[2]), 
            .I3(GND_net), .O(n17027));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14098_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n34118), .I3(GND_net), .O(n18887));   // verilog/coms.v(127[12] 300[6])
    defparam i14098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1708 (.I0(control_mode[0]), .I1(control_mode[1]), 
            .I2(n17027), .I3(GND_net), .O(n15_adj_4928));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i2_3_lut_adj_1708.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_72_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4928), .I3(n15_adj_4936), .O(motor_state_23__N_82[23]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_72_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i24_3_lut (.I0(encoder0_position_scaled[22]), .I1(motor_state_23__N_82[23]), 
            .I2(n15), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(165[5] 168[10])
    defparam mux_70_i24_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i14099_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n34118), .I3(GND_net), .O(n18888));   // verilog/coms.v(127[12] 300[6])
    defparam i14099_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14100_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n34118), .I3(GND_net), .O(n18889));   // verilog/coms.v(127[12] 300[6])
    defparam i14100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14101_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n34118), .I3(GND_net), .O(n18890));   // verilog/coms.v(127[12] 300[6])
    defparam i14101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4950));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4949));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14102_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n34118), .I3(GND_net), .O(n18891));   // verilog/coms.v(127[12] 300[6])
    defparam i14102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1373_3_lut (.I0(n2010), .I1(n2063), 
            .I2(n2026), .I3(GND_net), .O(n29_adj_5022));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14103_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n34118), .I3(GND_net), .O(n18892));   // verilog/coms.v(127[12] 300[6])
    defparam i14103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1374_3_lut (.I0(n2011), .I1(n2064), 
            .I2(n2026), .I3(GND_net), .O(n27_adj_5021));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1365_3_lut (.I0(n2002), .I1(n2055), 
            .I2(n2026), .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1381_3_lut (.I0(n2018), .I1(n2071), 
            .I2(n2026), .I3(GND_net), .O(n13_adj_5019));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14104_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n34118), .I3(GND_net), .O(n18893));   // verilog/coms.v(127[12] 300[6])
    defparam i14104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30575_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n32359));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i30575_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 encoder0_position_23__I_0_i1368_3_lut (.I0(n2005), .I1(n2058), 
            .I2(n2026), .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26744_3_lut (.I0(encoder0_position[18]), .I1(n33126), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n679));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut_adj_1709 (.I0(n2020), .I1(n35924), .I2(n2026), .I3(n2019), 
            .O(n5_adj_4886));
    defparam i16_4_lut_adj_1709.LUT_INIT = 16'hac0c;
    SB_LUT4 i29828_3_lut (.I0(n775), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n35956));
    defparam i29828_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 encoder0_position_23__I_0_i1363_3_lut (.I0(n2000), .I1(n2053), 
            .I2(n2026), .I3(GND_net), .O(n49));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1366_3_lut (.I0(n2003), .I1(n2056), 
            .I2(n2026), .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(n35956), .I1(n5_adj_4886), .I2(n35957), 
            .I3(n2026), .O(n30964));
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'h88c0;
    SB_LUT4 i14105_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n34118), .I3(GND_net), .O(n18894));   // verilog/coms.v(127[12] 300[6])
    defparam i14105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1711 (.I0(n2016), .I1(n29_adj_5022), .I2(n2069), 
            .I3(n2026), .O(n24_adj_4875));
    defparam i4_4_lut_adj_1711.LUT_INIT = 16'heefc;
    SB_LUT4 i2_4_lut_adj_1712 (.I0(n30964), .I1(n2001), .I2(n2054), .I3(n2026), 
            .O(n22_adj_4877));
    defparam i2_4_lut_adj_1712.LUT_INIT = 16'heefa;
    SB_LUT4 i14106_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n34118), .I3(GND_net), .O(n18895));   // verilog/coms.v(127[12] 300[6])
    defparam i14106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_adj_1713 (.I0(n2007), .I1(n49), .I2(n2060), .I3(n2026), 
            .O(n23_adj_4876));
    defparam i3_4_lut_adj_1713.LUT_INIT = 16'heefc;
    SB_LUT4 i21_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3379[2]), 
            .I3(r_SM_Main[0]), .O(n18223));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i21_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n2014), .I1(n43), .I2(n2067), .I3(n2026), 
            .O(n21_adj_4878));
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_23__I_0_i1369_3_lut (.I0(n2006), .I1(n2059), 
            .I2(n2026), .I3(GND_net), .O(n37_adj_5023));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14107_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n34118), .I3(GND_net), .O(n18896));   // verilog/coms.v(127[12] 300[6])
    defparam i14107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1376_3_lut (.I0(n2013), .I1(n2066), 
            .I2(n2026), .I3(GND_net), .O(n23_adj_5020));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i8_4_lut_adj_1715 (.I0(n2008), .I1(n27_adj_5021), .I2(n2061), 
            .I3(n2026), .O(n28));
    defparam i8_4_lut_adj_1715.LUT_INIT = 16'heefc;
    SB_LUT4 i14108_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n14410), .I3(GND_net), .O(n18897));   // verilog/coms.v(127[12] 300[6])
    defparam i14108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1716 (.I0(n2004), .I1(n45), .I2(n2057), .I3(n2026), 
            .O(n26));
    defparam i6_4_lut_adj_1716.LUT_INIT = 16'heefc;
    SB_LUT4 i7_4_lut_adj_1717 (.I0(n2012), .I1(n13_adj_5019), .I2(n2065), 
            .I3(n2026), .O(n27));
    defparam i7_4_lut_adj_1717.LUT_INIT = 16'heefc;
    SB_LUT4 i5_4_lut_adj_1718 (.I0(n2017), .I1(n23_adj_5020), .I2(n2070), 
            .I3(n2026), .O(n25_adj_4874));
    defparam i5_4_lut_adj_1718.LUT_INIT = 16'heefc;
    SB_LUT4 i14109_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n14410), .I3(GND_net), .O(n18898));   // verilog/coms.v(127[12] 300[6])
    defparam i14109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n18223), 
            .I3(rx_data_ready), .O(n31970));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i14110_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n14410), .I3(GND_net), .O(n18899));   // verilog/coms.v(127[12] 300[6])
    defparam i14110_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_17_lut (.I0(GND_net), .I1(n1534), 
            .I2(VCC_net), .I3(n28168), .O(n1587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1719 (.I0(n2009), .I1(n39), .I2(n2062), .I3(n2026), 
            .O(n30));
    defparam i10_4_lut_adj_1719.LUT_INIT = 16'heefc;
    SB_LUT4 i16_4_lut_adj_1720 (.I0(n21_adj_4878), .I1(n23_adj_4876), .I2(n22_adj_4877), 
            .I3(n24_adj_4875), .O(n36));
    defparam i16_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_23__I_0_add_1043_17 (.CI(n28168), .I0(n1534), 
            .I1(VCC_net), .CO(n28169));
    SB_LUT4 i14111_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n14410), .I3(GND_net), .O(n18900));   // verilog/coms.v(127[12] 300[6])
    defparam i14111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut_adj_1721 (.I0(n2015), .I1(n37_adj_5023), .I2(n2068), 
            .I3(n2026), .O(n29));
    defparam i9_4_lut_adj_1721.LUT_INIT = 16'heefc;
    SB_LUT4 i17_4_lut (.I0(n25_adj_4874), .I1(n27), .I2(n26), .I3(n28), 
            .O(n37));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30847_4_lut (.I0(n37), .I1(n29), .I2(n36), .I3(n30), .O(n24674));
    defparam i30847_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14112_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n14410), .I3(GND_net), .O(n18901));   // verilog/coms.v(127[12] 300[6])
    defparam i14112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14113_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n14410), .I3(GND_net), .O(n18902));   // verilog/coms.v(127[12] 300[6])
    defparam i14113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_16_lut (.I0(GND_net), .I1(n1535), 
            .I2(VCC_net), .I3(n28167), .O(n1588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4948));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14114_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n14410), .I3(GND_net), .O(n18903));   // verilog/coms.v(127[12] 300[6])
    defparam i14114_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1043_16 (.CI(n28167), .I0(n1535), 
            .I1(VCC_net), .CO(n28168));
    SB_LUT4 i14115_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n14410), .I3(GND_net), .O(n18904));   // verilog/coms.v(127[12] 300[6])
    defparam i14115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_15_lut (.I0(GND_net), .I1(n1536), 
            .I2(VCC_net), .I3(n28166), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_15 (.CI(n28166), .I0(n1536), 
            .I1(VCC_net), .CO(n28167));
    SB_LUT4 i14116_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n14410), .I3(GND_net), .O(n18905));   // verilog/coms.v(127[12] 300[6])
    defparam i14116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_14_lut (.I0(GND_net), .I1(n1537), 
            .I2(VCC_net), .I3(n28165), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_14 (.CI(n28165), .I0(n1537), 
            .I1(VCC_net), .CO(n28166));
    SB_LUT4 i14117_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n14410), .I3(GND_net), .O(n18906));   // verilog/coms.v(127[12] 300[6])
    defparam i14117_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_13_lut (.I0(GND_net), .I1(n1538), 
            .I2(VCC_net), .I3(n28164), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_13 (.CI(n28164), .I0(n1538), 
            .I1(VCC_net), .CO(n28165));
    SB_LUT4 encoder0_position_23__I_0_add_1043_12_lut (.I0(GND_net), .I1(n1539), 
            .I2(VCC_net), .I3(n28163), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_12 (.CI(n28163), .I0(n1539), 
            .I1(VCC_net), .CO(n28164));
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1043_11_lut (.I0(GND_net), .I1(n1540), 
            .I2(VCC_net), .I3(n28162), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_11 (.CI(n28162), .I0(n1540), 
            .I1(VCC_net), .CO(n28163));
    SB_LUT4 i14118_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n14410), .I3(GND_net), .O(n18907));   // verilog/coms.v(127[12] 300[6])
    defparam i14118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_10_lut (.I0(GND_net), .I1(n1541), 
            .I2(VCC_net), .I3(n28161), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_10 (.CI(n28161), .I0(n1541), 
            .I1(VCC_net), .CO(n28162));
    SB_LUT4 encoder0_position_23__I_0_add_1043_9_lut (.I0(GND_net), .I1(n1542), 
            .I2(VCC_net), .I3(n28160), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_9 (.CI(n28160), .I0(n1542), 
            .I1(VCC_net), .CO(n28161));
    SB_LUT4 encoder0_position_23__I_0_add_1043_8_lut (.I0(GND_net), .I1(n1543), 
            .I2(VCC_net), .I3(n28159), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30448_2_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(\ID_READOUT_FSM.state_2__N_207 ));   // verilog/TinyFPGA_B.v(241[7:11])
    defparam i30448_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_adj_1722 (.I0(n16906), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n16908));
    defparam i1_2_lut_adj_1722.LUT_INIT = 16'heeee;
    SB_LUT4 i29609_4_lut (.I0(n27_adj_4982), .I1(n15_adj_4976), .I2(n13_adj_4975), 
            .I3(n11_adj_4973), .O(n36005));
    defparam i29609_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY encoder0_position_23__I_0_add_1043_8 (.CI(n28159), .I0(n1543), 
            .I1(VCC_net), .CO(n28160));
    SB_LUT4 encoder0_position_23__I_0_add_1043_7_lut (.I0(GND_net), .I1(n1544), 
            .I2(GND_net), .I3(n28158), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_7 (.CI(n28158), .I0(n1544), 
            .I1(GND_net), .CO(n28159));
    SB_LUT4 encoder0_position_23__I_0_add_1043_6_lut (.I0(GND_net), .I1(n1545), 
            .I2(GND_net), .I3(n28157), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14119_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n14410), .I3(GND_net), .O(n18908));   // verilog/coms.v(127[12] 300[6])
    defparam i14119_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1043_6 (.CI(n28157), .I0(n1545), 
            .I1(GND_net), .CO(n28158));
    SB_LUT4 encoder0_position_23__I_0_add_1043_5_lut (.I0(GND_net), .I1(n1546), 
            .I2(VCC_net), .I3(n28156), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_5 (.CI(n28156), .I0(n1546), 
            .I1(VCC_net), .CO(n28157));
    SB_LUT4 i29903_4_lut (.I0(n9_adj_4971), .I1(n7_adj_4969), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n36300));
    defparam i29903_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 encoder0_position_23__I_0_add_1043_4_lut (.I0(GND_net), .I1(n1547), 
            .I2(GND_net), .I3(n28155), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_4 (.CI(n28155), .I0(n1547), 
            .I1(GND_net), .CO(n28156));
    SB_LUT4 encoder0_position_23__I_0_add_1043_3_lut (.I0(GND_net), .I1(n1548), 
            .I2(VCC_net), .I3(n28154), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30073_4_lut (.I0(n15_adj_4976), .I1(n13_adj_4975), .I2(n11_adj_4973), 
            .I3(n36300), .O(n36470));
    defparam i30073_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30071_4_lut (.I0(n21_adj_4979), .I1(n19_adj_4978), .I2(n17_adj_4977), 
            .I3(n36470), .O(n36468));
    defparam i30071_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY encoder0_position_23__I_0_add_1043_3 (.CI(n28154), .I0(n1548), 
            .I1(VCC_net), .CO(n28155));
    SB_LUT4 i29611_4_lut (.I0(n27_adj_4982), .I1(n25_adj_4981), .I2(n23_adj_4980), 
            .I3(n36468), .O(n36007));
    defparam i29611_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 encoder0_position_23__I_0_add_1043_2_lut (.I0(GND_net), .I1(n769), 
            .I2(GND_net), .I3(VCC_net), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_3291_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4914), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n513));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14120_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n14410), .I3(GND_net), .O(n18909));   // verilog/coms.v(127[12] 300[6])
    defparam i14120_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1043_2 (.CI(VCC_net), .I0(n769), 
            .I1(GND_net), .CO(n28154));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4947));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_732_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4967));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i30222_3_lut (.I0(n4_adj_4967), .I1(pwm_setpoint[13]), .I2(n27_adj_4982), 
            .I3(GND_net), .O(n36619));   // verilog/pwm.v(21[8:24])
    defparam i30222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_990_18_lut (.I0(GND_net), .I1(n1454), 
            .I2(VCC_net), .I3(n28153), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_990_17_lut (.I0(GND_net), .I1(n1455), 
            .I2(VCC_net), .I3(n28152), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_17 (.CI(n28152), .I0(n1455), 
            .I1(VCC_net), .CO(n28153));
    SB_LUT4 encoder0_position_23__I_0_add_990_16_lut (.I0(GND_net), .I1(n1456), 
            .I2(VCC_net), .I3(n28151), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_16 (.CI(n28151), .I0(n1456), 
            .I1(VCC_net), .CO(n28152));
    SB_LUT4 encoder0_position_23__I_0_add_990_15_lut (.I0(GND_net), .I1(n1457), 
            .I2(VCC_net), .I3(n28150), .O(n1510)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_732_i30_3_lut (.I0(n12_adj_4974), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30_adj_4984));   // verilog/pwm.v(21[8:24])
    defparam LessThan_732_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30223_3_lut (.I0(n36619), .I1(pwm_setpoint[14]), .I2(n29_adj_4983), 
            .I3(GND_net), .O(n36620));   // verilog/pwm.v(21[8:24])
    defparam i30223_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_15 (.CI(n28150), .I0(n1457), 
            .I1(VCC_net), .CO(n28151));
    SB_LUT4 encoder0_position_23__I_0_add_990_14_lut (.I0(GND_net), .I1(n1458), 
            .I2(VCC_net), .I3(n28149), .O(n1511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_14 (.CI(n28149), .I0(n1458), 
            .I1(VCC_net), .CO(n28150));
    SB_LUT4 mux_3291_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4915), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n425));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29605_4_lut (.I0(n33_adj_4986), .I1(n31_adj_4985), .I2(n29_adj_4983), 
            .I3(n36005), .O(n36001));
    defparam i29605_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30336_4_lut (.I0(n30_adj_4984), .I1(n10_adj_4972), .I2(n35), 
            .I3(n35999), .O(n36733));   // verilog/pwm.v(21[8:24])
    defparam i30336_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_23__I_0_add_990_13_lut (.I0(GND_net), .I1(n1459), 
            .I2(VCC_net), .I3(n28148), .O(n1512)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_13 (.CI(n28148), .I0(n1459), 
            .I1(VCC_net), .CO(n28149));
    SB_LUT4 encoder0_position_23__I_0_add_990_12_lut (.I0(GND_net), .I1(n1460), 
            .I2(VCC_net), .I3(n28147), .O(n1513)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30208_3_lut (.I0(n36620), .I1(pwm_setpoint[15]), .I2(n31_adj_4985), 
            .I3(GND_net), .O(n36605));   // verilog/pwm.v(21[8:24])
    defparam i30208_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_12 (.CI(n28147), .I0(n1460), 
            .I1(VCC_net), .CO(n28148));
    SB_LUT4 encoder0_position_23__I_0_add_990_11_lut (.I0(GND_net), .I1(n1461), 
            .I2(VCC_net), .I3(n28146), .O(n1514)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30224_3_lut (.I0(n6_adj_4968), .I1(pwm_setpoint[10]), .I2(n21_adj_4979), 
            .I3(GND_net), .O(n36621));   // verilog/pwm.v(21[8:24])
    defparam i30224_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_11 (.CI(n28146), .I0(n1461), 
            .I1(VCC_net), .CO(n28147));
    SB_LUT4 i30225_3_lut (.I0(n36621), .I1(pwm_setpoint[11]), .I2(n23_adj_4980), 
            .I3(GND_net), .O(n36622));   // verilog/pwm.v(21[8:24])
    defparam i30225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_990_10_lut (.I0(GND_net), .I1(n1462), 
            .I2(VCC_net), .I3(n28145), .O(n1515)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29893_4_lut (.I0(n23_adj_4980), .I1(n21_adj_4979), .I2(n19_adj_4978), 
            .I3(n36013), .O(n36290));
    defparam i29893_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY encoder0_position_23__I_0_add_990_10 (.CI(n28145), .I0(n1462), 
            .I1(VCC_net), .CO(n28146));
    SB_LUT4 i30147_3_lut (.I0(n8_adj_4970), .I1(pwm_setpoint[9]), .I2(n19_adj_4978), 
            .I3(GND_net), .O(n36544));   // verilog/pwm.v(21[8:24])
    defparam i30147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_990_9_lut (.I0(GND_net), .I1(n1463), 
            .I2(VCC_net), .I3(n28144), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_9 (.CI(n28144), .I0(n1463), 
            .I1(VCC_net), .CO(n28145));
    SB_LUT4 encoder0_position_23__I_0_add_990_8_lut (.I0(GND_net), .I1(n1464), 
            .I2(VCC_net), .I3(n28143), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30206_3_lut (.I0(n36622), .I1(pwm_setpoint[12]), .I2(n25_adj_4981), 
            .I3(GND_net), .O(n36603));   // verilog/pwm.v(21[8:24])
    defparam i30206_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_990_8 (.CI(n28143), .I0(n1464), 
            .I1(VCC_net), .CO(n28144));
    SB_LUT4 encoder0_position_23__I_0_add_990_7_lut (.I0(GND_net), .I1(n1465), 
            .I2(GND_net), .I3(n28142), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30153_4_lut (.I0(n33_adj_4986), .I1(n31_adj_4985), .I2(n29_adj_4983), 
            .I3(n36007), .O(n36550));
    defparam i30153_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_23__I_0_add_990_7 (.CI(n28142), .I0(n1465), 
            .I1(GND_net), .CO(n28143));
    SB_LUT4 i30387_4_lut (.I0(n36605), .I1(n36733), .I2(n35), .I3(n36001), 
            .O(n36784));   // verilog/pwm.v(21[8:24])
    defparam i30387_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30218_4_lut (.I0(n36603), .I1(n36544), .I2(n25_adj_4981), 
            .I3(n36290), .O(n36615));   // verilog/pwm.v(21[8:24])
    defparam i30218_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 encoder0_position_23__I_0_add_990_6_lut (.I0(GND_net), .I1(n1466), 
            .I2(GND_net), .I3(n28141), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30391_4_lut (.I0(n36615), .I1(n36784), .I2(n35), .I3(n36550), 
            .O(n36788));   // verilog/pwm.v(21[8:24])
    defparam i30391_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30392_3_lut (.I0(n36788), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n36789));   // verilog/pwm.v(21[8:24])
    defparam i30392_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_990_6 (.CI(n28141), .I0(n1466), 
            .I1(GND_net), .CO(n28142));
    SB_LUT4 encoder0_position_23__I_0_add_990_5_lut (.I0(GND_net), .I1(n1467), 
            .I2(VCC_net), .I3(n28140), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30390_3_lut (.I0(n36789), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n36787));   // verilog/pwm.v(21[8:24])
    defparam i30390_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_990_5 (.CI(n28140), .I0(n1467), 
            .I1(VCC_net), .CO(n28141));
    SB_LUT4 i30316_3_lut (.I0(n36787), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n36713));   // verilog/pwm.v(21[8:24])
    defparam i30316_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_add_990_4_lut (.I0(GND_net), .I1(n1468), 
            .I2(GND_net), .I3(n28139), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_4 (.CI(n28139), .I0(n1468), 
            .I1(GND_net), .CO(n28140));
    SB_LUT4 i30317_3_lut (.I0(n36713), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n36714));   // verilog/pwm.v(21[8:24])
    defparam i30317_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_add_990_3_lut (.I0(GND_net), .I1(n1469), 
            .I2(VCC_net), .I3(n28138), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_3 (.CI(n28138), .I0(n1469), 
            .I1(VCC_net), .CO(n28139));
    SB_LUT4 encoder0_position_23__I_0_add_990_2_lut (.I0(GND_net), .I1(n768), 
            .I2(GND_net), .I3(VCC_net), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_2 (.CI(VCC_net), .I0(n768), 
            .I1(GND_net), .CO(n28138));
    SB_LUT4 encoder0_position_23__I_0_add_937_17_lut (.I0(GND_net), .I1(n1376), 
            .I2(VCC_net), .I3(n28137), .O(n1429)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_937_16_lut (.I0(GND_net), .I1(n1377), 
            .I2(VCC_net), .I3(n28136), .O(n1430)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_16 (.CI(n28136), .I0(n1377), 
            .I1(VCC_net), .CO(n28137));
    SB_LUT4 encoder0_position_23__I_0_add_937_15_lut (.I0(GND_net), .I1(n1378), 
            .I2(VCC_net), .I3(n28135), .O(n1431)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_15 (.CI(n28135), .I0(n1378), 
            .I1(VCC_net), .CO(n28136));
    SB_LUT4 i30214_3_lut (.I0(n36714), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n36611));   // verilog/pwm.v(21[8:24])
    defparam i30214_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_add_937_14_lut (.I0(GND_net), .I1(n1379), 
            .I2(VCC_net), .I3(n28134), .O(n1432)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_14 (.CI(n28134), .I0(n1379), 
            .I1(VCC_net), .CO(n28135));
    SB_LUT4 encoder0_position_23__I_0_add_937_13_lut (.I0(GND_net), .I1(n1380), 
            .I2(VCC_net), .I3(n28133), .O(n1433)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_13 (.CI(n28133), .I0(n1380), 
            .I1(VCC_net), .CO(n28134));
    SB_LUT4 mux_3291_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4916), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_937_12_lut (.I0(GND_net), .I1(n1381), 
            .I2(VCC_net), .I3(n28132), .O(n1434)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_12 (.CI(n28132), .I0(n1381), 
            .I1(VCC_net), .CO(n28133));
    SB_LUT4 encoder0_position_23__I_0_add_937_11_lut (.I0(GND_net), .I1(n1382), 
            .I2(VCC_net), .I3(n28131), .O(n1435)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_11 (.CI(n28131), .I0(n1382), 
            .I1(VCC_net), .CO(n28132));
    SB_LUT4 encoder0_position_23__I_0_add_937_10_lut (.I0(GND_net), .I1(n1383), 
            .I2(VCC_net), .I3(n28130), .O(n1436)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_10 (.CI(n28130), .I0(n1383), 
            .I1(VCC_net), .CO(n28131));
    SB_LUT4 encoder0_position_23__I_0_add_937_9_lut (.I0(GND_net), .I1(n1384), 
            .I2(VCC_net), .I3(n28129), .O(n1437)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_9 (.CI(n28129), .I0(n1384), 
            .I1(VCC_net), .CO(n28130));
    SB_LUT4 encoder0_position_23__I_0_add_937_8_lut (.I0(GND_net), .I1(n1385), 
            .I2(VCC_net), .I3(n28128), .O(n1438)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_8 (.CI(n28128), .I0(n1385), 
            .I1(VCC_net), .CO(n28129));
    SB_LUT4 encoder0_position_23__I_0_add_937_7_lut (.I0(GND_net), .I1(n1386), 
            .I2(GND_net), .I3(n28127), .O(n1439)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_7 (.CI(n28127), .I0(n1386), 
            .I1(GND_net), .CO(n28128));
    SB_LUT4 encoder0_position_23__I_0_add_937_6_lut (.I0(GND_net), .I1(n1387), 
            .I2(GND_net), .I3(n28126), .O(n1440)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_6 (.CI(n28126), .I0(n1387), 
            .I1(GND_net), .CO(n28127));
    SB_LUT4 encoder0_position_23__I_0_add_937_5_lut (.I0(GND_net), .I1(n1388), 
            .I2(VCC_net), .I3(n28125), .O(n1441)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_5 (.CI(n28125), .I0(n1388), 
            .I1(VCC_net), .CO(n28126));
    SB_CARRY add_28_20 (.CI(n27652), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n27653));
    SB_LUT4 encoder0_position_23__I_0_add_937_4_lut (.I0(GND_net), .I1(n1389), 
            .I2(GND_net), .I3(n28124), .O(n1442)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_4 (.CI(n28124), .I0(n1389), 
            .I1(GND_net), .CO(n28125));
    SB_LUT4 encoder0_position_23__I_0_add_937_3_lut (.I0(GND_net), .I1(n1390), 
            .I2(VCC_net), .I3(n28123), .O(n1443)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_3 (.CI(n28123), .I0(n1390), 
            .I1(VCC_net), .CO(n28124));
    SB_LUT4 i14121_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n14410), .I3(GND_net), .O(n18910));   // verilog/coms.v(127[12] 300[6])
    defparam i14121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_937_2_lut (.I0(GND_net), .I1(n767), 
            .I2(GND_net), .I3(VCC_net), .O(n1444)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14122_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n14410), .I3(GND_net), .O(n18911));   // verilog/coms.v(127[12] 300[6])
    defparam i14122_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_937_2 (.CI(VCC_net), .I0(n767), 
            .I1(GND_net), .CO(n28123));
    SB_LUT4 encoder0_position_23__I_0_add_884_16_lut (.I0(GND_net), .I1(n1298), 
            .I2(VCC_net), .I3(n28122), .O(n1351)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14123_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n14410), .I3(GND_net), .O(n18912));   // verilog/coms.v(127[12] 300[6])
    defparam i14123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_884_15_lut (.I0(GND_net), .I1(n1299), 
            .I2(VCC_net), .I3(n28121), .O(n1352)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_15 (.CI(n28121), .I0(n1299), 
            .I1(VCC_net), .CO(n28122));
    SB_LUT4 encoder0_position_23__I_0_add_884_14_lut (.I0(GND_net), .I1(n1300), 
            .I2(VCC_net), .I3(n28120), .O(n1353)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_14 (.CI(n28120), .I0(n1300), 
            .I1(VCC_net), .CO(n28121));
    SB_LUT4 encoder0_position_23__I_0_add_884_13_lut (.I0(GND_net), .I1(n1301), 
            .I2(VCC_net), .I3(n28119), .O(n1354)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_13 (.CI(n28119), .I0(n1301), 
            .I1(VCC_net), .CO(n28120));
    SB_LUT4 encoder0_position_23__I_0_add_884_12_lut (.I0(GND_net), .I1(n1302), 
            .I2(VCC_net), .I3(n28118), .O(n1355)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_12 (.CI(n28118), .I0(n1302), 
            .I1(VCC_net), .CO(n28119));
    SB_LUT4 i14124_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n14410), .I3(GND_net), .O(n18913));   // verilog/coms.v(127[12] 300[6])
    defparam i14124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_884_11_lut (.I0(GND_net), .I1(n1303), 
            .I2(VCC_net), .I3(n28117), .O(n1356)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_11 (.CI(n28117), .I0(n1303), 
            .I1(VCC_net), .CO(n28118));
    SB_LUT4 encoder0_position_23__I_0_add_884_10_lut (.I0(GND_net), .I1(n1304), 
            .I2(VCC_net), .I3(n28116), .O(n1357)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n27640), .O(n612)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14125_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n14410), .I3(GND_net), .O(n18914));   // verilog/coms.v(127[12] 300[6])
    defparam i14125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14126_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n14410), .I3(GND_net), .O(n18915));   // verilog/coms.v(127[12] 300[6])
    defparam i14126_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_10 (.CI(n28116), .I0(n1304), 
            .I1(VCC_net), .CO(n28117));
    SB_LUT4 i14127_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n14410), .I3(GND_net), .O(n18916));   // verilog/coms.v(127[12] 300[6])
    defparam i14127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_884_9_lut (.I0(GND_net), .I1(n1305), 
            .I2(VCC_net), .I3(n28115), .O(n1358)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n27651), .O(n601)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14128_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n14410), .I3(GND_net), .O(n18917));   // verilog/coms.v(127[12] 300[6])
    defparam i14128_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_9 (.CI(n28115), .I0(n1305), 
            .I1(VCC_net), .CO(n28116));
    SB_CARRY add_28_19 (.CI(n27651), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n27652));
    SB_LUT4 i14129_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n14410), .I3(GND_net), .O(n18918));   // verilog/coms.v(127[12] 300[6])
    defparam i14129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_884_8_lut (.I0(GND_net), .I1(n1306), 
            .I2(VCC_net), .I3(n28114), .O(n1359)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_8 (.CI(n27640), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n27641));
    SB_LUT4 i14130_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n14410), .I3(GND_net), .O(n18919));   // verilog/coms.v(127[12] 300[6])
    defparam i14130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14131_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n14410), .I3(GND_net), .O(n18920));   // verilog/coms.v(127[12] 300[6])
    defparam i14131_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_8 (.CI(n28114), .I0(n1306), 
            .I1(VCC_net), .CO(n28115));
    SB_LUT4 encoder0_position_23__I_0_add_884_7_lut (.I0(GND_net), .I1(n1307), 
            .I2(GND_net), .I3(n28113), .O(n1360)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n1172), .I3(data_ready), .O(n31596));   // verilog/TinyFPGA_B.v(237[10] 261[6])
    defparam i12_4_lut_4_lut.LUT_INIT = 16'hce8a;
    SB_LUT4 i14132_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n14410), .I3(GND_net), .O(n18921));   // verilog/coms.v(127[12] 300[6])
    defparam i14132_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_7 (.CI(n28113), .I0(n1307), 
            .I1(GND_net), .CO(n28114));
    SB_LUT4 add_28_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n27639), .O(n613)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_884_6_lut (.I0(GND_net), .I1(n1308), 
            .I2(GND_net), .I3(n28112), .O(n1361)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14133_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n14410), .I3(GND_net), .O(n18922));   // verilog/coms.v(127[12] 300[6])
    defparam i14133_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_6 (.CI(n28112), .I0(n1308), 
            .I1(GND_net), .CO(n28113));
    SB_LUT4 encoder0_position_23__I_0_add_884_5_lut (.I0(GND_net), .I1(n1309), 
            .I2(VCC_net), .I3(n28111), .O(n1362)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_5 (.CI(n28111), .I0(n1309), 
            .I1(VCC_net), .CO(n28112));
    SB_LUT4 encoder0_position_23__I_0_add_884_4_lut (.I0(GND_net), .I1(n1310), 
            .I2(GND_net), .I3(n28110), .O(n1363)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_4 (.CI(n28110), .I0(n1310), 
            .I1(GND_net), .CO(n28111));
    SB_LUT4 i14134_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n14410), .I3(GND_net), .O(n18923));   // verilog/coms.v(127[12] 300[6])
    defparam i14134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_884_3_lut (.I0(GND_net), .I1(n1311), 
            .I2(VCC_net), .I3(n28109), .O(n1364)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14135_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n14410), .I3(GND_net), .O(n18924));   // verilog/coms.v(127[12] 300[6])
    defparam i14135_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_3 (.CI(n28109), .I0(n1311), 
            .I1(VCC_net), .CO(n28110));
    SB_LUT4 encoder0_position_23__I_0_add_884_2_lut (.I0(GND_net), .I1(n523), 
            .I2(GND_net), .I3(VCC_net), .O(n1365)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14136_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n14410), .I3(GND_net), .O(n18925));   // verilog/coms.v(127[12] 300[6])
    defparam i14136_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_884_2 (.CI(VCC_net), .I0(n523), 
            .I1(GND_net), .CO(n28109));
    SB_LUT4 encoder0_position_23__I_0_add_831_15_lut (.I0(GND_net), .I1(n1220), 
            .I2(VCC_net), .I3(n28108), .O(n1273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n27650), .O(n602)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_831_14_lut (.I0(GND_net), .I1(n1221), 
            .I2(VCC_net), .I3(n28107), .O(n1274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_14 (.CI(n28107), .I0(n1221), 
            .I1(VCC_net), .CO(n28108));
    SB_LUT4 encoder0_position_23__I_0_add_831_13_lut (.I0(GND_net), .I1(n1222), 
            .I2(VCC_net), .I3(n28106), .O(n1275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14137_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n14410), .I3(GND_net), .O(n18926));   // verilog/coms.v(127[12] 300[6])
    defparam i14137_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_28_18 (.CI(n27650), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n27651));
    SB_CARRY encoder0_position_23__I_0_add_831_13 (.CI(n28106), .I0(n1222), 
            .I1(VCC_net), .CO(n28107));
    SB_LUT4 add_28_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n27649), .O(n603)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_831_12_lut (.I0(GND_net), .I1(n1223), 
            .I2(VCC_net), .I3(n28105), .O(n1276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_12 (.CI(n28105), .I0(n1223), 
            .I1(VCC_net), .CO(n28106));
    SB_LUT4 encoder0_position_23__I_0_add_831_11_lut (.I0(GND_net), .I1(n1224), 
            .I2(VCC_net), .I3(n28104), .O(n1277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_11 (.CI(n28104), .I0(n1224), 
            .I1(VCC_net), .CO(n28105));
    SB_LUT4 i14138_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n14410), .I3(GND_net), .O(n18927));   // verilog/coms.v(127[12] 300[6])
    defparam i14138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_10_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n28103), .O(n1278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28598_1_lut (.I0(n4_adj_4962), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n34993));
    defparam i28598_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3291_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4917), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n510));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4873));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14139_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n14410), .I3(GND_net), .O(n18928));   // verilog/coms.v(127[12] 300[6])
    defparam i14139_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_28_17 (.CI(n27649), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n27650));
    SB_LUT4 i30415_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n15_adj_4867), .I3(GND_net), .O(n18163));   // verilog/TinyFPGA_B.v(251[7:11])
    defparam i30415_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_831_10 (.CI(n28103), .I0(n1225), 
            .I1(VCC_net), .CO(n28104));
    SB_LUT4 encoder0_position_23__I_0_add_831_9_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n28102), .O(n1279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_9 (.CI(n28102), .I0(n1226), 
            .I1(VCC_net), .CO(n28103));
    SB_LUT4 i14140_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n14410), .I3(GND_net), .O(n18929));   // verilog/coms.v(127[12] 300[6])
    defparam i14140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14141_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n14410), .I3(GND_net), .O(n18930));   // verilog/coms.v(127[12] 300[6])
    defparam i14141_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_28_3 (.CI(n27635), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n27636));
    SB_LUT4 add_28_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n618)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14142_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n14410), .I3(GND_net), .O(n18931));   // verilog/coms.v(127[12] 300[6])
    defparam i14142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14143_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n14410), .I3(GND_net), .O(n18932));   // verilog/coms.v(127[12] 300[6])
    defparam i14143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5111[1]), .I1(r_SM_Main_adj_5111[0]), 
            .I2(r_SM_Main_adj_5111[2]), .I3(r_SM_Main_2__N_3450[1]), .O(n37939));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i14144_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n14410), .I3(GND_net), .O(n18933));   // verilog/coms.v(127[12] 300[6])
    defparam i14144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14145_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n14410), .I3(GND_net), .O(n18934));   // verilog/coms.v(127[12] 300[6])
    defparam i14145_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_28_7 (.CI(n27639), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n27640));
    SB_LUT4 encoder0_position_23__I_0_add_831_8_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n28101), .O(n1280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_8 (.CI(n28101), .I0(n1227), 
            .I1(VCC_net), .CO(n28102));
    SB_LUT4 encoder0_position_23__I_0_add_831_7_lut (.I0(GND_net), .I1(n1228), 
            .I2(GND_net), .I3(n28100), .O(n1281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n27648), .O(n604)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_7 (.CI(n28100), .I0(n1228), 
            .I1(GND_net), .CO(n28101));
    SB_LUT4 i14146_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n14410), .I3(GND_net), .O(n18935));   // verilog/coms.v(127[12] 300[6])
    defparam i14146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14147_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n14410), .I3(GND_net), .O(n18936));   // verilog/coms.v(127[12] 300[6])
    defparam i14147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14148_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n14410), .I3(GND_net), .O(n18937));   // verilog/coms.v(127[12] 300[6])
    defparam i14148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_831_6_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n28099), .O(n1282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_6 (.CI(n28099), .I0(n1229), 
            .I1(GND_net), .CO(n28100));
    SB_LUT4 i14149_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n14410), .I3(GND_net), .O(n18938));   // verilog/coms.v(127[12] 300[6])
    defparam i14149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14150_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n14410), .I3(GND_net), .O(n18939));   // verilog/coms.v(127[12] 300[6])
    defparam i14150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13837_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n34304), .I3(GND_net), .O(n18626));   // verilog/coms.v(127[12] 300[6])
    defparam i13837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_831_5_lut (.I0(GND_net), .I1(n1230), 
            .I2(VCC_net), .I3(n28098), .O(n1283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_5 (.CI(n28098), .I0(n1230), 
            .I1(VCC_net), .CO(n28099));
    SB_LUT4 encoder0_position_23__I_0_add_831_4_lut (.I0(GND_net), .I1(n1231), 
            .I2(GND_net), .I3(n28097), .O(n1284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_4 (.CI(n28097), .I0(n1231), 
            .I1(GND_net), .CO(n28098));
    SB_LUT4 encoder0_position_23__I_0_add_831_3_lut (.I0(GND_net), .I1(n1232), 
            .I2(VCC_net), .I3(n28096), .O(n1285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_3 (.CI(n28096), .I0(n1232), 
            .I1(VCC_net), .CO(n28097));
    SB_LUT4 i13843_4_lut (.I0(state_7__N_3877[3]), .I1(data[7]), .I2(n23726), 
            .I3(n17058), .O(n18632));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13843_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_23__I_0_add_831_2_lut (.I0(GND_net), .I1(n765), 
            .I2(GND_net), .I3(VCC_net), .O(n1286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_2 (.CI(VCC_net), .I0(n765), 
            .I1(GND_net), .CO(n28096));
    SB_LUT4 i14151_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n14410), .I3(GND_net), .O(n18940));   // verilog/coms.v(127[12] 300[6])
    defparam i14151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14152_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n14410), .I3(GND_net), .O(n18941));   // verilog/coms.v(127[12] 300[6])
    defparam i14152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_778_14_lut (.I0(GND_net), .I1(n1142), 
            .I2(VCC_net), .I3(n28095), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_778_13_lut (.I0(GND_net), .I1(n1143), 
            .I2(VCC_net), .I3(n28094), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26737_3_lut (.I0(encoder0_position[19]), .I1(n33118), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n678));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26737_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_778_13 (.CI(n28094), .I0(n1143), 
            .I1(VCC_net), .CO(n28095));
    SB_LUT4 i14153_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n14410), .I3(GND_net), .O(n18942));   // verilog/coms.v(127[12] 300[6])
    defparam i14153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14154_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n14410), .I3(GND_net), .O(n18943));   // verilog/coms.v(127[12] 300[6])
    defparam i14154_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14155_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n14410), .I3(GND_net), .O(n18944));   // verilog/coms.v(127[12] 300[6])
    defparam i14155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14156_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n14410), 
            .I3(GND_net), .O(n18945));   // verilog/coms.v(127[12] 300[6])
    defparam i14156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_778_12_lut (.I0(GND_net), .I1(n1144), 
            .I2(VCC_net), .I3(n28093), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_12 (.CI(n28093), .I0(n1144), 
            .I1(VCC_net), .CO(n28094));
    SB_LUT4 i14157_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n14410), 
            .I3(GND_net), .O(n18946));   // verilog/coms.v(127[12] 300[6])
    defparam i14157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14158_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n14410), 
            .I3(GND_net), .O(n18947));   // verilog/coms.v(127[12] 300[6])
    defparam i14158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_778_11_lut (.I0(GND_net), .I1(n1145), 
            .I2(VCC_net), .I3(n28092), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_11 (.CI(n28092), .I0(n1145), 
            .I1(VCC_net), .CO(n28093));
    SB_LUT4 i29827_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(n26386), 
            .I2(start), .I3(state[0]), .O(n35879));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29827_3_lut_4_lut.LUT_INIT = 16'hf0f4;
    SB_LUT4 i13844_4_lut (.I0(state_7__N_3877[3]), .I1(data[6]), .I2(n23726), 
            .I3(n17053), .O(n18633));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i13844_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4872));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13845_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18634));   // verilog/coms.v(127[12] 300[6])
    defparam i13845_3_lut.LUT_INIT = 16'hcaca;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 encoder0_position_23__I_0_add_778_10_lut (.I0(GND_net), .I1(n1146), 
            .I2(VCC_net), .I3(n28091), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_10 (.CI(n28091), .I0(n1146), 
            .I1(VCC_net), .CO(n28092));
    SB_LUT4 encoder0_position_23__I_0_add_778_9_lut (.I0(GND_net), .I1(n1147), 
            .I2(VCC_net), .I3(n28090), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_9_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_CARRY encoder0_position_23__I_0_add_778_9 (.CI(n28090), .I0(n1147), 
            .I1(VCC_net), .CO(n28091));
    SB_LUT4 i13846_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n34304), 
            .I3(GND_net), .O(n18635));   // verilog/coms.v(127[12] 300[6])
    defparam i13846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_8_lut (.I0(GND_net), .I1(n1148), 
            .I2(VCC_net), .I3(n28089), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13847_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n34304), 
            .I3(GND_net), .O(n18636));   // verilog/coms.v(127[12] 300[6])
    defparam i13847_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_778_8 (.CI(n28089), .I0(n1148), 
            .I1(VCC_net), .CO(n28090));
    SB_LUT4 encoder0_position_23__I_0_add_778_7_lut (.I0(GND_net), .I1(n1149), 
            .I2(GND_net), .I3(n28088), .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_16 (.CI(n27648), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n27649));
    SB_CARRY encoder0_position_23__I_0_add_778_7 (.CI(n28088), .I0(n1149), 
            .I1(GND_net), .CO(n28089));
    SB_LUT4 encoder0_position_23__I_0_add_778_6_lut (.I0(GND_net), .I1(n1150), 
            .I2(GND_net), .I3(n28087), .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_6 (.CI(n28087), .I0(n1150), 
            .I1(GND_net), .CO(n28088));
    SB_LUT4 encoder0_position_23__I_0_add_778_5_lut (.I0(GND_net), .I1(n1151), 
            .I2(VCC_net), .I3(n28086), .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_5 (.CI(n28086), .I0(n1151), 
            .I1(VCC_net), .CO(n28087));
    SB_LUT4 i13848_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n34118), .I3(GND_net), .O(n18637));   // verilog/coms.v(127[12] 300[6])
    defparam i13848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_778_4_lut (.I0(GND_net), .I1(n1152), 
            .I2(GND_net), .I3(n28085), .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_4 (.CI(n28085), .I0(n1152), 
            .I1(GND_net), .CO(n28086));
    SB_LUT4 encoder0_position_23__I_0_add_778_3_lut (.I0(GND_net), .I1(n1153), 
            .I2(VCC_net), .I3(n28084), .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_3 (.CI(n28084), .I0(n1153), 
            .I1(VCC_net), .CO(n28085));
    SB_LUT4 encoder0_position_23__I_0_add_778_2_lut (.I0(GND_net), .I1(n521), 
            .I2(GND_net), .I3(VCC_net), .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13850_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n34304), .I3(GND_net), .O(n18639));   // verilog/coms.v(127[12] 300[6])
    defparam i13850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13851_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n34304), .I3(GND_net), .O(n18640));   // verilog/coms.v(127[12] 300[6])
    defparam i13851_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_778_2 (.CI(VCC_net), .I0(n521), 
            .I1(GND_net), .CO(n28084));
    SB_LUT4 i14159_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n14410), 
            .I3(GND_net), .O(n18948));   // verilog/coms.v(127[12] 300[6])
    defparam i14159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14160_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n14410), 
            .I3(GND_net), .O(n18949));   // verilog/coms.v(127[12] 300[6])
    defparam i14160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14161_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n14410), 
            .I3(GND_net), .O(n18950));   // verilog/coms.v(127[12] 300[6])
    defparam i14161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14162_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n14410), 
            .I3(GND_net), .O(n18951));   // verilog/coms.v(127[12] 300[6])
    defparam i14162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14163_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n14410), 
            .I3(GND_net), .O(n18952));   // verilog/coms.v(127[12] 300[6])
    defparam i14163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14164_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n14410), 
            .I3(GND_net), .O(n18953));   // verilog/coms.v(127[12] 300[6])
    defparam i14164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14165_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n14410), 
            .I3(GND_net), .O(n18954));   // verilog/coms.v(127[12] 300[6])
    defparam i14165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14166_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n14410), 
            .I3(GND_net), .O(n18955));   // verilog/coms.v(127[12] 300[6])
    defparam i14166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14167_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n14410), 
            .I3(GND_net), .O(n18956));   // verilog/coms.v(127[12] 300[6])
    defparam i14167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14168_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n14410), 
            .I3(GND_net), .O(n18957));   // verilog/coms.v(127[12] 300[6])
    defparam i14168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14169_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n14410), 
            .I3(GND_net), .O(n18958));   // verilog/coms.v(127[12] 300[6])
    defparam i14169_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_28_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n27635));
    SB_LUT4 encoder0_position_23__I_0_add_725_13_lut (.I0(GND_net), .I1(n1064), 
            .I2(VCC_net), .I3(n28075), .O(n1117)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_12_lut (.I0(GND_net), .I1(n1065), 
            .I2(VCC_net), .I3(n28074), .O(n1118)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_12 (.CI(n28074), .I0(n1065), 
            .I1(VCC_net), .CO(n28075));
    SB_LUT4 encoder0_position_23__I_0_add_725_11_lut (.I0(GND_net), .I1(n1066), 
            .I2(VCC_net), .I3(n28073), .O(n1119)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_11 (.CI(n28073), .I0(n1066), 
            .I1(VCC_net), .CO(n28074));
    SB_LUT4 i14170_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n14410), 
            .I3(GND_net), .O(n18959));   // verilog/coms.v(127[12] 300[6])
    defparam i14170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14171_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n14410), 
            .I3(GND_net), .O(n18960));   // verilog/coms.v(127[12] 300[6])
    defparam i14171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_725_10_lut (.I0(GND_net), .I1(n1067), 
            .I2(VCC_net), .I3(n28072), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_10 (.CI(n28072), .I0(n1067), 
            .I1(VCC_net), .CO(n28073));
    SB_LUT4 add_28_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n27647), .O(n605)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_9_lut (.I0(GND_net), .I1(n1068), 
            .I2(VCC_net), .I3(n28071), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_9 (.CI(n28071), .I0(n1068), 
            .I1(VCC_net), .CO(n28072));
    SB_LUT4 encoder0_position_23__I_0_add_725_8_lut (.I0(GND_net), .I1(n1069), 
            .I2(VCC_net), .I3(n28070), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_8 (.CI(n28070), .I0(n1069), 
            .I1(VCC_net), .CO(n28071));
    SB_LUT4 i14172_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n14410), 
            .I3(GND_net), .O(n18961));   // verilog/coms.v(127[12] 300[6])
    defparam i14172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14173_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n14410), 
            .I3(GND_net), .O(n18962));   // verilog/coms.v(127[12] 300[6])
    defparam i14173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_725_7_lut (.I0(GND_net), .I1(n1070), 
            .I2(GND_net), .I3(n28069), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_15 (.CI(n27647), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n27648));
    SB_CARRY encoder0_position_23__I_0_add_725_7 (.CI(n28069), .I0(n1070), 
            .I1(GND_net), .CO(n28070));
    SB_LUT4 encoder0_position_23__I_0_add_725_6_lut (.I0(GND_net), .I1(n1071), 
            .I2(GND_net), .I3(n28068), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_6 (.CI(n28068), .I0(n1071), 
            .I1(GND_net), .CO(n28069));
    SB_LUT4 encoder0_position_23__I_0_add_725_5_lut (.I0(GND_net), .I1(n1072), 
            .I2(VCC_net), .I3(n28067), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_5 (.CI(n28067), .I0(n1072), 
            .I1(VCC_net), .CO(n28068));
    SB_LUT4 encoder0_position_23__I_0_add_725_4_lut (.I0(GND_net), .I1(n1073), 
            .I2(GND_net), .I3(n28066), .O(n1126)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_4 (.CI(n28066), .I0(n1073), 
            .I1(GND_net), .CO(n28067));
    SB_LUT4 encoder0_position_23__I_0_add_725_3_lut (.I0(GND_net), .I1(n1074), 
            .I2(VCC_net), .I3(n28065), .O(n1127)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_3 (.CI(n28065), .I0(n1074), 
            .I1(VCC_net), .CO(n28066));
    SB_LUT4 encoder0_position_23__I_0_add_725_2_lut (.I0(GND_net), .I1(n763), 
            .I2(GND_net), .I3(VCC_net), .O(n1128)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14174_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n14410), 
            .I3(GND_net), .O(n18963));   // verilog/coms.v(127[12] 300[6])
    defparam i14174_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_725_2 (.CI(VCC_net), .I0(n763), 
            .I1(GND_net), .CO(n28065));
    SB_LUT4 i14175_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n14410), 
            .I3(GND_net), .O(n18964));   // verilog/coms.v(127[12] 300[6])
    defparam i14175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_672_12_lut (.I0(GND_net), .I1(n986), 
            .I2(VCC_net), .I3(n28064), .O(n1039)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_672_11_lut (.I0(GND_net), .I1(n987), 
            .I2(VCC_net), .I3(n28063), .O(n1040)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n27646), .O(n606)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_11 (.CI(n28063), .I0(n987), 
            .I1(VCC_net), .CO(n28064));
    SB_LUT4 encoder0_position_23__I_0_add_672_10_lut (.I0(GND_net), .I1(n988), 
            .I2(VCC_net), .I3(n28062), .O(n1041)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_10 (.CI(n28062), .I0(n988), 
            .I1(VCC_net), .CO(n28063));
    SB_LUT4 encoder0_position_23__I_0_add_672_9_lut (.I0(GND_net), .I1(n989), 
            .I2(VCC_net), .I3(n28061), .O(n1042)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_9 (.CI(n28061), .I0(n989), 
            .I1(VCC_net), .CO(n28062));
    SB_LUT4 i14176_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n14410), 
            .I3(GND_net), .O(n18965));   // verilog/coms.v(127[12] 300[6])
    defparam i14176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_672_8_lut (.I0(GND_net), .I1(n990), 
            .I2(VCC_net), .I3(n28060), .O(n1043)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_28_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n27638), .O(n614)) /* synthesis syn_instantiated=1 */ ;
    defparam add_28_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_8 (.CI(n28060), .I0(n990), 
            .I1(VCC_net), .CO(n28061));
    SB_LUT4 i14177_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n14410), 
            .I3(GND_net), .O(n18966));   // verilog/coms.v(127[12] 300[6])
    defparam i14177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_672_7_lut (.I0(GND_net), .I1(n991), 
            .I2(GND_net), .I3(n28059), .O(n1044)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_7_lut.LUT_INIT = 16'hC33C;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .data_o({quadA_debounced_adj_4922, quadB_debounced_adj_4923}), 
            .GND_net(GND_net), .n34883(n34883), .reg_B({reg_B_adj_5120}), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .VCC_net(VCC_net), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n18645(n18645), .n19185(n19185)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(193[15] 198[4])
    SB_CARRY encoder0_position_23__I_0_add_672_7 (.CI(n28059), .I0(n991), 
            .I1(GND_net), .CO(n28060));
    SB_LUT4 encoder0_position_23__I_0_add_672_6_lut (.I0(GND_net), .I1(n992), 
            .I2(GND_net), .I3(n28058), .O(n1045)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_6 (.CI(n28058), .I0(n992), 
            .I1(GND_net), .CO(n28059));
    SB_LUT4 encoder0_position_23__I_0_add_672_5_lut (.I0(GND_net), .I1(n993), 
            .I2(VCC_net), .I3(n28057), .O(n1046)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_5 (.CI(n28057), .I0(n993), 
            .I1(VCC_net), .CO(n28058));
    SB_CARRY add_28_6 (.CI(n27638), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n27639));
    SB_LUT4 encoder0_position_23__I_0_add_672_4_lut (.I0(GND_net), .I1(n994), 
            .I2(GND_net), .I3(n28056), .O(n1047)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_4 (.CI(n28056), .I0(n994), 
            .I1(GND_net), .CO(n28057));
    SB_LUT4 encoder0_position_23__I_0_add_672_3_lut (.I0(GND_net), .I1(n995), 
            .I2(VCC_net), .I3(n28055), .O(n1048)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_3 (.CI(n28055), .I0(n995), 
            .I1(VCC_net), .CO(n28056));
    SB_LUT4 encoder0_position_23__I_0_add_672_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n1049)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14178_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n14410), 
            .I3(GND_net), .O(n18967));   // verilog/coms.v(127[12] 300[6])
    defparam i14178_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_672_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n28055));
    SB_LUT4 i14179_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n14410), 
            .I3(GND_net), .O(n18968));   // verilog/coms.v(127[12] 300[6])
    defparam i14179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14180_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n14410), .I3(GND_net), .O(n18969));   // verilog/coms.v(127[12] 300[6])
    defparam i14180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_619_11_lut (.I0(GND_net), .I1(n908), 
            .I2(VCC_net), .I3(n28054), .O(n961)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_619_10_lut (.I0(GND_net), .I1(n909), 
            .I2(VCC_net), .I3(n28053), .O(n962)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_10 (.CI(n28053), .I0(n909), 
            .I1(VCC_net), .CO(n28054));
    SB_LUT4 i14181_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n14410), .I3(GND_net), .O(n18970));   // verilog/coms.v(127[12] 300[6])
    defparam i14181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_619_9_lut (.I0(GND_net), .I1(n910), 
            .I2(VCC_net), .I3(n28052), .O(n963)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14182_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n14410), .I3(GND_net), .O(n18971));   // verilog/coms.v(127[12] 300[6])
    defparam i14182_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_619_9 (.CI(n28052), .I0(n910), 
            .I1(VCC_net), .CO(n28053));
    SB_LUT4 i14183_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n14410), .I3(GND_net), .O(n18972));   // verilog/coms.v(127[12] 300[6])
    defparam i14183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_619_8_lut (.I0(GND_net), .I1(n911), 
            .I2(VCC_net), .I3(n28051), .O(n964)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_8 (.CI(n28051), .I0(n911), 
            .I1(VCC_net), .CO(n28052));
    SB_LUT4 encoder0_position_23__I_0_add_619_7_lut (.I0(GND_net), .I1(n912), 
            .I2(GND_net), .I3(n28050), .O(n965)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14184_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n14410), .I3(GND_net), .O(n18973));   // verilog/coms.v(127[12] 300[6])
    defparam i14184_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_619_7 (.CI(n28050), .I0(n912), 
            .I1(GND_net), .CO(n28051));
    SB_LUT4 encoder0_position_23__I_0_add_619_6_lut (.I0(GND_net), .I1(n913), 
            .I2(GND_net), .I3(n28049), .O(n966)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_28_14 (.CI(n27646), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n27647));
    SB_CARRY encoder0_position_23__I_0_add_619_6 (.CI(n28049), .I0(n913), 
            .I1(GND_net), .CO(n28050));
    SB_LUT4 encoder0_position_23__I_0_add_619_5_lut (.I0(GND_net), .I1(n914), 
            .I2(VCC_net), .I3(n28048), .O(n967)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_5 (.CI(n28048), .I0(n914), 
            .I1(VCC_net), .CO(n28049));
    SB_LUT4 encoder0_position_23__I_0_add_619_4_lut (.I0(GND_net), .I1(n915), 
            .I2(GND_net), .I3(n28047), .O(n968)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_4 (.CI(n28047), .I0(n915), 
            .I1(GND_net), .CO(n28048));
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 encoder0_position_23__I_0_add_619_3_lut (.I0(GND_net), .I1(n916), 
            .I2(VCC_net), .I3(n28046), .O(n969)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_3 (.CI(n28046), .I0(n916), 
            .I1(VCC_net), .CO(n28047));
    SB_LUT4 i26733_3_lut (.I0(encoder0_position[20]), .I1(n33114), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n677));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_619_2_lut (.I0(GND_net), .I1(n518), 
            .I2(GND_net), .I3(VCC_net), .O(n970)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_2_lut.LUT_INIT = 16'hC33C;
    motorControl control (.\Ki[8] (Ki[8]), .GND_net(GND_net), .IntegralLimit({IntegralLimit}), 
            .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), .\Ki[12] (Ki[12]), 
            .PWMLimit({PWMLimit}), .duty({duty}), .n37310(n37310), .\Ki[1] (Ki[1]), 
            .\Ki[0] (Ki[0]), .\Ki[2] (Ki[2]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), .\Kp[14] (Kp[14]), 
            .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), .\Kp[2] (Kp[2]), .\Ki[3] (Ki[3]), 
            .clk32MHz(clk32MHz), .\Kp[3] (Kp[3]), .\Kp[4] (Kp[4]), .\Ki[4] (Ki[4]), 
            .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), .VCC_net(VCC_net), 
            .\Kp[15] (Kp[15]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), 
            .setpoint({setpoint}), .motor_state({motor_state})) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(170[16] 182[4])
    SB_CARRY encoder0_position_23__I_0_add_619_2 (.CI(VCC_net), .I0(n518), 
            .I1(GND_net), .CO(n28046));
    SB_LUT4 encoder0_position_23__I_0_add_566_10_lut (.I0(GND_net), .I1(n830), 
            .I2(VCC_net), .I3(n28045), .O(n883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_566_9_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n28044), .O(n884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_9 (.CI(n28044), .I0(n831), 
            .I1(VCC_net), .CO(n28045));
    SB_LUT4 encoder0_position_23__I_0_add_566_8_lut (.I0(GND_net), .I1(n832), 
            .I2(VCC_net), .I3(n28043), .O(n885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_8 (.CI(n28043), .I0(n832), 
            .I1(VCC_net), .CO(n28044));
    SB_LUT4 encoder0_position_23__I_0_add_566_7_lut (.I0(GND_net), .I1(n833), 
            .I2(GND_net), .I3(n28042), .O(n886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_7 (.CI(n28042), .I0(n833), 
            .I1(GND_net), .CO(n28043));
    SB_LUT4 i19894_4_lut (.I0(n515), .I1(n677), .I2(n678), .I3(n679), 
            .O(n24676));
    defparam i19894_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 encoder0_position_23__I_0_add_566_6_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(n28041), .O(n887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_6 (.CI(n28041), .I0(n834), 
            .I1(GND_net), .CO(n28042));
    SB_LUT4 encoder0_position_23__I_0_add_566_5_lut (.I0(GND_net), .I1(n835), 
            .I2(VCC_net), .I3(n28040), .O(n888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_5 (.CI(n28040), .I0(n835), 
            .I1(VCC_net), .CO(n28041));
    SB_LUT4 encoder0_position_23__I_0_add_566_4_lut (.I0(GND_net), .I1(n836), 
            .I2(GND_net), .I3(n28039), .O(n889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_4 (.CI(n28039), .I0(n836), 
            .I1(GND_net), .CO(n28040));
    SB_LUT4 encoder0_position_23__I_0_add_566_3_lut (.I0(GND_net), .I1(n837), 
            .I2(VCC_net), .I3(n28038), .O(n890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_3 (.CI(n28038), .I0(n837), 
            .I1(VCC_net), .CO(n28039));
    SB_LUT4 encoder0_position_23__I_0_add_566_2_lut (.I0(GND_net), .I1(n517), 
            .I2(GND_net), .I3(VCC_net), .O(n891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_2 (.CI(VCC_net), .I0(n517), 
            .I1(GND_net), .CO(n28038));
    SB_LUT4 i14185_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n14410), .I3(GND_net), .O(n18974));   // verilog/coms.v(127[12] 300[6])
    defparam i14185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14186_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n14410), .I3(GND_net), .O(n18975));   // verilog/coms.v(127[12] 300[6])
    defparam i14186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14187_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n14410), .I3(GND_net), .O(n18976));   // verilog/coms.v(127[12] 300[6])
    defparam i14187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30858_4_lut (.I0(n676), .I1(n674), .I2(n675), .I3(n24676), 
            .O(n700));
    defparam i30858_4_lut.LUT_INIT = 16'h1333;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4946));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14188_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n14410), .I3(GND_net), .O(n18977));   // verilog/coms.v(127[12] 300[6])
    defparam i14188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14189_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n14410), .I3(GND_net), .O(n18978));   // verilog/coms.v(127[12] 300[6])
    defparam i14189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14190_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n14410), .I3(GND_net), .O(n18979));   // verilog/coms.v(127[12] 300[6])
    defparam i14190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4945));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4944));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14191_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n14410), .I3(GND_net), .O(n18980));   // verilog/coms.v(127[12] 300[6])
    defparam i14191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14192_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n14410), .I3(GND_net), .O(n18981));   // verilog/coms.v(127[12] 300[6])
    defparam i14192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4943));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14193_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n14410), .I3(GND_net), .O(n18982));   // verilog/coms.v(127[12] 300[6])
    defparam i14193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14194_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n14410), .I3(GND_net), .O(n18983));   // verilog/coms.v(127[12] 300[6])
    defparam i14194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14195_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n14410), .I3(GND_net), .O(n18984));   // verilog/coms.v(127[12] 300[6])
    defparam i14195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14196_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n14410), .I3(GND_net), .O(n18985));   // verilog/coms.v(127[12] 300[6])
    defparam i14196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14197_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n14410), .I3(GND_net), .O(n18986));   // verilog/coms.v(127[12] 300[6])
    defparam i14197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14198_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n14410), .I3(GND_net), .O(n18987));   // verilog/coms.v(127[12] 300[6])
    defparam i14198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14199_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n14410), .I3(GND_net), .O(n18988));   // verilog/coms.v(127[12] 300[6])
    defparam i14199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14200_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n14410), .I3(GND_net), .O(n18989));   // verilog/coms.v(127[12] 300[6])
    defparam i14200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14201_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n14410), .I3(GND_net), .O(n18990));   // verilog/coms.v(127[12] 300[6])
    defparam i14201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3291_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4912), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n515));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14202_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n14410), .I3(GND_net), .O(n18991));   // verilog/coms.v(127[12] 300[6])
    defparam i14202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14203_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n14410), .I3(GND_net), .O(n18992));   // verilog/coms.v(127[12] 300[6])
    defparam i14203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14204_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n14410), .I3(GND_net), .O(n18993));   // verilog/coms.v(127[12] 300[6])
    defparam i14204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14205_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n14410), .I3(GND_net), .O(n18994));   // verilog/coms.v(127[12] 300[6])
    defparam i14205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14206_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4893), 
            .I3(n17079), .O(n18995));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14206_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14207_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n14410), .I3(GND_net), .O(n18996));   // verilog/coms.v(127[12] 300[6])
    defparam i14207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14208_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n14410), .I3(GND_net), .O(n18997));   // verilog/coms.v(127[12] 300[6])
    defparam i14208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14209_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n14410), .I3(GND_net), .O(n18998));   // verilog/coms.v(127[12] 300[6])
    defparam i14209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14210_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n14410), .I3(GND_net), .O(n18999));   // verilog/coms.v(127[12] 300[6])
    defparam i14210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14211_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n14410), .I3(GND_net), .O(n19000));   // verilog/coms.v(127[12] 300[6])
    defparam i14211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14212_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n14410), .I3(GND_net), .O(n19001));   // verilog/coms.v(127[12] 300[6])
    defparam i14212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14213_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n14410), .I3(GND_net), .O(n19002));   // verilog/coms.v(127[12] 300[6])
    defparam i14213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14214_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n14410), .I3(GND_net), .O(n19003));   // verilog/coms.v(127[12] 300[6])
    defparam i14214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14215_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n14410), .I3(GND_net), .O(n19004));   // verilog/coms.v(127[12] 300[6])
    defparam i14215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14216_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n14410), .I3(GND_net), .O(n19005));   // verilog/coms.v(127[12] 300[6])
    defparam i14216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4871));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14217_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n14410), .I3(GND_net), .O(n19006));   // verilog/coms.v(127[12] 300[6])
    defparam i14217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14218_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n14410), .I3(GND_net), .O(n19007));   // verilog/coms.v(127[12] 300[6])
    defparam i14218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4870));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i468_3_lut (.I0(n515), .I1(n733), 
            .I2(n700), .I3(GND_net), .O(n758));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3291_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4911), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3291_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19406_2_lut (.I0(n516), .I1(n758), .I2(GND_net), .I3(GND_net), 
            .O(n24181));
    defparam i19406_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14219_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n14410), .I3(GND_net), .O(n19008));   // verilog/coms.v(127[12] 300[6])
    defparam i14219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14220_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n14410), .I3(GND_net), .O(n19009));   // verilog/coms.v(127[12] 300[6])
    defparam i14220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4942));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14221_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n14410), .I3(GND_net), .O(n19010));   // verilog/coms.v(127[12] 300[6])
    defparam i14221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14222_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n14410), .I3(GND_net), .O(n19011));   // verilog/coms.v(127[12] 300[6])
    defparam i14222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14223_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n14410), .I3(GND_net), .O(n19012));   // verilog/coms.v(127[12] 300[6])
    defparam i14223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14224_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n14410), .I3(GND_net), .O(n19013));   // verilog/coms.v(127[12] 300[6])
    defparam i14224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14225_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n14410), .I3(GND_net), .O(n19014));   // verilog/coms.v(127[12] 300[6])
    defparam i14225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14226_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n14410), .I3(GND_net), .O(n19015));   // verilog/coms.v(127[12] 300[6])
    defparam i14226_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14227_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n14410), .I3(GND_net), .O(n19016));   // verilog/coms.v(127[12] 300[6])
    defparam i14227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n754), .I1(n24181), .I2(n756), .I3(n757), 
            .O(n4_adj_5031));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'ha8a0;
    SB_LUT4 i14228_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n14410), .I3(GND_net), .O(n19017));   // verilog/coms.v(127[12] 300[6])
    defparam i14228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14229_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n14410), .I3(GND_net), .O(n19018));   // verilog/coms.v(127[12] 300[6])
    defparam i14229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14230_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n14410), .I3(GND_net), .O(n19019));   // verilog/coms.v(127[12] 300[6])
    defparam i14230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4941));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14231_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n14410), .I3(GND_net), .O(n19020));   // verilog/coms.v(127[12] 300[6])
    defparam i14231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14232_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n14410), .I3(GND_net), .O(n19021));   // verilog/coms.v(127[12] 300[6])
    defparam i14232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14233_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n14410), .I3(GND_net), .O(n19022));   // verilog/coms.v(127[12] 300[6])
    defparam i14233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14234_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n14410), .I3(GND_net), .O(n19023));   // verilog/coms.v(127[12] 300[6])
    defparam i14234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14235_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n14410), .I3(GND_net), .O(n19024));   // verilog/coms.v(127[12] 300[6])
    defparam i14235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14236_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n14410), .I3(GND_net), .O(n19025));   // verilog/coms.v(127[12] 300[6])
    defparam i14236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14237_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n14410), .I3(GND_net), .O(n19026));   // verilog/coms.v(127[12] 300[6])
    defparam i14237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14238_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n14410), .I3(GND_net), .O(n19027));   // verilog/coms.v(127[12] 300[6])
    defparam i14238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14239_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n14410), .I3(GND_net), .O(n19028));   // verilog/coms.v(127[12] 300[6])
    defparam i14239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14240_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n14410), .I3(GND_net), .O(n19029));   // verilog/coms.v(127[12] 300[6])
    defparam i14240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14241_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n14410), .I3(GND_net), .O(n19030));   // verilog/coms.v(127[12] 300[6])
    defparam i14241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14242_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n14410), .I3(GND_net), .O(n19031));   // verilog/coms.v(127[12] 300[6])
    defparam i14242_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4940));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14243_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n14410), .I3(GND_net), .O(n19032));   // verilog/coms.v(127[12] 300[6])
    defparam i14243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14244_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n14410), .I3(GND_net), .O(n19033));   // verilog/coms.v(127[12] 300[6])
    defparam i14244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14245_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[22]), 
            .I2(n14410), .I3(GND_net), .O(n19034));   // verilog/coms.v(127[12] 300[6])
    defparam i14245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14246_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n14410), .I3(GND_net), .O(n19035));   // verilog/coms.v(127[12] 300[6])
    defparam i14246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14247_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[22]), 
            .I2(n14410), .I3(GND_net), .O(n19036));   // verilog/coms.v(127[12] 300[6])
    defparam i14247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14248_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n14410), .I3(GND_net), .O(n19037));   // verilog/coms.v(127[12] 300[6])
    defparam i14248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14249_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n14410), .I3(GND_net), .O(n19038));   // verilog/coms.v(127[12] 300[6])
    defparam i14249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14250_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n14410), .I3(GND_net), .O(n19039));   // verilog/coms.v(127[12] 300[6])
    defparam i14250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14251_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n14410), .I3(GND_net), .O(n19040));   // verilog/coms.v(127[12] 300[6])
    defparam i14251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14252_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n14410), .I3(GND_net), .O(n19041));   // verilog/coms.v(127[12] 300[6])
    defparam i14252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14253_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n14410), .I3(GND_net), .O(n19042));   // verilog/coms.v(127[12] 300[6])
    defparam i14253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14254_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n14410), .I3(GND_net), .O(n19043));   // verilog/coms.v(127[12] 300[6])
    defparam i14254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14255_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n14410), .I3(GND_net), .O(n19044));   // verilog/coms.v(127[12] 300[6])
    defparam i14255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14256_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n14410), .I3(GND_net), .O(n19045));   // verilog/coms.v(127[12] 300[6])
    defparam i14256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14257_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n14410), .I3(GND_net), .O(n19046));   // verilog/coms.v(127[12] 300[6])
    defparam i14257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14258_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n14410), .I3(GND_net), .O(n19047));   // verilog/coms.v(127[12] 300[6])
    defparam i14258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14259_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n14410), .I3(GND_net), .O(n19048));   // verilog/coms.v(127[12] 300[6])
    defparam i14259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14260_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n14410), .I3(GND_net), .O(n19049));   // verilog/coms.v(127[12] 300[6])
    defparam i14260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14261_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n14410), 
            .I3(GND_net), .O(n19050));   // verilog/coms.v(127[12] 300[6])
    defparam i14261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14262_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n14410), 
            .I3(GND_net), .O(n19051));   // verilog/coms.v(127[12] 300[6])
    defparam i14262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14263_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n14410), 
            .I3(GND_net), .O(n19052));   // verilog/coms.v(127[12] 300[6])
    defparam i14263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14264_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n14410), 
            .I3(GND_net), .O(n19053));   // verilog/coms.v(127[12] 300[6])
    defparam i14264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14265_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n14410), 
            .I3(GND_net), .O(n19054));   // verilog/coms.v(127[12] 300[6])
    defparam i14265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14266_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n14410), 
            .I3(GND_net), .O(n19055));   // verilog/coms.v(127[12] 300[6])
    defparam i14266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14267_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n14410), 
            .I3(GND_net), .O(n19056));   // verilog/coms.v(127[12] 300[6])
    defparam i14267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14268_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n14410), 
            .I3(GND_net), .O(n19057));   // verilog/coms.v(127[12] 300[6])
    defparam i14268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14269_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n34304), 
            .I3(GND_net), .O(n19058));   // verilog/coms.v(127[12] 300[6])
    defparam i14269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14270_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n34304), 
            .I3(GND_net), .O(n19059));   // verilog/coms.v(127[12] 300[6])
    defparam i14270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14271_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n34304), 
            .I3(GND_net), .O(n19060));   // verilog/coms.v(127[12] 300[6])
    defparam i14271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14272_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n34304), 
            .I3(GND_net), .O(n19061));   // verilog/coms.v(127[12] 300[6])
    defparam i14272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14273_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n34304), 
            .I3(GND_net), .O(n19062));   // verilog/coms.v(127[12] 300[6])
    defparam i14273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14274_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n34304), 
            .I3(GND_net), .O(n19063));   // verilog/coms.v(127[12] 300[6])
    defparam i14274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14275_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n34304), 
            .I3(GND_net), .O(n19064));   // verilog/coms.v(127[12] 300[6])
    defparam i14275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14276_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n34304), 
            .I3(GND_net), .O(n19065));   // verilog/coms.v(127[12] 300[6])
    defparam i14276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14277_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n34304), 
            .I3(GND_net), .O(n19066));   // verilog/coms.v(127[12] 300[6])
    defparam i14277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14278_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n34304), 
            .I3(GND_net), .O(n19067));   // verilog/coms.v(127[12] 300[6])
    defparam i14278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14279_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n34304), 
            .I3(GND_net), .O(n19068));   // verilog/coms.v(127[12] 300[6])
    defparam i14279_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4939));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30559_4_lut (.I0(n752), .I1(n755), .I2(n753), .I3(n4_adj_5031), 
            .O(n778));
    defparam i30559_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4938));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14280_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n34304), 
            .I3(GND_net), .O(n19069));   // verilog/coms.v(127[12] 300[6])
    defparam i14280_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14281_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n34304), 
            .I3(GND_net), .O(n19070));   // verilog/coms.v(127[12] 300[6])
    defparam i14281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14282_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n34304), 
            .I3(GND_net), .O(n19071));   // verilog/coms.v(127[12] 300[6])
    defparam i14282_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14283_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n34304), 
            .I3(GND_net), .O(n19072));   // verilog/coms.v(127[12] 300[6])
    defparam i14283_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14284_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n34304), 
            .I3(GND_net), .O(n19073));   // verilog/coms.v(127[12] 300[6])
    defparam i14284_3_lut.LUT_INIT = 16'hacac;
    EEPROM eeprom (.CLK_c(CLK_c), .GND_net(GND_net), .\state[3] (state_adj_5132[3]), 
           .n6(n6_adj_5055), .n3567({n3568}), .\state[1] (state_adj_5104[1]), 
           .\state[0] (state_adj_5104[0]), .enable_slow_N_3964(enable_slow_N_3964), 
           .n33160(n33160), .n32413(n32413), .read(read), .n23704(n23704), 
           .\state[2] (state_adj_5132[2]), .n7(n7_adj_5043), .n18643(n18643), 
           .rw(rw), .n32166(n32166), .data_ready(data_ready), .n32068(n32068), 
           .n32064(n32064), .n10(n10_adj_4926), .n17058(n17058), .n17053(n17053), 
           .n4867(n4867), .\saved_addr[0] (saved_addr[0]), .\state[0]_adj_13 (state_adj_5132[0]), 
           .\state_7__N_3861[0] (state_7__N_3861[0]), .n4(n4_adj_4927), 
           .n35900(n35900), .n4_adj_14(n4_adj_4865), .scl_enable(scl_enable), 
           .sda_enable(sda_enable), .\state_7__N_3877[3] (state_7__N_3877[3]), 
           .VCC_net(VCC_net), .scl(scl), .sda_out(sda_out), .n10_adj_15(n10_adj_4966), 
           .n5300(n5300), .n8(n8_adj_5030), .n18652(n18652), .data({data}), 
           .n18650(n18650), .n18649(n18649), .n18648(n18648), .n18647(n18647), 
           .n18646(n18646), .n19174(n19174), .n23726(n23726), .n18633(n18633), 
           .n18632(n18632)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(263[10] 274[6])
    SB_LUT4 i14285_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n34304), 
            .I3(GND_net), .O(n19074));   // verilog/coms.v(127[12] 300[6])
    defparam i14285_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14286_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n34304), 
            .I3(GND_net), .O(n19075));   // verilog/coms.v(127[12] 300[6])
    defparam i14286_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14287_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n34304), 
            .I3(GND_net), .O(n19076));   // verilog/coms.v(127[12] 300[6])
    defparam i14287_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14288_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n34304), 
            .I3(GND_net), .O(n19077));   // verilog/coms.v(127[12] 300[6])
    defparam i14288_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14289_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n34304), 
            .I3(GND_net), .O(n19078));   // verilog/coms.v(127[12] 300[6])
    defparam i14289_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14290_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n34304), 
            .I3(GND_net), .O(n19079));   // verilog/coms.v(127[12] 300[6])
    defparam i14290_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.clk32MHz(clk32MHz), .\data_in_frame[1] ({\data_in_frame[1] }), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .rx_data({rx_data}), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[25] ({\data_out_frame[25] }), 
         .\data_out_frame[24] ({\data_out_frame[24] }), .GND_net(GND_net), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .\data_out_frame[18] ({\data_out_frame[18] }), .n32658(n32658), 
         .\data_in_frame[19] ({\data_in_frame[19] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n30832(n30832), .n32385(n32385), .n32397(n32397), .n30803(n30803), 
         .n32722(n32722), .n32920(n32920), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n32699(n32699), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n32403(n32403), .n32412(n32412), .n66(n66), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[17] ({\data_in_frame[17] }), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .\data_in_frame[11] ({\data_in_frame[11] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .\data_in_frame[18] ({\data_in_frame[18] }), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n63(n63), .\FRAME_MATCHER.i_31__N_2461 (\FRAME_MATCHER.i_31__N_2461 ), 
         .n3303(n3303), .n4452(n4452), .n34405(n34405), .rx_data_ready(rx_data_ready), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .setpoint({setpoint}), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .n123(n123), .n1(n1_adj_4965), 
         .n18735(n18735), .n18734(n18734), .n18733(n18733), .n18732(n18732), 
         .n18731(n18731), .n18730(n18730), .n18729(n18729), .n18728(n18728), 
         .n18727(n18727), .n18726(n18726), .n18725(n18725), .n18724(n18724), 
         .n18723(n18723), .n18722(n18722), .n18721(n18721), .n18720(n18720), 
         .n18719(n18719), .n18718(n18718), .n18717(n18717), .n18716(n18716), 
         .n18715(n18715), .n18714(n18714), .n18713(n18713), .n18712(n18712), 
         .n18703(n18703), .n18702(n18702), .n18701(n18701), .n18700(n18700), 
         .n18699(n18699), .n18698(n18698), .n18697(n18697), .n18693(n18693), 
         .n18692(n18692), .control_mode({control_mode}), .n18691(n18691), 
         .n18690(n18690), .n18689(n18689), .n18688(n18688), .n18687(n18687), 
         .n18686(n18686), .\data_in[0] ({\data_in[0] }), .\data_in[1] ({\data_in[1] }), 
         .\data_in[2] ({\data_in[2] }), .\data_in[3] ({\data_in[3] }), .n18685(n18685), 
         .PWMLimit({PWMLimit}), .tx_active(tx_active), .\state[0] (state_adj_5132[0]), 
         .\state[2] (state_adj_5132[2]), .\state[3] (state_adj_5132[3]), 
         .n5300(n5300), .n32404(n32404), .n34118(n34118), .n34304(n34304), 
         .DE_c(DE_c), .n18684(n18684), .LED_c(LED_c), .n18683(n18683), 
         .n18682(n18682), .n18681(n18681), .n18680(n18680), .n18679(n18679), 
         .n18678(n18678), .ID({ID}), .n18677(n18677), .n18676(n18676), 
         .n18675(n18675), .n18674(n18674), .n18673(n18673), .n18672(n18672), 
         .n18671(n18671), .n18670(n18670), .n18669(n18669), .n18668(n18668), 
         .n18667(n18667), .n18666(n18666), .n18665(n18665), .n18664(n18664), 
         .n18663(n18663), .n37934(n37934), .n19173(n19173), .IntegralLimit({IntegralLimit}), 
         .n19172(n19172), .n19171(n19171), .n19170(n19170), .n19169(n19169), 
         .n19168(n19168), .n19167(n19167), .n19166(n19166), .n19165(n19165), 
         .n19164(n19164), .n19163(n19163), .n19162(n19162), .n19161(n19161), 
         .n19160(n19160), .n19159(n19159), .n19158(n19158), .n19157(n19157), 
         .n19156(n19156), .n19155(n19155), .n19154(n19154), .n19153(n19153), 
         .n19152(n19152), .n19151(n19151), .n19118(n19118), .n19117(n19117), 
         .n19116(n19116), .n19115(n19115), .n19114(n19114), .n19113(n19113), 
         .n19112(n19112), .n19111(n19111), .n19110(n19110), .n19109(n19109), 
         .n19108(n19108), .n19107(n19107), .n19106(n19106), .n19105(n19105), 
         .n19104(n19104), .n19103(n19103), .n19102(n19102), .n19101(n19101), 
         .n19100(n19100), .n19099(n19099), .n19098(n19098), .n19097(n19097), 
         .n19096(n19096), .n19095(n19095), .n19094(n19094), .n19093(n19093), 
         .n19092(n19092), .n19091(n19091), .n19090(n19090), .n19089(n19089), 
         .n19088(n19088), .n19087(n19087), .\Kp[1] (Kp[1]), .n19086(n19086), 
         .\Kp[2] (Kp[2]), .n19085(n19085), .\Kp[3] (Kp[3]), .n19084(n19084), 
         .\Kp[4] (Kp[4]), .n19083(n19083), .\Kp[5] (Kp[5]), .n19082(n19082), 
         .\Kp[6] (Kp[6]), .n19081(n19081), .\Kp[7] (Kp[7]), .n19080(n19080), 
         .\Kp[8] (Kp[8]), .n19079(n19079), .\Kp[9] (Kp[9]), .n19078(n19078), 
         .\Kp[10] (Kp[10]), .n19077(n19077), .\Kp[11] (Kp[11]), .n19076(n19076), 
         .\Kp[12] (Kp[12]), .n19075(n19075), .\Kp[13] (Kp[13]), .n19074(n19074), 
         .\Kp[14] (Kp[14]), .n19073(n19073), .\Kp[15] (Kp[15]), .n19072(n19072), 
         .\Ki[1] (Ki[1]), .n19071(n19071), .\Ki[2] (Ki[2]), .n19070(n19070), 
         .\Ki[3] (Ki[3]), .n19069(n19069), .\Ki[4] (Ki[4]), .n19068(n19068), 
         .\Ki[5] (Ki[5]), .n19067(n19067), .\Ki[6] (Ki[6]), .n19066(n19066), 
         .\Ki[7] (Ki[7]), .n19065(n19065), .\Ki[8] (Ki[8]), .n19064(n19064), 
         .\Ki[9] (Ki[9]), .n19063(n19063), .\Ki[10] (Ki[10]), .n19062(n19062), 
         .\Ki[11] (Ki[11]), .n19061(n19061), .\Ki[12] (Ki[12]), .n19060(n19060), 
         .\Ki[13] (Ki[13]), .n19059(n19059), .\Ki[14] (Ki[14]), .n19058(n19058), 
         .\Ki[15] (Ki[15]), .n19057(n19057), .n19056(n19056), .n19055(n19055), 
         .n19054(n19054), .n19053(n19053), .n19052(n19052), .n19051(n19051), 
         .n19050(n19050), .n19049(n19049), .n19048(n19048), .n19047(n19047), 
         .n19046(n19046), .n19045(n19045), .n19044(n19044), .n19043(n19043), 
         .n19042(n19042), .n19041(n19041), .n19040(n19040), .n19039(n19039), 
         .n19038(n19038), .n19037(n19037), .n19036(n19036), .n19035(n19035), 
         .n19034(n19034), .n19033(n19033), .n19032(n19032), .n19031(n19031), 
         .n19030(n19030), .n19029(n19029), .n19028(n19028), .n19027(n19027), 
         .n19026(n19026), .n19025(n19025), .n19024(n19024), .n19023(n19023), 
         .n19022(n19022), .n19021(n19021), .n19020(n19020), .n19019(n19019), 
         .n19018(n19018), .n19017(n19017), .n19016(n19016), .n19015(n19015), 
         .n19014(n19014), .n19013(n19013), .n19012(n19012), .n19011(n19011), 
         .n19010(n19010), .n19009(n19009), .n19008(n19008), .n19007(n19007), 
         .n19006(n19006), .n19005(n19005), .n19004(n19004), .n19003(n19003), 
         .n19002(n19002), .n19001(n19001), .n19000(n19000), .n18999(n18999), 
         .n18998(n18998), .n18997(n18997), .n18996(n18996), .n18994(n18994), 
         .n18993(n18993), .n18992(n18992), .n18991(n18991), .n18990(n18990), 
         .n18989(n18989), .n18988(n18988), .n18987(n18987), .n18986(n18986), 
         .n18985(n18985), .n18984(n18984), .n18983(n18983), .n18982(n18982), 
         .n32395(n32395), .n32400(n32400), .n18981(n18981), .n32409(n32409), 
         .n18980(n18980), .n18979(n18979), .n18978(n18978), .n18977(n18977), 
         .n18976(n18976), .n18975(n18975), .n18974(n18974), .n18973(n18973), 
         .n18972(n18972), .n18971(n18971), .n18970(n18970), .n18969(n18969), 
         .n18968(n18968), .n18967(n18967), .n18966(n18966), .n18965(n18965), 
         .n18964(n18964), .n18963(n18963), .n18962(n18962), .n18961(n18961), 
         .n18960(n18960), .n18959(n18959), .n18958(n18958), .n18957(n18957), 
         .n18956(n18956), .n18955(n18955), .n18954(n18954), .n18953(n18953), 
         .n18952(n18952), .n18951(n18951), .n18950(n18950), .n18949(n18949), 
         .n18948(n18948), .n18640(n18640), .n18639(n18639), .n18637(n18637), 
         .neopxl_color({neopxl_color}), .n18636(n18636), .\Ki[0] (Ki[0]), 
         .n18635(n18635), .\Kp[0] (Kp[0]), .n18634(n18634), .n18947(n18947), 
         .n18946(n18946), .n18945(n18945), .n18944(n18944), .n18943(n18943), 
         .n18942(n18942), .n18941(n18941), .n18940(n18940), .n18626(n18626), 
         .n18939(n18939), .n18938(n18938), .n18937(n18937), .n18936(n18936), 
         .n18935(n18935), .n18934(n18934), .n18933(n18933), .n18932(n18932), 
         .n18931(n18931), .n18930(n18930), .n18929(n18929), .n18928(n18928), 
         .n18927(n18927), .n18926(n18926), .n18925(n18925), .n18924(n18924), 
         .n18923(n18923), .n18922(n18922), .n18921(n18921), .n18920(n18920), 
         .n18919(n18919), .n18918(n18918), .n18917(n18917), .n18916(n18916), 
         .n18915(n18915), .n18914(n18914), .n18913(n18913), .n18912(n18912), 
         .n18911(n18911), .n18910(n18910), .n18909(n18909), .n18908(n18908), 
         .n18907(n18907), .n18906(n18906), .n18905(n18905), .n18904(n18904), 
         .n18903(n18903), .n18902(n18902), .n18901(n18901), .n18900(n18900), 
         .n18899(n18899), .n18898(n18898), .n18897(n18897), .n18896(n18896), 
         .n18895(n18895), .n18894(n18894), .n18893(n18893), .n18892(n18892), 
         .n18891(n18891), .n18890(n18890), .n18889(n18889), .n18888(n18888), 
         .n18887(n18887), .n18886(n18886), .n18885(n18885), .n18884(n18884), 
         .n18883(n18883), .n18882(n18882), .n18881(n18881), .n18880(n18880), 
         .n18879(n18879), .n18878(n18878), .n18877(n18877), .n18876(n18876), 
         .n18875(n18875), .n18874(n18874), .n18866(n18866), .n18865(n18865), 
         .n18864(n18864), .n18863(n18863), .n18862(n18862), .n18861(n18861), 
         .n18860(n18860), .n18859(n18859), .n18850(n18850), .n18849(n18849), 
         .n18848(n18848), .n18847(n18847), .n18846(n18846), .n18845(n18845), 
         .n18844(n18844), .n18843(n18843), .n18834(n18834), .n18833(n18833), 
         .n18832(n18832), .n18831(n18831), .n18830(n18830), .n18829(n18829), 
         .n18828(n18828), .n18827(n18827), .n18802(n18802), .n18801(n18801), 
         .n18800(n18800), .n18799(n18799), .n18798(n18798), .n18797(n18797), 
         .n18796(n18796), .n18795(n18795), .n18786(n18786), .n18785(n18785), 
         .n18784(n18784), .n18783(n18783), .n32831(n32831), .n18782(n18782), 
         .n18781(n18781), .n18780(n18780), .n18779(n18779), .n18770(n18770), 
         .n18769(n18769), .n18768(n18768), .n18767(n18767), .n18766(n18766), 
         .n18765(n18765), .n18764(n18764), .n18763(n18763), .n29929(n29929), 
         .n32394(n32394), .n32410(n32410), .n32402(n32402), .n14410(n14410), 
         .r_SM_Main({r_SM_Main_adj_5111}), .n10125(n10125), .tx_o(tx_o), 
         .\r_SM_Main_2__N_3450[1] (r_SM_Main_2__N_3450[1]), .\r_Bit_Index[0] (r_Bit_Index_adj_5113[0]), 
         .n18336(n18336), .n18590(n18590), .VCC_net(VCC_net), .n4(n4_adj_5053), 
         .n18644(n18644), .n18660(n18660), .n37939(n37939), .tx_enable(tx_enable), 
         .n23776(n23776), .n4_adj_3(n4_adj_4921), .\r_Bit_Index[0]_adj_4 (r_Bit_Index[0]), 
         .n17079(n17079), .n4_adj_5(n4), .r_SM_Main_adj_10({r_SM_Main}), 
         .\r_SM_Main_2__N_3379[2] (r_SM_Main_2__N_3379[2]), .n17084(n17084), 
         .n4_adj_9(n4_adj_4893), .n31970(n31970), .r_Rx_Data(r_Rx_Data), 
         .RX_N_10(RX_N_10), .n33211(n33211), .n33251(n33251), .n19204(n19204), 
         .n19202(n19202), .n19201(n19201), .n19200(n19200), .n19199(n19199), 
         .n19198(n19198), .n19197(n19197), .n18696(n18696), .n18995(n18995), 
         .n32359(n32359)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(137[8] 160[4])
    SB_LUT4 i14291_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n34304), 
            .I3(GND_net), .O(n19080));   // verilog/coms.v(127[12] 300[6])
    defparam i14291_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14292_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n34304), 
            .I3(GND_net), .O(n19081));   // verilog/coms.v(127[12] 300[6])
    defparam i14292_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14293_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n34304), 
            .I3(GND_net), .O(n19082));   // verilog/coms.v(127[12] 300[6])
    defparam i14293_3_lut.LUT_INIT = 16'hacac;
    pwm PWM (.n36611(n36611), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n16908(n16908), .pwm_counter({pwm_counter}), .n16906(n16906), 
        .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, clk32MHz, data_o, 
            GND_net, n34934, reg_B, VCC_net, ENCODER0_B_c_0, n18641, 
            n19175, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input clk32MHz;
    output [1:0]data_o;
    input GND_net;
    output n34934;
    output [1:0]reg_B;
    input VCC_net;
    input ENCODER0_B_c_0;
    input n18641;
    input n19175;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n3124;
    
    wire count_enable, B_delayed, A_delayed, count_direction, n3120, 
        n27846, n27845, n27844, n27843, n27842, n27841, n27840, 
        n27839, n27838, n27837, n27836, n27835, n27834, n27833, 
        n27832, n27831, n27830, n27829, n27828, n27827, n27826, 
        n27825, n27824, n27823;
    
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n3124[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_729_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n3120), 
            .I3(n27846), .O(n3124[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_729_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n3120), 
            .I3(n27845), .O(n3124[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_24 (.CI(n27845), .I0(encoder0_position[22]), .I1(n3120), 
            .CO(n27846));
    SB_LUT4 add_729_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n3120), 
            .I3(n27844), .O(n3124[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_23 (.CI(n27844), .I0(encoder0_position[21]), .I1(n3120), 
            .CO(n27845));
    SB_LUT4 add_729_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n3120), 
            .I3(n27843), .O(n3124[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_22 (.CI(n27843), .I0(encoder0_position[20]), .I1(n3120), 
            .CO(n27844));
    SB_LUT4 add_729_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n3120), 
            .I3(n27842), .O(n3124[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_21 (.CI(n27842), .I0(encoder0_position[19]), .I1(n3120), 
            .CO(n27843));
    SB_LUT4 add_729_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n3120), 
            .I3(n27841), .O(n3124[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_20 (.CI(n27841), .I0(encoder0_position[18]), .I1(n3120), 
            .CO(n27842));
    SB_LUT4 add_729_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n3120), 
            .I3(n27840), .O(n3124[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_19 (.CI(n27840), .I0(encoder0_position[17]), .I1(n3120), 
            .CO(n27841));
    SB_LUT4 add_729_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n3120), 
            .I3(n27839), .O(n3124[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_729_18 (.CI(n27839), .I0(encoder0_position[16]), .I1(n3120), 
            .CO(n27840));
    SB_LUT4 add_729_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n3120), 
            .I3(n27838), .O(n3124[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_17 (.CI(n27838), .I0(encoder0_position[15]), .I1(n3120), 
            .CO(n27839));
    SB_LUT4 add_729_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n3120), 
            .I3(n27837), .O(n3124[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_16 (.CI(n27837), .I0(encoder0_position[14]), .I1(n3120), 
            .CO(n27838));
    SB_LUT4 add_729_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n3120), 
            .I3(n27836), .O(n3124[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_15 (.CI(n27836), .I0(encoder0_position[13]), .I1(n3120), 
            .CO(n27837));
    SB_LUT4 add_729_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n3120), 
            .I3(n27835), .O(n3124[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_14 (.CI(n27835), .I0(encoder0_position[12]), .I1(n3120), 
            .CO(n27836));
    SB_LUT4 add_729_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n3120), 
            .I3(n27834), .O(n3124[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_13 (.CI(n27834), .I0(encoder0_position[11]), .I1(n3120), 
            .CO(n27835));
    SB_LUT4 add_729_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n3120), 
            .I3(n27833), .O(n3124[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_12 (.CI(n27833), .I0(encoder0_position[10]), .I1(n3120), 
            .CO(n27834));
    SB_LUT4 add_729_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n3120), 
            .I3(n27832), .O(n3124[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_11 (.CI(n27832), .I0(encoder0_position[9]), .I1(n3120), 
            .CO(n27833));
    SB_LUT4 add_729_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n3120), 
            .I3(n27831), .O(n3124[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_10 (.CI(n27831), .I0(encoder0_position[8]), .I1(n3120), 
            .CO(n27832));
    SB_LUT4 add_729_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n3120), 
            .I3(n27830), .O(n3124[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_9 (.CI(n27830), .I0(encoder0_position[7]), .I1(n3120), 
            .CO(n27831));
    SB_LUT4 add_729_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n3120), 
            .I3(n27829), .O(n3124[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_8 (.CI(n27829), .I0(encoder0_position[6]), .I1(n3120), 
            .CO(n27830));
    SB_LUT4 add_729_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n3120), 
            .I3(n27828), .O(n3124[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_7 (.CI(n27828), .I0(encoder0_position[5]), .I1(n3120), 
            .CO(n27829));
    SB_LUT4 add_729_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n3120), 
            .I3(n27827), .O(n3124[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_6 (.CI(n27827), .I0(encoder0_position[4]), .I1(n3120), 
            .CO(n27828));
    SB_LUT4 add_729_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n3120), 
            .I3(n27826), .O(n3124[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_5 (.CI(n27826), .I0(encoder0_position[3]), .I1(n3120), 
            .CO(n27827));
    SB_LUT4 add_729_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n3120), 
            .I3(n27825), .O(n3124[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_4 (.CI(n27825), .I0(encoder0_position[2]), .I1(n3120), 
            .CO(n27826));
    SB_LUT4 add_729_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n3120), 
            .I3(n27824), .O(n3124[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_3 (.CI(n27824), .I0(encoder0_position[1]), .I1(n3120), 
            .CO(n27825));
    SB_LUT4 add_729_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n27823), .O(n3124[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_729_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_729_2 (.CI(n27823), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n27824));
    SB_CARRY add_729_1 (.CI(GND_net), .I0(n3120), .I1(n3120), .CO(n27823));
    SB_LUT4 i1161_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n3120));   // quad.v(37[5] 40[8])
    defparam i1161_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,100)_U0  debounce (.n34934(n34934), .reg_B({reg_B}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .ENCODER0_B_c_0(ENCODER0_B_c_0), .n18641(n18641), .data_o({data_o}), 
            .n19175(n19175), .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (n34934, reg_B, GND_net, clk32MHz, 
            VCC_net, ENCODER0_B_c_0, n18641, data_o, n19175, ENCODER0_A_c_1);
    output n34934;
    output [1:0]reg_B;
    input GND_net;
    input clk32MHz;
    input VCC_net;
    input ENCODER0_B_c_0;
    input n18641;
    output [1:0]data_o;
    input n19175;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3693;
    wire [6:0]n33;
    
    wire n28434, n28433, n28432, n28431, n28430, n28429;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[4]), .I3(cnt_reg[2]), 
            .O(n34934));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n34934), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1550_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n28434), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1550_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1550_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n28433), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1550_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1550_add_4_7 (.CI(n28433), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n28434));
    SB_LUT4 cnt_reg_1550_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n28432), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1550_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1550_add_4_6 (.CI(n28432), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n28433));
    SB_LUT4 cnt_reg_1550_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n28431), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1550_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1550_add_4_5 (.CI(n28431), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n28432));
    SB_LUT4 cnt_reg_1550_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n28430), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1550_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1550_add_4_4 (.CI(n28430), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n28431));
    SB_LUT4 cnt_reg_1550_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n28429), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1550_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1550_add_4_3 (.CI(n28429), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n28430));
    SB_LUT4 cnt_reg_1550_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1550_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1550_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n28429));
    SB_DFFSR cnt_reg_1550__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n18641));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n19175));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1550__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1550__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1550__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1550__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1550__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1550__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (GND_net, \neo_pixel_transmitter.t0 , \neo_pixel_transmitter.done , 
            clk32MHz, VCC_net, n6, n33407, \state[0] , \state[1] , 
            start, n5, n2134, timer, n4, n26386, LED_c, neopxl_color, 
            n31374, n19149, n19148, n19147, n19146, n19145, n19144, 
            n19143, n19142, n19141, n19140, n19139, n19138, n19137, 
            n19136, n19135, n19134, n19133, n19132, n19131, n19130, 
            n19129, n19128, n19127, n19126, n19125, n19124, n19123, 
            n19122, n19121, n19120, n19119, NEOPXL_c, n18625) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    input VCC_net;
    output n6;
    output n33407;
    output \state[0] ;
    output \state[1] ;
    output start;
    output n5;
    output n2134;
    output [31:0]timer;
    output n4;
    output n26386;
    input LED_c;
    input [23:0]neopxl_color;
    input n31374;
    input n19149;
    input n19148;
    input n19147;
    input n19146;
    input n19145;
    input n19144;
    input n19143;
    input n19142;
    input n19141;
    input n19140;
    input n19139;
    input n19138;
    input n19137;
    input n19136;
    input n19135;
    input n19134;
    input n19133;
    input n19132;
    input n19131;
    input n19130;
    input n19129;
    input n19128;
    input n19127;
    input n19126;
    input n19125;
    input n19124;
    input n19123;
    input n19122;
    input n19121;
    input n19120;
    input n19119;
    output NEOPXL_c;
    input n18625;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n2500, n2401, n2423, n28586, n1806, n1803, n1798, n1805, 
        n24, n28587, n1808, n1804, n1802, n1807, n22, n1800, 
        n1799, n1797, n1801, n23, n1796;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n1809, n21, n1829, n1730, n37309;
    wire [31:0]n56;
    
    wire n2501, n2402, n28585, n1998, n2004, n18, n2003, n1999, 
        n1996, n2007, n28, n1997, n2005, n2000, n2002, n26, 
        n2502, n2403, n28584, n2001, n2008, n1994, n1995, n27, 
        n2503, n2404, n28583, n2006, n2009, n25, n2027, n2504, 
        n2405, n28582, \neo_pixel_transmitter.done_N_573 , n32362, n2505, 
        n2406, n28581, n2506, n2407, n28580, n1699, n1709, n17, 
        n1698, n1707, n1703, n1705, n21_adj_4709, n1704, n1701, 
        n1708, n20, n2507, n2408, n28579, n1702, n1697, n24_adj_4710, 
        n1700, n1706, n2693, n2704, n28_adj_4711, n2699, n2706, 
        n2694, n2691, n38, n2709, n24514, n2701, n2696, n2697, 
        n36, n2700, n2705, n42, n2702, n2690, n2689, n2708, 
        n40, n2687, n2703, n2695, n41, n2688, n2698, n2692, 
        n2707, n39, n2720, n1631, n37307, n2508, n2409, n37298, 
        n28578, n2509;
    wire [31:0]n255;
    
    wire n18162, n18520, n34978, n2588, n2489, n2522, n28577, 
        n2589, n2490, n28576, n2590, n2491, n28575, n2591, n2492, 
        n28574, n2592, n2493, n28573, n2593, n2494, n28572, n28646, 
        n2204, n2225, n28647, n2304, n2205, n28645, n2305, n2206, 
        n28644, n2594, n2495, n28571, n2595, n2496, n28570, n2596, 
        n2497, n28569, n2306, n2207, n28643, n2597, n2498, n28568, 
        n2307, n2208, n28642, n2308, n2209, n37300, n28641, n2598, 
        n2499, n28567, n27671, n27672, n2599, n28566, n27861, 
        n27862, n25_adj_4714, n27860;
    wire [31:0]one_wire_N_516;
    
    wire n2600, n28565, n2601, n28564, n2602, n28563, n1608, n1606, 
        n1604, n1603, n20_adj_4717, n1602, n1609, n13, n1598, 
        n1600, n18_adj_4718, n1605, n1599, n22_adj_4719, n1601, 
        n1607, n1532, n37306, n1334, n37304, n1506, n1503, n1500, 
        n1501, n18_adj_4722, n1504, n1502, n1499, n20_adj_4723, 
        n1505, n1509, n15, n1508, n1507, n1136, n37305, n2324, 
        n37302, n1109, n24484, n1105, n1103, n1108, n12, n1107, 
        n1106, n1104, n1037, n37303, n2;
    wire [31:0]n971;
    
    wire n1007, n2621, n37301, n1006, n27670, n24_adj_4726, n27859, 
        n2603, n28562, n2604, n28561, n2605, n28560, n2606, n28559, 
        n2309, n2607, n28558, n2608, n37299, n28557, n2609, n28556, 
        n27_adj_4728, n27858, n28555, n28554, n2390, n2291, n28640, 
        n2391, n2292, n28639, n28553, n28552, n2392, n2293, n28638, 
        n28551, n28550, n28549, n28548, n28547, n28546, n28545, 
        n28544, n2393, n2294, n28637, n28543, n28542, n2394, n2295, 
        n28636, n28541, n33146, n4_adj_4730, n28769, n2395, n2296, 
        n28635, n28540, n21_adj_4731, n23_adj_4732, n22_adj_4733, 
        n36_adj_4734, n26_adj_4735, n28_adj_4736, n37, n29_adj_4737, 
        n30_adj_4738, n17063, n1400, n1301, n28030, n9, n7, n8, 
        n1, n1005, n28768, n2396, n2297, n28634, n28539, n2397, 
        n2298, n28633, n28538, n1928, n37313, n28537, n28536, 
        n33550, n2398, n2299, n28632, n26370, n2399, n2300, n28631, 
        n2400, n2301, n28630, n2302, n28629, n28767, n2907, n2909, 
        n33_adj_4739, n2900, n2891, n2897, n2888, n41_adj_4740, 
        n2906, n2887, n2892, n38_adj_4741, n1401, n1302, n28029, 
        n28535, n28766, n2896, n2885, n2905, n2902, n43, n2899, 
        n2890, n2898, n2908, n40_adj_4742, n27857, n2303, n28628, 
        n2889, n2901, n46, n2886, n2894, n2895, n2903, n39_adj_4743, 
        n2904, n2893, n47, n1008, n28765, n2918, n28627;
    wire [31:0]n133;
    
    wire n28534, n28533, n28626, n26341, n1009, n28764, n28625, 
        n28532, n1402, n1303, n28028, n33_adj_4744, n28624, n1202, 
        n28763, n1403, n1304, n28027, n28531, n2819, n37314, n1433, 
        n37312, n28530, n28623, n1404, n1305, n28026, n28529, 
        n3209, n24526, n35871, n35, n11, n29_adj_4745, n51, n48, 
        n37_adj_4746, n23_adj_4747, n53, n39_adj_4748, n46_adj_4749, 
        n27_adj_4750, n57, n63, n43_adj_4751, n47_adj_4752, n25_adj_4753, 
        n33_adj_4754, n47_adj_4755, n61, n45, n59, n17_adj_4756, 
        n15_adj_4757, n55, n44, n28528, n31_adj_4758, n41_adj_4759, 
        n49, n43_adj_4760, n1405, n1306, n28025, n54, n45_adj_4761, 
        n13_adj_4762, n19_adj_4763, n21_adj_4764, n49_adj_4765, n29565, 
        n26387, n2798, n2804, n2791, n2795, n40_adj_4766, n28527, 
        n2796, n2793, n2788, n2808, n38_adj_4767, n2789, n2800, 
        n2803, n2805, n39_adj_4768, n27856, n2792, n2787, n2801, 
        n2799, n37_adj_4769, n10, n26337, n2786, n2797, n34, n1406, 
        n1307, n28024, n26348, n7_adj_4770, n38250, n28622, n2794, 
        n2806, n2807, n2790, n42_adj_4771, n46_adj_4772;
    wire [4:0]color_bit_N_559;
    
    wire n2802, n2809, n33_adj_4773, n1203, n28762, n37541, n37427, 
        n22_adj_4774, n37337, color_bit, n28526, n1204, n28761, 
        n1205, n28760, n28525, n1206, n28759, n28524, n1207, n28758, 
        n1208, n28757, n28523, n28522, n1209, n28756, n28755, 
        n28521, n28520, n28519, n1407, n1308, n28023, n27855, 
        n28518, n28754, n1895, n1902, n1899, n1897, n26_adj_4775, 
        n1907, n1909, n19_adj_4776, n1908, n1900, n16, n28517, 
        n1904, n1901, n1906, n1898, n24_adj_4777, n1905, n1903, 
        n28_adj_4778, n28516, n1896, n37311, n28515, n28514, n1408, 
        n1309, n28022, n28513, n28753, n28512, n28511, n28510, 
        n28509, n28508, n28507, n28752, n28506, n1409, n28505, 
        n28504, n28751, n28750, n27854, n28749, n28748, n27669, 
        n28747, n28746, n27679, n27680, n28745, n28744, n27853, 
        n28743, n33241, n28742, n28741, n28740, n27852, n28739, 
        n28738, n27851, n10_adj_4779, n12_adj_4780, n16_adj_4781, 
        n906, n807, n60, n838, n739, n15594, n708, n33188, n24530, 
        n16_adj_4782, n17_adj_4783, n37308, n28737, n28736, n27678, 
        n27850, n28735, n28734, n28597, n28457, n28596, n28456, 
        n28595, n28455, n28454, n28453, n28594, n28452, n28733, 
        n27677, n28593, n28732, n28592, n28731, n28451, n27668, 
        n28730, n28591, n27849, n28590, n28729, n28588, n28450, 
        n28728, n28449, n28727, n28726, n28725, n27848, n4_adj_4784, 
        n27847, n27676, n28724, n28448, n28447, n28723, n28446, 
        n28589, n28722, n28721, n28720, n28719, n28445, n28444, 
        n28718, n28443, n28442, n608, n7966, n29899, n33158, n15590, 
        n905, n4_adj_4786, n18398, n33247, n28441, n28440, n46_adj_4787, 
        n44_adj_4788, n45_adj_4789, n43_adj_4790, n42_adj_4791, n28717, 
        n28439, n28438, n41_adj_4792, n28437, n52, n47_adj_4793, 
        n28716, n28436, n14682, n6_adj_4794, n35911, n28435, n28715, 
        n28008, n27784, n28714, n28713, n28712, n28711, n28710, 
        n28709, n28708, n28707, n28706, n28007, n28705, n28704, 
        n28703, n28006, n28702, n28417, n28416, n28415, n28414, 
        n28413, n28005, n28412, n28411, n28410, n28409, n28408, 
        n28407, n28406, n28405, n28404, n28004, n28701, n28403, 
        n28402, n28003, n28002, n28001, n28401, n27783, n28700, 
        n28400, n28699, n28399, n28698, n28000, n27999, n28398, 
        n28697, n28397, n35012, n6_adj_4797, n28696, n28396, n28395, 
        n28695, n28394, n2984, n28393, n28694, n2985, n28392, 
        n2986, n28391, n2987, n28390, n2988, n28389, n27782, n2989, 
        n28388, n2990, n28387, n2991, n28386, n2992, n28385, n28693, 
        n2993, n28384, n28692, n2994, n28383, n2995, n28382, n2996, 
        n28381, n27675, n2997, n28380, n1235, n37320, n2998, n28379, 
        n2999, n28378, n3000, n28377, n3001, n28376, n3002, n28375, 
        n3003, n28374, n27781, n2093, n28691, n2094, n28690, n3004, 
        n28373, n2095, n28689, n3005, n28372, n3006, n28371, n3007, 
        n28370, n2096, n28688, n2097, n28687, n2098, n28686, n3008, 
        n37315, n28369, n3009, n2099, n28685, n2100, n28684, n3083, 
        n3017, n28368, n3084, n28367, n27780, n3085, n28366, n3086, 
        n28365, n2101, n28683, n3087, n28364, n3088, n28363, n3089, 
        n28362, n3090, n28361, n3091, n28360, n2102, n28682, n22_adj_4799, 
        n30_adj_4800, n34_adj_4801, n32_adj_4802, n33_adj_4803, n31_adj_4804, 
        n3092, n28359, n2103, n28681, n27674, n3093, n28358, n27667, 
        n2104, n28680, n27673, n2105, n28679, n3094, n28357, n36_adj_4805, 
        n25_adj_4806, n34_adj_4807, n40_adj_4808, n38_adj_4809, n39_adj_4810, 
        n37_adj_4811, n3095, n28356, n3096, n28355, n3097, n28354, 
        n2106, n28678, n3098, n28353, n3099, n28352, n3100, n28351, 
        n3101, n28350, n3102, n28349, n3103, n28348, n2193, n2194, 
        n28_adj_4812, n2203, n32_adj_4813, n2201, n2192, n2196, 
        n30_adj_4814, n3104, n28347, n3105, n28346, n3106, n28345, 
        n3107, n28344, n3108, n37317, n28343, n3109, n2107, n28677, 
        n2108, n37316, n28676, n3116, n28342, n28341, n28340, 
        n28339, n2195, n2199, n31_adj_4815, n2202, n2197, n2198, 
        n2200, n29_adj_4816, n28338, n28337, n28336, n28335, n2109, 
        n28334, n28333, n28332, n28331, n24_adj_4817, n34_adj_4818, 
        n22_adj_4819, n38_adj_4820, n36_adj_4821, n37_adj_4822, n28330, 
        n28329, n28328, n28327, n27666, n2126, n28675, n28326, 
        n28325, n35_adj_4823, n28324, n28323, n28322, n28321, n28320, 
        n28319, n28318, n28317, n37318, n28316, n28674, n37538, 
        n14_adj_4824, n9_adj_4825, n37478, n35154, n37472, n35157, 
        n34915, n37460, n35163, n27696, n27695, n37424, n27694, 
        n28673, n27693, n27692, n28672, n28671, n28670, n27691, 
        n28669, n27690, n27689, n28668, n27688, n28667, n28666, 
        n27687, n27_adj_4826, n33_adj_4827, n28665;
    wire [3:0]state_3__N_365;
    
    wire n27686, n28664, n27685, n28663, n27684, n28662, n28661, 
        n28660, n32_adj_4830, n31_adj_4831, n35_adj_4832, n37_adj_4833, 
        n37319, n28659, n27877, n27876, n27875, n27874, n27683, 
        n28658, n28657, n27873, n27682, n28656, n27872, n28655, 
        \neo_pixel_transmitter.done_N_579 , n33275, n27871, n27681, 
        n28654, n27870, n28653, n27869, n26349, n11_adj_4842, n28652, 
        n27868, n28651, n27867, n28083, n28082, n28081, n28080, 
        n28079, n28078, n28077, n28650, n28076, n27866, n28649, 
        n27865, n28648, n27864, n27863, n36260, n36176, n33261, 
        n18_adj_4843, n24500, n30_adj_4844, n28_adj_4845, n29_adj_4846, 
        n27_adj_4847, n37_adj_4848, n45_adj_4849, n42_adj_4850, n32_adj_4851, 
        n44_adj_4852, n50, n48_adj_4853, n49_adj_4854, n47_adj_4855, 
        n37340, n36546, n37334, n40_adj_4856, n44_adj_4857, n42_adj_4858, 
        n43_adj_4859, n41_adj_4860, n38_adj_4861, n46_adj_4862, n50_adj_4863, 
        n37_adj_4864;
    
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n28586), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i10_4_lut (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_11 (.CI(n28586), .I0(n2401), .I1(n2423), .CO(n28587));
    SB_LUT4 i8_4_lut (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n21));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut (.I0(n21), .I1(n23), .I2(n22), .I3(n24), .O(n1829));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30914_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37309));
    defparam i30914_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n28585), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n28585), .I0(n2402), .I1(n2423), .CO(n28586));
    SB_LUT4 i2_2_lut (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1513 (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26));
    defparam i10_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n28584), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n28584), .I0(n2403), .I1(n2423), .CO(n28585));
    SB_LUT4 i11_4_lut (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n28583), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_4_lut_adj_1514 (.I0(bit_ctr[15]), .I1(n18), .I2(n2006), 
            .I3(n2009), .O(n25));
    defparam i9_4_lut_adj_1514.LUT_INIT = 16'hfefc;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n2027));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_8 (.CI(n28583), .I0(n2404), .I1(n2423), .CO(n28584));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n28582), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n28582), .I0(n2405), .I1(n2423), .CO(n28583));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n32362), .D(\neo_pixel_transmitter.done_N_573 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n28581), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n28581), .I0(n2406), .I1(n2423), .CO(n28582));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n28580), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), .I3(GND_net), 
            .O(n17));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1515 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4709));
    defparam i8_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1516 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20));
    defparam i7_3_lut_adj_1516.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_1674_5 (.CI(n28580), .I0(n2407), .I1(n2423), .CO(n28581));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n28579), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_1517 (.I0(n21_adj_4709), .I1(n17), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4710));
    defparam i11_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1518 (.I0(n1700), .I1(n24_adj_4710), .I2(n20), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_4 (.CI(n28579), .I0(n2408), .I1(n2423), .CO(n28580));
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4711));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1519 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38));
    defparam i15_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i19733_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n24514));
    defparam i19733_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1520 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n24514), 
            .O(n36));
    defparam i13_4_lut_adj_1520.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n2700), .I1(n38), .I2(n28_adj_4711), .I3(n2705), 
            .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n2687), .I1(n36), .I2(n2703), .I3(n2695), 
            .O(n41));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30912_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37307));
    defparam i30912_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n37298), 
            .I3(n28578), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n28578), .I0(n2409), .I1(n37298), .CO(n28579));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n37298), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n18162), 
            .D(n255[1]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n18162), 
            .D(n255[2]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n18162), 
            .D(n255[3]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n18162), 
            .D(n255[4]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n18162), 
            .D(n255[5]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n18162), 
            .D(n255[6]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n18162), 
            .D(n255[7]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n18162), 
            .D(n255[8]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n18162), 
            .D(n255[9]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n18162), 
            .D(n255[10]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n18162), 
            .D(n255[11]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n18162), 
            .D(n255[12]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n18162), 
            .D(n255[13]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n18162), 
            .D(n255[14]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n18162), 
            .D(n255[15]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n18162), 
            .D(n255[16]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n18162), 
            .D(n255[17]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n18162), 
            .D(n255[18]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n18162), 
            .D(n255[19]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n18162), 
            .D(n255[20]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n18162), 
            .D(n255[21]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n18162), 
            .D(n255[22]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i21610_4_lut (.I0(n6), .I1(n33407), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n34978));   // verilog/neopixel.v(16[20:25])
    defparam i21610_4_lut.LUT_INIT = 16'hacca;
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n18162), 
            .D(n255[23]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n18162), 
            .D(n255[24]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(start), .I2(n5), .I3(n34978), 
            .O(n2134));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_4_lut.LUT_INIT = 16'h5554;
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n18162), 
            .D(n255[25]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n37298), 
            .CO(n28578));
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n18162), 
            .D(n255[26]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n18162), 
            .D(n255[27]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n18162), 
            .D(n255[28]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n18162), 
            .D(n255[29]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n18162), 
            .D(n255[30]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n18162), 
            .D(n255[31]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n28577), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n28576), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n28576), .I0(n2490), .I1(n2522), .CO(n28577));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n28575), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n28575), .I0(n2491), .I1(n2522), .CO(n28576));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n28574), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n28574), .I0(n2492), .I1(n2522), .CO(n28575));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n28573), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n28573), .I0(n2493), .I1(n2522), .CO(n28574));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n28572), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n28646), .I0(n2204), .I1(n2225), .CO(n28647));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n28645), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n28572), .I0(n2494), .I1(n2522), .CO(n28573));
    SB_CARRY mod_5_add_1540_7 (.CI(n28645), .I0(n2205), .I1(n2225), .CO(n28646));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n28644), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n28571), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n28571), .I0(n2495), .I1(n2522), .CO(n28572));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n28570), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n28644), .I0(n2206), .I1(n2225), .CO(n28645));
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_16 (.CI(n28570), .I0(n2496), .I1(n2522), .CO(n28571));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n28569), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n28569), .I0(n2497), .I1(n2522), .CO(n28570));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n28643), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n28643), .I0(n2207), .I1(n2225), .CO(n28644));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n28568), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n28642), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n28642), .I0(n2208), .I1(n2225), .CO(n28643));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n37300), 
            .I3(n28641), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_14 (.CI(n28568), .I0(n2498), .I1(n2522), .CO(n28569));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n28567), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n27671), .I0(bit_ctr[6]), .I1(GND_net), .CO(n27672));
    SB_CARRY mod_5_add_1741_13 (.CI(n28567), .I0(n2499), .I1(n2522), .CO(n28568));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n28566), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n28566), .I0(n2500), .I1(n2522), .CO(n28567));
    SB_CARRY sub_14_add_2_17 (.CI(n27861), .I0(timer[15]), .I1(n56[15]), 
            .CO(n27862));
    SB_LUT4 sub_14_add_2_16_lut (.I0(one_wire_N_516[21]), .I1(timer[14]), 
            .I2(n56[14]), .I3(n27860), .O(n25_adj_4714)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n28565), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_16 (.CI(n27860), .I0(timer[14]), .I1(n56[14]), 
            .CO(n27861));
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_11 (.CI(n28565), .I0(n2501), .I1(n2522), .CO(n28566));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n28564), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n28564), .I0(n2502), .I1(n2522), .CO(n28565));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n28563), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1521 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4717));
    defparam i8_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), .I3(GND_net), 
            .O(n13));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4718));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1522 (.I0(n13), .I1(n20_adj_4717), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4719));
    defparam i10_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1523 (.I0(n1601), .I1(n22_adj_4719), .I2(n18_adj_4718), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i30911_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37306));
    defparam i30911_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30909_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37304));
    defparam i30909_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4722));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1524 (.I0(n1504), .I1(n18_adj_4722), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4723));
    defparam i9_4_lut_adj_1524.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1525 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15));
    defparam i4_3_lut_adj_1525.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1526 (.I0(n15), .I1(n20_adj_4723), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1526.LUT_INIT = 16'hfffe;
    SB_LUT4 i30910_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37305));
    defparam i30910_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30907_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37302));
    defparam i30907_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19703_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n24484));
    defparam i19703_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n24484), .I3(n1108), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1107), .I1(n12), .I2(n1106), .I3(n1104), 
            .O(n1136));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30908_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37303));
    defparam i30908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30525_2_lut (.I0(n2), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i30525_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i30906_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37301));
    defparam i30906_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30523_2_lut (.I0(n2), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i30523_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n27670), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_15_lut (.I0(one_wire_N_516[22]), .I1(timer[13]), 
            .I2(n56[13]), .I3(n27859), .O(n24_adj_4726)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1741_9 (.CI(n28563), .I0(n2503), .I1(n2522), .CO(n28564));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n28562), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n28562), .I0(n2504), .I1(n2522), .CO(n28563));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n28561), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n28561), .I0(n2505), .I1(n2522), .CO(n28562));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n28560), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n28560), .I0(n2506), .I1(n2522), .CO(n28561));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n28559), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n28559), .I0(n2507), .I1(n2522), .CO(n28560));
    SB_CARRY mod_5_add_1540_3 (.CI(n28641), .I0(n2209), .I1(n37300), .CO(n28642));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n37300), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n28558), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_4 (.CI(n28558), .I0(n2508), .I1(n2522), .CO(n28559));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n37299), 
            .I3(n28557), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_3 (.CI(n28557), .I0(n2509), .I1(n37299), .CO(n28558));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n37299), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n37299), 
            .CO(n28557));
    SB_CARRY sub_14_add_2_15 (.CI(n27859), .I0(timer[13]), .I1(n56[13]), 
            .CO(n27860));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n28556), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_516[17]), .I1(timer[12]), 
            .I2(n56[12]), .I3(n27858), .O(n27_adj_4728)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_516[2]), .I1(one_wire_N_516[4]), .I2(one_wire_N_516[3]), 
            .I3(GND_net), .O(n33407));   // verilog/neopixel.v(6[16:24])
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n28555), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n28555), .I0(n2589), .I1(n2621), .CO(n28556));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n28554), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n37300), 
            .CO(n28641));
    SB_CARRY mod_5_add_1808_22 (.CI(n28554), .I0(n2590), .I1(n2621), .CO(n28555));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n28640), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n28639), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n28639), .I0(n2292), .I1(n2324), .CO(n28640));
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n28553), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n28553), .I0(n2591), .I1(n2621), .CO(n28554));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n28552), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_20 (.CI(n28552), .I0(n2592), .I1(n2621), .CO(n28553));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n28638), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n28551), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n28551), .I0(n2593), .I1(n2621), .CO(n28552));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n28550), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n28550), .I0(n2594), .I1(n2621), .CO(n28551));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n28549), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n28549), .I0(n2595), .I1(n2621), .CO(n28550));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n28548), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n28548), .I0(n2596), .I1(n2621), .CO(n28549));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n28547), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n28547), .I0(n2597), .I1(n2621), .CO(n28548));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n28546), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n28546), .I0(n2598), .I1(n2621), .CO(n28547));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n28545), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n28545), .I0(n2599), .I1(n2621), .CO(n28546));
    SB_CARRY mod_5_add_1607_19 (.CI(n28638), .I0(n2293), .I1(n2324), .CO(n28639));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n28544), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n28544), .I0(n2600), .I1(n2621), .CO(n28545));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n28637), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n28543), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n28543), .I0(n2601), .I1(n2621), .CO(n28544));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n28542), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n28542), .I0(n2602), .I1(n2621), .CO(n28543));
    SB_CARRY mod_5_add_1607_18 (.CI(n28637), .I0(n2294), .I1(n2324), .CO(n28638));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n28636), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n28636), .I0(n2295), .I1(n2324), .CO(n28637));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n28541), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i26763_2_lut (.I0(\state[1] ), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n33146));
    defparam i26763_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1808_9 (.CI(n28541), .I0(n2603), .I1(n2621), .CO(n28542));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4730), .I1(n4_adj_4730), .I2(n1037), 
            .I3(n28769), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n28635), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n28540), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1527 (.I0(n21_adj_4731), .I1(n23_adj_4732), .I2(n22_adj_4733), 
            .I3(n24_adj_4726), .O(n36_adj_4734));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1527.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1528 (.I0(n25_adj_4714), .I1(n27_adj_4728), .I2(n26_adj_4735), 
            .I3(n28_adj_4736), .O(n37));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1808_8 (.CI(n28540), .I0(n2604), .I1(n2621), .CO(n28541));
    SB_LUT4 i19_4_lut_adj_1529 (.I0(n37), .I1(n29_adj_4737), .I2(n36_adj_4734), 
            .I3(n30_adj_4738), .O(n17063));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28030), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i5_3_lut (.I0(n9), .I1(n7), .I2(n8), .I3(GND_net), .O(n1));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_1607_16 (.CI(n28635), .I0(n2296), .I1(n2324), .CO(n28636));
    SB_CARRY sub_14_add_2_14 (.CI(n27858), .I0(timer[12]), .I1(n56[12]), 
            .CO(n27859));
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n28768), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n28768), .I0(n1005), .I1(n1037), .CO(n28769));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n28634), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n28634), .I0(n2297), .I1(n2324), .CO(n28635));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n28539), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n28633), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n28539), .I0(n2605), .I1(n2621), .CO(n28540));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n28538), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n28538), .I0(n2606), .I1(n2621), .CO(n28539));
    SB_CARRY mod_5_add_1607_14 (.CI(n28633), .I0(n2298), .I1(n2324), .CO(n28634));
    SB_LUT4 i30918_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37313));
    defparam i30918_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n28537), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n28537), .I0(n2607), .I1(n2621), .CO(n28538));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n28536), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_adj_1530 (.I0(n33550), .I1(one_wire_N_516[4]), .I2(one_wire_N_516[3]), 
            .I3(GND_net), .O(n6));   // verilog/neopixel.v(6[16:24])
    defparam i2_3_lut_adj_1530.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n28632), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n5), .I1(n6), .I2(GND_net), .I3(GND_net), 
            .O(n26370));   // verilog/neopixel.v(6[16:24])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1607_13 (.CI(n28632), .I0(n2299), .I1(n2324), .CO(n28633));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n28631), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n28631), .I0(n2300), .I1(n2324), .CO(n28632));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n28630), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n28630), .I0(n2301), .I1(n2324), .CO(n28631));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n28629), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n28767), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n28767), .I0(n1006), .I1(n1037), .CO(n28768));
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4739));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1531 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_4740));
    defparam i16_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_4741));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28029), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n28536), .I0(n2608), .I1(n2621), .CO(n28537));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n37301), 
            .I3(n28535), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n28766), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_3 (.CI(n28535), .I0(n2609), .I1(n37301), .CO(n28536));
    SB_LUT4 i18_4_lut_adj_1532 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43));
    defparam i18_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_736_5 (.CI(n28766), .I0(n1007), .I1(n1037), .CO(n28767));
    SB_LUT4 i15_4_lut_adj_1533 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_4742));
    defparam i15_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n56[11]), 
            .I3(n27857), .O(one_wire_N_516[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n28629), .I0(n2302), .I1(n2324), .CO(n28630));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n28628), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n37301), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i21_4_lut (.I0(n41_adj_4740), .I1(n33_adj_4739), .I2(n2889), 
            .I3(n2901), .O(n46));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39_adj_4743));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1534 (.I0(n43), .I1(n2904), .I2(n38_adj_4741), 
            .I3(n2893), .O(n47));
    defparam i22_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n28765), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_13 (.CI(n27857), .I0(timer[11]), .I1(n56[11]), 
            .CO(n27858));
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n37301), 
            .CO(n28535));
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39_adj_4743), .I2(n46), .I3(n40_adj_4742), 
            .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_736_4 (.CI(n28765), .I0(n1008), .I1(n1037), .CO(n28766));
    SB_CARRY mod_5_add_1607_9 (.CI(n28628), .I0(n2303), .I1(n2324), .CO(n28629));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n28627), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1544_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n28534), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_10 (.CI(n28029), .I0(n1302), .I1(n1334), .CO(n28030));
    SB_CARRY mod_5_add_1607_8 (.CI(n28627), .I0(n2304), .I1(n2324), .CO(n28628));
    SB_LUT4 timer_1544_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n28533), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n28626), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n28626), .I0(n2305), .I1(n2324), .CO(n28627));
    SB_LUT4 i1_2_lut_adj_1535 (.I0(n33407), .I1(n5), .I2(GND_net), .I3(GND_net), 
            .O(n26341));   // verilog/neopixel.v(6[16:24])
    defparam i1_2_lut_adj_1535.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n37303), 
            .I3(n28764), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n28625), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n28625), .I0(n2306), .I1(n2324), .CO(n28626));
    SB_CARRY timer_1544_add_4_32 (.CI(n28533), .I0(GND_net), .I1(timer[30]), 
            .CO(n28534));
    SB_CARRY mod_5_add_736_3 (.CI(n28764), .I0(n1009), .I1(n37303), .CO(n28765));
    SB_LUT4 timer_1544_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n28532), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28028), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n37303), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_4_lut_adj_1536 (.I0(n26341), .I1(n26370), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n33_adj_4744));
    defparam i1_4_lut_adj_1536.LUT_INIT = 16'h3553;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n37303), 
            .CO(n28764));
    SB_CARRY timer_1544_add_4_31 (.CI(n28532), .I0(GND_net), .I1(timer[29]), 
            .CO(n28533));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n28624), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n28624), .I0(n2307), .I1(n2324), .CO(n28625));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28763), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n28028), .I0(n1303), .I1(n1334), .CO(n28029));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28027), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1544_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n28531), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30919_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37314));
    defparam i30919_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30917_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37312));
    defparam i30917_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1544_add_4_30 (.CI(n28531), .I0(GND_net), .I1(timer[28]), 
            .CO(n28532));
    SB_LUT4 timer_1544_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n28530), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_8 (.CI(n28027), .I0(n1304), .I1(n1334), .CO(n28028));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n28623), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1544_add_4_29 (.CI(n28530), .I0(GND_net), .I1(timer[27]), 
            .CO(n28531));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28026), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1544_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n28529), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_4 (.CI(n28623), .I0(n2308), .I1(n2324), .CO(n28624));
    SB_CARRY timer_1544_add_4_28 (.CI(n28529), .I0(GND_net), .I1(timer[26]), 
            .CO(n28530));
    SB_CARRY mod_5_add_937_7 (.CI(n28026), .I0(n1305), .I1(n1334), .CO(n28027));
    SB_LUT4 i19745_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n24526));
    defparam i19745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29840_2_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n26386), 
            .I3(GND_net), .O(n35871));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29840_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i30400_2_lut (.I0(n33_adj_4744), .I1(n33146), .I2(GND_net), 
            .I3(GND_net), .O(n32362));
    defparam i30400_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n11), .I2(n29_adj_4745), .I3(n51), 
            .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1537 (.I0(n37_adj_4746), .I1(n23_adj_4747), .I2(n53), 
            .I3(n39_adj_4748), .O(n46_adj_4749));
    defparam i18_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1538 (.I0(n27_adj_4750), .I1(n57), .I2(n63), 
            .I3(n43_adj_4751), .O(n47_adj_4752));
    defparam i19_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1539 (.I0(n25_adj_4753), .I1(n33_adj_4754), .I2(n47_adj_4755), 
            .I3(n61), .O(n45));
    defparam i17_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1540 (.I0(n59), .I1(n17_adj_4756), .I2(n15_adj_4757), 
            .I3(n55), .O(n44));
    defparam i16_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1544_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n28528), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1541 (.I0(n31_adj_4758), .I1(n41_adj_4759), .I2(n49), 
            .I3(n24526), .O(n43_adj_4760));
    defparam i15_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28025), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47_adj_4752), .I2(n46_adj_4749), 
            .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1542 (.I0(n45_adj_4761), .I1(n13_adj_4762), .I2(n19_adj_4763), 
            .I3(n21_adj_4764), .O(n49_adj_4765));
    defparam i21_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4765), .I1(n54), .I2(n43_adj_4760), 
            .I3(n44), .O(n29565));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1543 (.I0(\neo_pixel_transmitter.done ), .I1(n26386), 
            .I2(GND_net), .I3(GND_net), .O(n26387));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_adj_1543.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1544 (.I0(n17063), .I1(one_wire_N_516[11]), .I2(one_wire_N_516[9]), 
            .I3(one_wire_N_516[10]), .O(n26386));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1544.LUT_INIT = 16'heeea;
    SB_LUT4 i16_4_lut_adj_1545 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4766));
    defparam i16_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1544_add_4_27 (.CI(n28528), .I0(GND_net), .I1(timer[25]), 
            .CO(n28529));
    SB_LUT4 timer_1544_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n28527), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_1546 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4767));
    defparam i14_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1547 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4768));
    defparam i15_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n56[10]), 
            .I3(n27856), .O(one_wire_N_516[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut_adj_1548 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4769));
    defparam i13_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_937_6 (.CI(n28025), .I0(n1306), .I1(n1334), .CO(n28026));
    SB_LUT4 i23_4_lut (.I0(n35871), .I1(n10), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n26337));   // verilog/neopixel.v(16[20:25])
    defparam i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28024), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut_adj_1549 (.I0(n26348), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(n26387), .O(n7_adj_4770));
    defparam i15_4_lut_adj_1549.LUT_INIT = 16'hfaca;
    SB_LUT4 i1_rep_288_2_lut (.I0(bit_ctr[3]), .I1(n29565), .I2(GND_net), 
            .I3(GND_net), .O(n38250));
    defparam i1_rep_288_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n37302), 
            .I3(n28622), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1544_add_4_26 (.CI(n28527), .I0(GND_net), .I1(timer[24]), 
            .CO(n28528));
    SB_LUT4 i18_4_lut_adj_1550 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4771));
    defparam i18_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1551 (.I0(n37_adj_4769), .I1(n39_adj_4768), .I2(n38_adj_4767), 
            .I3(n40_adj_4766), .O(n46_adj_4772));
    defparam i22_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2239_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n29565), 
            .I3(GND_net), .O(color_bit_N_559[4]));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2239_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4773));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28762), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i23_4_lut_adj_1552 (.I0(n33_adj_4773), .I1(n46_adj_4772), .I2(n42_adj_4771), 
            .I3(n34), .O(n2819));
    defparam i23_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_LUT4 i2011675_i1_3_lut (.I0(n37541), .I1(n37427), .I2(bit_ctr[2]), 
            .I3(GND_net), .O(n22_adj_4774));
    defparam i2011675_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 color_bit_I_0_i31_4_lut (.I0(n37337), .I1(n22_adj_4774), .I2(color_bit_N_559[4]), 
            .I3(n38250), .O(color_bit));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i31_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY mod_5_add_803_8 (.CI(n28762), .I0(n1104), .I1(n1136), .CO(n28763));
    SB_LUT4 timer_1544_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n28526), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28761), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n28761), .I0(n1105), .I1(n1136), .CO(n28762));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28760), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n28760), .I0(n1106), .I1(n1136), .CO(n28761));
    SB_CARRY mod_5_add_1607_3 (.CI(n28622), .I0(n2309), .I1(n37302), .CO(n28623));
    SB_CARRY timer_1544_add_4_25 (.CI(n28526), .I0(GND_net), .I1(timer[23]), 
            .CO(n28527));
    SB_LUT4 timer_1544_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n28525), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n37302), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n37302), 
            .CO(n28622));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28759), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n28759), .I0(n1107), .I1(n1136), .CO(n28760));
    SB_CARRY timer_1544_add_4_24 (.CI(n28525), .I0(GND_net), .I1(timer[22]), 
            .CO(n28526));
    SB_LUT4 timer_1544_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n28524), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_23 (.CI(n28524), .I0(GND_net), .I1(timer[21]), 
            .CO(n28525));
    SB_CARRY add_21_7 (.CI(n27670), .I0(bit_ctr[5]), .I1(GND_net), .CO(n27671));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28758), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n28758), .I0(n1108), .I1(n1136), .CO(n28759));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n37305), 
            .I3(n28757), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n28757), .I0(n1109), .I1(n37305), .CO(n28758));
    SB_LUT4 timer_1544_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n28523), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n27856), .I0(timer[10]), .I1(n56[10]), 
            .CO(n27857));
    SB_CARRY timer_1544_add_4_22 (.CI(n28523), .I0(GND_net), .I1(timer[20]), 
            .CO(n28524));
    SB_LUT4 timer_1544_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n28522), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n37305), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n37305), 
            .CO(n28757));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n28756), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1544_add_4_21 (.CI(n28522), .I0(GND_net), .I1(timer[19]), 
            .CO(n28523));
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n28755), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n28024), .I0(n1307), .I1(n1334), .CO(n28025));
    SB_LUT4 timer_1544_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n28521), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_20 (.CI(n28521), .I0(GND_net), .I1(timer[18]), 
            .CO(n28522));
    SB_LUT4 timer_1544_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n28520), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_19 (.CI(n28520), .I0(GND_net), .I1(timer[17]), 
            .CO(n28521));
    SB_LUT4 timer_1544_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n28519), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28023), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1544_add_4_18 (.CI(n28519), .I0(GND_net), .I1(timer[16]), 
            .CO(n28520));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n56[9]), 
            .I3(n27855), .O(one_wire_N_516[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_12 (.CI(n28755), .I0(n1500), .I1(n1532), .CO(n28756));
    SB_LUT4 timer_1544_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n28518), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_4 (.CI(n28023), .I0(n1308), .I1(n1334), .CO(n28024));
    SB_CARRY timer_1544_add_4_17 (.CI(n28518), .I0(GND_net), .I1(timer[15]), 
            .CO(n28519));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n28754), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_11 (.CI(n28754), .I0(n1501), .I1(n1532), .CO(n28755));
    SB_LUT4 i11_4_lut_adj_1553 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4775));
    defparam i11_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1554 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19_adj_4776));
    defparam i4_3_lut_adj_1554.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1555 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16));
    defparam i1_2_lut_adj_1555.LUT_INIT = 16'heeee;
    SB_LUT4 timer_1544_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n28517), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1556 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4777));
    defparam i9_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1544_add_4_16 (.CI(n28517), .I0(GND_net), .I1(timer[14]), 
            .CO(n28518));
    SB_LUT4 i13_4_lut_adj_1557 (.I0(n19_adj_4776), .I1(n26_adj_4775), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4778));
    defparam i13_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1544_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n28516), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_15 (.CI(n28516), .I0(GND_net), .I1(timer[13]), 
            .CO(n28517));
    SB_LUT4 i14_4_lut_adj_1558 (.I0(n1896), .I1(n28_adj_4778), .I2(n24_adj_4777), 
            .I3(n16), .O(n1928));
    defparam i14_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i30916_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37311));
    defparam i30916_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1544_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n28515), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_14 (.CI(n28515), .I0(GND_net), .I1(timer[12]), 
            .CO(n28516));
    SB_LUT4 timer_1544_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n28514), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_13 (.CI(n28514), .I0(GND_net), .I1(timer[11]), 
            .CO(n28515));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n37304), 
            .I3(n28022), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1544_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n28513), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_12 (.CI(n28513), .I0(GND_net), .I1(timer[10]), 
            .CO(n28514));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n28753), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1544_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n28512), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_11 (.CI(n28512), .I0(GND_net), .I1(timer[9]), 
            .CO(n28513));
    SB_LUT4 timer_1544_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n28511), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_3 (.CI(n28022), .I0(n1309), .I1(n37304), .CO(n28023));
    SB_CARRY sub_14_add_2_11 (.CI(n27855), .I0(timer[9]), .I1(n56[9]), 
            .CO(n27856));
    SB_CARRY timer_1544_add_4_10 (.CI(n28511), .I0(GND_net), .I1(timer[8]), 
            .CO(n28512));
    SB_LUT4 timer_1544_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n28510), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_9 (.CI(n28510), .I0(GND_net), .I1(timer[7]), 
            .CO(n28511));
    SB_LUT4 timer_1544_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n28509), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_8 (.CI(n28509), .I0(GND_net), .I1(timer[6]), 
            .CO(n28510));
    SB_LUT4 timer_1544_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n28508), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_7 (.CI(n28508), .I0(GND_net), .I1(timer[5]), 
            .CO(n28509));
    SB_LUT4 timer_1544_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n28507), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_10 (.CI(n28753), .I0(n1502), .I1(n1532), .CO(n28754));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n28752), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1544_add_4_6 (.CI(n28507), .I0(GND_net), .I1(timer[4]), 
            .CO(n28508));
    SB_CARRY mod_5_add_1071_9 (.CI(n28752), .I0(n1503), .I1(n1532), .CO(n28753));
    SB_LUT4 timer_1544_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n28506), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_5 (.CI(n28506), .I0(GND_net), .I1(timer[3]), 
            .CO(n28507));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n37304), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n37304), 
            .CO(n28022));
    SB_LUT4 timer_1544_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n28505), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_4 (.CI(n28505), .I0(GND_net), .I1(timer[2]), 
            .CO(n28506));
    SB_LUT4 timer_1544_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n28504), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_3 (.CI(n28504), .I0(GND_net), .I1(timer[1]), 
            .CO(n28505));
    SB_LUT4 timer_1544_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1544_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1544_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n28504));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n28751), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n28751), .I0(n1504), .I1(n1532), .CO(n28752));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n28750), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_10_lut (.I0(one_wire_N_516[11]), .I1(timer[8]), 
            .I2(n56[8]), .I3(n27854), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1071_7 (.CI(n28750), .I0(n1505), .I1(n1532), .CO(n28751));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n28749), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_10 (.CI(n27854), .I0(timer[8]), .I1(n56[8]), 
            .CO(n27855));
    SB_CARRY mod_5_add_1071_6 (.CI(n28749), .I0(n1506), .I1(n1532), .CO(n28750));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n28748), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n28748), .I0(n1507), .I1(n1532), .CO(n28749));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n27669), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n28747), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n28747), .I0(n1508), .I1(n1532), .CO(n28748));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n37306), 
            .I3(n28746), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_3 (.CI(n28746), .I0(n1509), .I1(n37306), .CO(n28747));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n37306), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n37306), 
            .CO(n28746));
    SB_CARRY add_21_16 (.CI(n27679), .I0(bit_ctr[14]), .I1(GND_net), .CO(n27680));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n28745), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n28744), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_9_lut (.I0(one_wire_N_516[10]), .I1(timer[7]), 
            .I2(n56[7]), .I3(n27853), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1138_13 (.CI(n28744), .I0(n1599), .I1(n1631), .CO(n28745));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n28743), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_4_lut (.I0(n17063), .I1(one_wire_N_516[9]), .I2(n6), 
            .I3(n1), .O(n33241));   // verilog/neopixel.v(53[15:25])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_9 (.CI(n27853), .I0(timer[7]), .I1(n56[7]), 
            .CO(n27854));
    SB_CARRY mod_5_add_1138_12 (.CI(n28743), .I0(n1600), .I1(n1631), .CO(n28744));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n28742), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n28742), .I0(n1601), .I1(n1631), .CO(n28743));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n28741), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_2_lut_3_lut (.I0(n17063), .I1(one_wire_N_516[9]), .I2(n1), 
            .I3(GND_net), .O(n5));   // verilog/neopixel.v(53[15:25])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_CARRY mod_5_add_1138_10 (.CI(n28741), .I0(n1602), .I1(n1631), .CO(n28742));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n28740), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n28740), .I0(n1603), .I1(n1631), .CO(n28741));
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_516[5]), .I1(timer[6]), .I2(n56[6]), 
            .I3(n27852), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n28739), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_8 (.CI(n27852), .I0(timer[6]), .I1(n56[6]), 
            .CO(n27853));
    SB_CARRY mod_5_add_1138_8 (.CI(n28739), .I0(n1604), .I1(n1631), .CO(n28740));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n28738), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n28738), .I0(n1605), .I1(n1631), .CO(n28739));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n56[5]), 
            .I3(n27851), .O(one_wire_N_516[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1559 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4779));
    defparam i1_2_lut_adj_1559.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12_adj_4780));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1560 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4779), 
            .O(n16_adj_4781));
    defparam i7_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1561 (.I0(n1307), .I1(n16_adj_4781), .I2(n12_adj_4780), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(bit_ctr[28]), .I1(n739), .I2(GND_net), 
            .I3(GND_net), .O(n15594));
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h6666;
    SB_LUT4 mod_5_i538_3_lut (.I0(n708), .I1(n33188), .I2(n739), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut.LUT_INIT = 16'ha9a9;
    SB_CARRY sub_14_add_2_7 (.CI(n27851), .I0(timer[5]), .I1(n56[5]), 
            .CO(n27852));
    SB_LUT4 i19749_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n24530));
    defparam i19749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1563 (.I0(n1405), .I1(n24530), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4782));
    defparam i6_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1564 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4783));
    defparam i7_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1565 (.I0(n17_adj_4783), .I1(n1408), .I2(n16_adj_4782), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i30913_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37308));
    defparam i30913_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n28737), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n28737), .I0(n1606), .I1(n1631), .CO(n28738));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n28736), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n27678), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n56[4]), 
            .I3(n27850), .O(one_wire_N_516[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_5 (.CI(n28736), .I0(n1607), .I1(n1631), .CO(n28737));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n28735), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n28735), .I0(n1608), .I1(n1631), .CO(n28736));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n37307), 
            .I3(n28734), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n28597), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i21657_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_573 ));   // verilog/neopixel.v(16[20:25])
    defparam i21657_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n28457), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n28596), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_3 (.CI(n28734), .I0(n1609), .I1(n37307), .CO(n28735));
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n28456), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n37307), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_21 (.CI(n28596), .I0(n2391), .I1(n2423), .CO(n28597));
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n37307), 
            .CO(n28734));
    SB_CARRY mod_5_add_1875_24 (.CI(n28456), .I0(n2688), .I1(n2720), .CO(n28457));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n28595), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n28455), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n28455), .I0(n2689), .I1(n2720), .CO(n28456));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n28454), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_22 (.CI(n28454), .I0(n2690), .I1(n2720), .CO(n28455));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n28453), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n28453), .I0(n2691), .I1(n2720), .CO(n28454));
    SB_CARRY mod_5_add_1674_20 (.CI(n28595), .I0(n2392), .I1(n2423), .CO(n28596));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n28594), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n28452), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n28594), .I0(n2393), .I1(n2423), .CO(n28595));
    SB_CARRY add_21_15 (.CI(n27678), .I0(bit_ctr[13]), .I1(GND_net), .CO(n27679));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n28733), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n27677), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n28593), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_20 (.CI(n28452), .I0(n2692), .I1(n2720), .CO(n28453));
    SB_CARRY mod_5_add_1674_18 (.CI(n28593), .I0(n2394), .I1(n2423), .CO(n28594));
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n28732), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n28732), .I0(n1698), .I1(n1730), .CO(n28733));
    SB_CARRY add_21_6 (.CI(n27669), .I0(bit_ctr[4]), .I1(GND_net), .CO(n27670));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n28592), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_6 (.CI(n27850), .I0(timer[4]), .I1(n56[4]), 
            .CO(n27851));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n28731), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n28731), .I0(n1699), .I1(n1730), .CO(n28732));
    SB_CARRY mod_5_add_1674_17 (.CI(n28592), .I0(n2395), .I1(n2423), .CO(n28593));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n28451), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n27668), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n28730), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_5 (.CI(n27668), .I0(bit_ctr[3]), .I1(GND_net), .CO(n27669));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n28591), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_14 (.CI(n27677), .I0(bit_ctr[12]), .I1(GND_net), .CO(n27678));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n56[3]), 
            .I3(n27849), .O(one_wire_N_516[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_12 (.CI(n28730), .I0(n1700), .I1(n1730), .CO(n28731));
    SB_CARRY mod_5_add_1875_19 (.CI(n28451), .I0(n2693), .I1(n2720), .CO(n28452));
    SB_CARRY mod_5_add_1674_16 (.CI(n28591), .I0(n2396), .I1(n2423), .CO(n28592));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n28590), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n28729), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n28590), .I0(n2397), .I1(n2423), .CO(n28591));
    SB_CARRY mod_5_add_1674_12 (.CI(n28587), .I0(n2400), .I1(n2423), .CO(n28588));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n28450), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_18 (.CI(n28450), .I0(n2694), .I1(n2720), .CO(n28451));
    SB_CARRY mod_5_add_1205_11 (.CI(n28729), .I0(n1701), .I1(n1730), .CO(n28730));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n28728), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n28728), .I0(n1702), .I1(n1730), .CO(n28729));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n28449), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n28449), .I0(n2695), .I1(n2720), .CO(n28450));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n28727), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n28727), .I0(n1703), .I1(n1730), .CO(n28728));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n28726), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n28726), .I0(n1704), .I1(n1730), .CO(n28727));
    SB_CARRY sub_14_add_2_5 (.CI(n27849), .I0(timer[3]), .I1(n56[3]), 
            .CO(n27850));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n28725), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n56[2]), 
            .I3(n27848), .O(one_wire_N_516[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n27848), .I0(timer[2]), .I1(n56[2]), 
            .CO(n27849));
    SB_CARRY mod_5_add_1205_7 (.CI(n28725), .I0(n1705), .I1(n1730), .CO(n28726));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_516[2]), .I1(timer[1]), .I2(n56[1]), 
            .I3(n27847), .O(n4_adj_4784)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n27676), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_3 (.CI(n27847), .I0(timer[1]), .I1(n56[1]), 
            .CO(n27848));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n28724), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n28448), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_2_lut (.I0(n4_adj_4784), .I1(timer[0]), .I2(n56[0]), 
            .I3(VCC_net), .O(n33550)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1875_16 (.CI(n28448), .I0(n2696), .I1(n2720), .CO(n28449));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n28447), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n28724), .I0(n1706), .I1(n1730), .CO(n28725));
    SB_CARRY mod_5_add_1875_15 (.CI(n28447), .I0(n2697), .I1(n2720), .CO(n28448));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n28723), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n28723), .I0(n1707), .I1(n1730), .CO(n28724));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n28446), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n56[0]), 
            .CO(n27847));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n28587), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n28588), .I0(n2399), .I1(n2423), .CO(n28589));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n28588), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n28722), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n28722), .I0(n1708), .I1(n1730), .CO(n28723));
    SB_CARRY mod_5_add_1674_14 (.CI(n28589), .I0(n2398), .I1(n2423), .CO(n28590));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n28589), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n28446), .I0(n2698), .I1(n2720), .CO(n28447));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n37309), 
            .I3(n28721), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n28721), .I0(n1709), .I1(n37309), .CO(n28722));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n37309), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n37309), 
            .CO(n28721));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n28720), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n28719), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n28445), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n28719), .I0(n1797), .I1(n1829), .CO(n28720));
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1875_13 (.CI(n28445), .I0(n2699), .I1(n2720), .CO(n28446));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n28444), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n28444), .I0(n2700), .I1(n2720), .CO(n28445));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n28718), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i24_4_lut_adj_1566 (.I0(start), .I1(n26370), .I2(\state[0] ), 
            .I3(n26341), .O(n10));   // verilog/neopixel.v(16[20:25])
    defparam i24_4_lut_adj_1566.LUT_INIT = 16'h4540;
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n28443), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n28718), .I0(n1798), .I1(n1829), .CO(n28719));
    SB_CARRY mod_5_add_1875_11 (.CI(n28443), .I0(n2701), .I1(n2720), .CO(n28444));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n28442), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n28442), .I0(n2702), .I1(n2720), .CO(n28443));
    SB_LUT4 i1_2_lut_adj_1567 (.I0(\neo_pixel_transmitter.done ), .I1(n10), 
            .I2(GND_net), .I3(GND_net), .O(n26348));   // verilog/neopixel.v(16[20:25])
    defparam i1_2_lut_adj_1567.LUT_INIT = 16'h8888;
    SB_LUT4 i19636_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i19636_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n608), .I2(n33188), .I3(n7966), 
            .O(n739));
    defparam i2_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 i29731_3_lut (.I0(n29899), .I1(bit_ctr[28]), .I2(n739), .I3(GND_net), 
            .O(n33158));
    defparam i29731_3_lut.LUT_INIT = 16'ha6a6;
    SB_LUT4 i1_2_lut_adj_1568 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n15590));
    defparam i1_2_lut_adj_1568.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i1_3_lut_adj_1569 (.I0(n905), .I1(bit_ctr[26]), .I2(n15590), 
            .I3(GND_net), .O(n4_adj_4786));   // verilog/neopixel.v(22[26:36])
    defparam i1_3_lut_adj_1569.LUT_INIT = 16'h1515;
    SB_LUT4 i2_4_lut_adj_1570 (.I0(n18398), .I1(n906), .I2(n33247), .I3(n4_adj_4786), 
            .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i2_4_lut_adj_1570.LUT_INIT = 16'h0100;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n15590), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n28441), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n28441), .I0(n2703), .I1(n2720), .CO(n28442));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n28440), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n28440), .I0(n2704), .I1(n2720), .CO(n28441));
    SB_LUT4 i19_4_lut_adj_1571 (.I0(bit_ctr[23]), .I1(bit_ctr[16]), .I2(bit_ctr[20]), 
            .I3(bit_ctr[7]), .O(n46_adj_4787));   // verilog/neopixel.v(38[12:22])
    defparam i19_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1572 (.I0(bit_ctr[14]), .I1(bit_ctr[9]), .I2(bit_ctr[25]), 
            .I3(bit_ctr[10]), .O(n44_adj_4788));   // verilog/neopixel.v(38[12:22])
    defparam i17_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1573 (.I0(bit_ctr[27]), .I1(bit_ctr[12]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[29]), .O(n45_adj_4789));   // verilog/neopixel.v(38[12:22])
    defparam i18_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1574 (.I0(bit_ctr[6]), .I1(bit_ctr[31]), .I2(bit_ctr[19]), 
            .I3(bit_ctr[21]), .O(n43_adj_4790));   // verilog/neopixel.v(38[12:22])
    defparam i16_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1575 (.I0(bit_ctr[17]), .I1(bit_ctr[28]), .I2(bit_ctr[11]), 
            .I3(bit_ctr[5]), .O(n42_adj_4791));   // verilog/neopixel.v(38[12:22])
    defparam i15_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n28717), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n28439), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n28717), .I0(n1799), .I1(n1829), .CO(n28718));
    SB_CARRY mod_5_add_1875_7 (.CI(n28439), .I0(n2705), .I1(n2720), .CO(n28440));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n28438), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n28438), .I0(n2706), .I1(n2720), .CO(n28439));
    SB_LUT4 i14_3_lut (.I0(bit_ctr[26]), .I1(bit_ctr[13]), .I2(bit_ctr[22]), 
            .I3(GND_net), .O(n41_adj_4792));   // verilog/neopixel.v(38[12:22])
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n28437), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i25_4_lut (.I0(n43_adj_4790), .I1(n45_adj_4789), .I2(n44_adj_4788), 
            .I3(n46_adj_4787), .O(n52));   // verilog/neopixel.v(38[12:22])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_5 (.CI(n28437), .I0(n2707), .I1(n2720), .CO(n28438));
    SB_LUT4 i20_4_lut_adj_1576 (.I0(bit_ctr[30]), .I1(bit_ctr[18]), .I2(bit_ctr[24]), 
            .I3(bit_ctr[8]), .O(n47_adj_4793));   // verilog/neopixel.v(38[12:22])
    defparam i20_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n28716), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n28436), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n28716), .I0(n1800), .I1(n1829), .CO(n28717));
    SB_LUT4 i26_4_lut_adj_1577 (.I0(n47_adj_4793), .I1(n52), .I2(n41_adj_4792), 
            .I3(n42_adj_4791), .O(n14682));   // verilog/neopixel.v(38[12:22])
    defparam i26_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1578 (.I0(start), .I1(n26341), .I2(\state[1] ), 
            .I3(\state[0] ), .O(n6_adj_4794));   // verilog/neopixel.v(16[20:25])
    defparam i2_4_lut_adj_1578.LUT_INIT = 16'h0544;
    SB_LUT4 i13760_4_lut (.I0(n18162), .I1(\neo_pixel_transmitter.done ), 
            .I2(n6_adj_4794), .I3(n26370), .O(n18520));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13760_4_lut.LUT_INIT = 16'h2aaa;
    SB_LUT4 i21603_4_lut (.I0(n26348), .I1(n35911), .I2(\state[1] ), .I3(\state[0] ), 
            .O(n18162));   // verilog/neopixel.v(16[20:25])
    defparam i21603_4_lut.LUT_INIT = 16'hca0a;
    SB_CARRY mod_5_add_1875_4 (.CI(n28436), .I0(n2708), .I1(n2720), .CO(n28437));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n37308), 
            .I3(n28435), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n28715), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_3 (.CI(n28435), .I0(n2709), .I1(n37308), .CO(n28436));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n37308), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n37308), 
            .CO(n28435));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n28008), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_13 (.CI(n27676), .I0(bit_ctr[11]), .I1(GND_net), .CO(n27677));
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n27784), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1272_11 (.CI(n28715), .I0(n1801), .I1(n1829), .CO(n28716));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n28714), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n28714), .I0(n1802), .I1(n1829), .CO(n28715));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n28713), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n28713), .I0(n1803), .I1(n1829), .CO(n28714));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n28712), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n28712), .I0(n1804), .I1(n1829), .CO(n28713));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n28711), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n28711), .I0(n1805), .I1(n1829), .CO(n28712));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n28710), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n28710), .I0(n1806), .I1(n1829), .CO(n28711));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n28709), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n28709), .I0(n1807), .I1(n1829), .CO(n28710));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n28708), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n28708), .I0(n1808), .I1(n1829), .CO(n28709));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n37311), 
            .I3(n28707), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n28707), .I0(n1809), .I1(n37311), .CO(n28708));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n37311), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n37311), 
            .CO(n28707));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n28706), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n28007), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n28007), .I0(n1401), .I1(n1433), .CO(n28008));
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n28705), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n28705), .I0(n1896), .I1(n1928), .CO(n28706));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n28704), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n28704), .I0(n1897), .I1(n1928), .CO(n28705));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n28703), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n28703), .I0(n1898), .I1(n1928), .CO(n28704));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n28006), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n28702), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n28702), .I0(n1899), .I1(n1928), .CO(n28703));
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n28417), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n28416), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n28416), .I0(n2787), .I1(n2819), .CO(n28417));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n28415), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n28415), .I0(n2788), .I1(n2819), .CO(n28416));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n28414), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n28414), .I0(n2789), .I1(n2819), .CO(n28415));
    SB_CARRY mod_5_add_1004_10 (.CI(n28006), .I0(n1402), .I1(n1433), .CO(n28007));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n28413), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n28005), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n28413), .I0(n2790), .I1(n2819), .CO(n28414));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n28412), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n28412), .I0(n2791), .I1(n2819), .CO(n28413));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n28411), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n28411), .I0(n2792), .I1(n2819), .CO(n28412));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n28410), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n28410), .I0(n2793), .I1(n2819), .CO(n28411));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n28409), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n28409), .I0(n2794), .I1(n2819), .CO(n28410));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n28408), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_17 (.CI(n28408), .I0(n2795), .I1(n2819), .CO(n28409));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n28407), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n28407), .I0(n2796), .I1(n2819), .CO(n28408));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n28406), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n28406), .I0(n2797), .I1(n2819), .CO(n28407));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n28405), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n28405), .I0(n2798), .I1(n2819), .CO(n28406));
    SB_CARRY mod_5_add_1004_9 (.CI(n28005), .I0(n1403), .I1(n1433), .CO(n28006));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n28404), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n28404), .I0(n2799), .I1(n2819), .CO(n28405));
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n28004), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n28701), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n28403), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_12 (.CI(n28403), .I0(n2800), .I1(n2819), .CO(n28404));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n28402), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_11 (.CI(n28402), .I0(n2801), .I1(n2819), .CO(n28403));
    SB_CARRY mod_5_add_1004_8 (.CI(n28004), .I0(n1404), .I1(n1433), .CO(n28005));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n28003), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n28003), .I0(n1405), .I1(n1433), .CO(n28004));
    SB_CARRY mod_5_add_1339_12 (.CI(n28701), .I0(n1900), .I1(n1928), .CO(n28702));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n28002), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n28002), .I0(n1406), .I1(n1433), .CO(n28003));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n28001), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n28401), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n27783), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_10 (.CI(n28401), .I0(n2802), .I1(n2819), .CO(n28402));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n28700), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n28400), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_9 (.CI(n28400), .I0(n2803), .I1(n2819), .CO(n28401));
    SB_CARRY mod_5_add_1339_11 (.CI(n28700), .I0(n1901), .I1(n1928), .CO(n28701));
    SB_CARRY mod_5_add_1004_5 (.CI(n28001), .I0(n1407), .I1(n1433), .CO(n28002));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n28699), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n28699), .I0(n1902), .I1(n1928), .CO(n28700));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n28399), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n28698), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n28698), .I0(n1903), .I1(n1928), .CO(n28699));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n28000), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n28000), .I0(n1408), .I1(n1433), .CO(n28001));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n37312), 
            .I3(n27999), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_8 (.CI(n28399), .I0(n2804), .I1(n2819), .CO(n28400));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n28398), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n28697), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_7 (.CI(n28398), .I0(n2805), .I1(n2819), .CO(n28399));
    SB_CARRY mod_5_add_1339_8 (.CI(n28697), .I0(n1904), .I1(n1928), .CO(n28698));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n28397), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n28397), .I0(n2806), .I1(n2819), .CO(n28398));
    SB_LUT4 i28616_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n35012));
    defparam i28616_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1579 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_4797));
    defparam i2_3_lut_adj_1579.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut (.I0(n2), .I1(n6_adj_4797), .I2(n1005), .I3(n35012), 
            .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i30581_2_lut (.I0(n2), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4730));   // verilog/neopixel.v(22[26:36])
    defparam i30581_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n28696), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n28396), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n28396), .I0(n2807), .I1(n2819), .CO(n28397));
    SB_CARRY mod_5_add_1339_7 (.CI(n28696), .I0(n1905), .I1(n1928), .CO(n28697));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n28395), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_6 (.CI(n27783), .I0(n906), .I1(VCC_net), .CO(n27784));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n28695), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n28395), .I0(n2808), .I1(n2819), .CO(n28396));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n37314), 
            .I3(n28394), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n28394), .I0(n2809), .I1(n37314), .CO(n28395));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n37314), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n37314), 
            .CO(n28394));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n28393), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n28695), .I0(n1906), .I1(n1928), .CO(n28696));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n28694), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n28392), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n28392), .I0(n2886), .I1(n2918), .CO(n28393));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n28391), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n28391), .I0(n2887), .I1(n2918), .CO(n28392));
    SB_LUT4 i4816_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n33158), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i4816_2_lut_3_lut_4_lut.LUT_INIT = 16'hff90;
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n28390), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n28390), .I0(n2888), .I1(n2918), .CO(n28391));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n28389), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n28389), .I0(n2889), .I1(n2918), .CO(n28390));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n33247), .I2(VCC_net), 
            .I3(n27782), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n28388), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n28694), .I0(n1907), .I1(n1928), .CO(n28695));
    SB_CARRY mod_5_add_2009_22 (.CI(n28388), .I0(n2890), .I1(n2918), .CO(n28389));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n28387), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_21 (.CI(n28387), .I0(n2891), .I1(n2918), .CO(n28388));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n28386), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n28386), .I0(n2892), .I1(n2918), .CO(n28387));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n28385), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_19 (.CI(n28385), .I0(n2893), .I1(n2918), .CO(n28386));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n28693), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n28384), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n28693), .I0(n1908), .I1(n1928), .CO(n28694));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n37313), 
            .I3(n28692), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_18 (.CI(n28384), .I0(n2894), .I1(n2918), .CO(n28385));
    SB_CARRY mod_5_add_1339_3 (.CI(n28692), .I0(n1909), .I1(n37313), .CO(n28693));
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n28383), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n28383), .I0(n2895), .I1(n2918), .CO(n28384));
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n28382), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_16 (.CI(n28382), .I0(n2896), .I1(n2918), .CO(n28383));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n28381), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n28381), .I0(n2897), .I1(n2918), .CO(n28382));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n27675), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n28380), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30925_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37320));
    defparam i30925_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_14 (.CI(n28380), .I0(n2898), .I1(n2918), .CO(n28381));
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n7966), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[29]), .O(n29899));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h45ba;
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n37313), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n28379), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(n7966), .I1(bit_ctr[30]), 
            .I2(bit_ctr[31]), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hb60c;
    SB_CARRY mod_5_add_2009_13 (.CI(n28379), .I0(n2899), .I1(n2918), .CO(n28380));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n28378), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_5 (.CI(n27782), .I0(n33247), .I1(VCC_net), 
            .CO(n27783));
    SB_CARRY mod_5_add_1004_3 (.CI(n27999), .I0(n1409), .I1(n37312), .CO(n28000));
    SB_CARRY mod_5_add_2009_12 (.CI(n28378), .I0(n2900), .I1(n2918), .CO(n28379));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n28377), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n28377), .I0(n2901), .I1(n2918), .CO(n28378));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n28376), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n37312), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_10 (.CI(n28376), .I0(n2902), .I1(n2918), .CO(n28377));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n28375), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_9 (.CI(n28375), .I0(n2903), .I1(n2918), .CO(n28376));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n28374), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n18398), .I2(VCC_net), 
            .I3(n27781), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n37313), 
            .CO(n28692));
    SB_DFF timer_1544__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n28691), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n28690), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n28690), .I0(n1995), .I1(n2027), .CO(n28691));
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n37312), 
            .CO(n27999));
    SB_CARRY mod_5_add_2009_8 (.CI(n28374), .I0(n2904), .I1(n2918), .CO(n28375));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n28373), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n28373), .I0(n2905), .I1(n2918), .CO(n28374));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n28689), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n28689), .I0(n1996), .I1(n2027), .CO(n28690));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n28372), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n28372), .I0(n2906), .I1(n2918), .CO(n28373));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n28371), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n28371), .I0(n2907), .I1(n2918), .CO(n28372));
    SB_CARRY mod_5_add_669_4 (.CI(n27781), .I0(n18398), .I1(VCC_net), 
            .CO(n27782));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n28370), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n28688), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_4 (.CI(n28370), .I0(n2908), .I1(n2918), .CO(n28371));
    SB_CARRY mod_5_add_1406_15 (.CI(n28688), .I0(n1997), .I1(n2027), .CO(n28689));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n28687), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n28687), .I0(n1998), .I1(n2027), .CO(n28688));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n28686), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n28686), .I0(n1999), .I1(n2027), .CO(n28687));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n37315), 
            .I3(n28369), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n28369), .I0(n2909), .I1(n37315), .CO(n28370));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n37315), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n37315), 
            .CO(n28369));
    SB_CARRY add_21_12 (.CI(n27675), .I0(bit_ctr[10]), .I1(GND_net), .CO(n27676));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n28685), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n28685), .I0(n2000), .I1(n2027), .CO(n28686));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n28684), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n28684), .I0(n2001), .I1(n2027), .CO(n28685));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n28368), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n28367), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n28367), .I0(n2985), .I1(n3017), .CO(n28368));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n15590), .I2(GND_net), 
            .I3(n27780), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n28366), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n28366), .I0(n2986), .I1(n3017), .CO(n28367));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n28365), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n28683), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n28365), .I0(n2987), .I1(n3017), .CO(n28366));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n28364), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n28683), .I0(n2002), .I1(n2027), .CO(n28684));
    SB_CARRY mod_5_add_2076_24 (.CI(n28364), .I0(n2988), .I1(n3017), .CO(n28365));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n28363), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n28363), .I0(n2989), .I1(n3017), .CO(n28364));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n28362), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n28362), .I0(n2990), .I1(n3017), .CO(n28363));
    SB_CARRY mod_5_add_669_3 (.CI(n27780), .I0(n15590), .I1(GND_net), 
            .CO(n27781));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n28361), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n28361), .I0(n2991), .I1(n3017), .CO(n28362));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n28360), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n28360), .I0(n2992), .I1(n3017), .CO(n28361));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n28682), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_9 (.CI(n28682), .I0(n2003), .I1(n2027), .CO(n28683));
    SB_LUT4 i3_2_lut_adj_1580 (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4799));
    defparam i3_2_lut_adj_1580.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut_adj_1581 (.I0(bit_ctr[12]), .I1(n22_adj_4799), .I2(n2299), 
            .I3(n2309), .O(n30_adj_4800));
    defparam i11_4_lut_adj_1581.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut_adj_1582 (.I0(n2294), .I1(n30_adj_4800), .I2(n2306), 
            .I3(n2297), .O(n34_adj_4801));
    defparam i15_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1583 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4802));
    defparam i13_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1584 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4803));
    defparam i14_4_lut_adj_1584.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1585 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4804));
    defparam i12_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1586 (.I0(n31_adj_4804), .I1(n33_adj_4803), .I2(n32_adj_4802), 
            .I3(n34_adj_4801), .O(n2324));
    defparam i18_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n28359), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_19 (.CI(n28359), .I0(n2993), .I1(n3017), .CO(n28360));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n28681), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n27674), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n28358), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n27667), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_18 (.CI(n28358), .I0(n2994), .I1(n3017), .CO(n28359));
    SB_CARRY mod_5_add_1406_8 (.CI(n28681), .I0(n2004), .I1(n2027), .CO(n28682));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n28680), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n28680), .I0(n2005), .I1(n2027), .CO(n28681));
    SB_CARRY add_21_9 (.CI(n27672), .I0(bit_ctr[7]), .I1(GND_net), .CO(n27673));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n28679), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n28357), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n28679), .I0(n2006), .I1(n2027), .CO(n28680));
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1587 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4805));
    defparam i14_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1588 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4806));
    defparam i3_3_lut_adj_1588.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1589 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4807));
    defparam i12_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1590 (.I0(n25_adj_4806), .I1(n36_adj_4805), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4808));
    defparam i18_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1591 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4809));
    defparam i16_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4807), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4810));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1592 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4811));
    defparam i15_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1593 (.I0(n37_adj_4811), .I1(n39_adj_4810), .I2(n38_adj_4809), 
            .I3(n40_adj_4808), .O(n2621));
    defparam i21_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i30904_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37299));
    defparam i30904_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_17 (.CI(n28357), .I0(n2995), .I1(n3017), .CO(n28358));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n28356), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n28356), .I0(n2996), .I1(n3017), .CO(n28357));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n28355), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n28355), .I0(n2997), .I1(n3017), .CO(n28356));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n28354), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n28678), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n28354), .I0(n2998), .I1(n3017), .CO(n28355));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n28353), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_4 (.CI(n27667), .I0(bit_ctr[2]), .I1(GND_net), .CO(n27668));
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n27780));
    SB_CARRY mod_5_add_2076_13 (.CI(n28353), .I0(n2999), .I1(n3017), .CO(n28354));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n28352), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n28352), .I0(n3000), .I1(n3017), .CO(n28353));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n28351), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n28351), .I0(n3001), .I1(n3017), .CO(n28352));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n28350), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n28350), .I0(n3002), .I1(n3017), .CO(n28351));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n28349), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n28349), .I0(n3003), .I1(n3017), .CO(n28350));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n28348), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30905_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37300));
    defparam i30905_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1594 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4812));
    defparam i10_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1595 (.I0(n2203), .I1(n28_adj_4812), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4813));
    defparam i14_4_lut_adj_1595.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1596 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4814));
    defparam i12_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2076_8 (.CI(n28348), .I0(n3004), .I1(n3017), .CO(n28349));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n28347), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_7 (.CI(n28347), .I0(n3005), .I1(n3017), .CO(n28348));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n28346), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n28346), .I0(n3006), .I1(n3017), .CO(n28347));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n28345), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n28345), .I0(n3007), .I1(n3017), .CO(n28346));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n28344), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n28344), .I0(n3008), .I1(n3017), .CO(n28345));
    SB_CARRY mod_5_add_1406_5 (.CI(n28678), .I0(n2007), .I1(n2027), .CO(n28679));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n37317), 
            .I3(n28343), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n28343), .I0(n3009), .I1(n37317), .CO(n28344));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n37317), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n28677), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n28677), .I0(n2008), .I1(n2027), .CO(n28678));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n37317), 
            .CO(n28343));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n37316), 
            .I3(n28676), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n28342), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n27673), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n28341), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n28341), .I0(n3084), .I1(n3116), .CO(n28342));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n28340), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n28340), .I0(n3085), .I1(n3116), .CO(n28341));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n28339), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut_adj_1597 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4815));
    defparam i13_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1598 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4816));
    defparam i11_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1599 (.I0(n29_adj_4816), .I1(n31_adj_4815), .I2(n30_adj_4814), 
            .I3(n32_adj_4813), .O(n2225));
    defparam i17_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_26 (.CI(n28339), .I0(n3086), .I1(n3116), .CO(n28340));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n28338), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n28338), .I0(n3087), .I1(n3116), .CO(n28339));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n28337), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n28337), .I0(n3088), .I1(n3116), .CO(n28338));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n28336), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n28336), .I0(n3089), .I1(n3116), .CO(n28337));
    SB_CARRY add_21_10 (.CI(n27673), .I0(bit_ctr[8]), .I1(GND_net), .CO(n27674));
    SB_CARRY mod_5_add_1406_3 (.CI(n28676), .I0(n2009), .I1(n37316), .CO(n28677));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n28335), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n28335), .I0(n3090), .I1(n3116), .CO(n28336));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n37316), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n28334), .O(n47_adj_4755)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n28334), .I0(n3091), .I1(n3116), .CO(n28335));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n28333), .O(n45_adj_4761)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n28333), .I0(n3092), .I1(n3116), .CO(n28334));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n28332), .O(n43_adj_4751)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n28332), .I0(n3093), .I1(n3116), .CO(n28333));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n28331), .O(n41_adj_4759)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n28331), .I0(n3094), .I1(n3116), .CO(n28332));
    SB_LUT4 i3_2_lut_adj_1600 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4817));
    defparam i3_2_lut_adj_1600.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1601 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4818));
    defparam i13_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1602 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4819));
    defparam i1_3_lut_adj_1602.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1603 (.I0(n2490), .I1(n34_adj_4818), .I2(n24_adj_4817), 
            .I3(n2494), .O(n38_adj_4820));
    defparam i17_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1604 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4821));
    defparam i15_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1605 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4819), 
            .O(n37_adj_4822));
    defparam i16_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n28330), .O(n39_adj_4748)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n37316), 
            .CO(n28676));
    SB_CARRY mod_5_add_2143_17 (.CI(n28330), .I0(n3095), .I1(n3116), .CO(n28331));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n28329), .O(n37_adj_4746)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n28329), .I0(n3096), .I1(n3116), .CO(n28330));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n28328), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n28328), .I0(n3097), .I1(n3116), .CO(n28329));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n28327), .O(n33_adj_4754)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n27666), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_14 (.CI(n28327), .I0(n3098), .I1(n3116), .CO(n28328));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n28675), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n28326), .O(n31_adj_4758)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n28326), .I0(n3099), .I1(n3116), .CO(n28327));
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n28325), .O(n29_adj_4745)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1606 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4823));
    defparam i14_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2143_12 (.CI(n28325), .I0(n3100), .I1(n3116), .CO(n28326));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n28324), .O(n27_adj_4750)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n28324), .I0(n3101), .I1(n3116), .CO(n28325));
    SB_CARRY add_21_3 (.CI(n27666), .I0(bit_ctr[1]), .I1(GND_net), .CO(n27667));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n28323), .O(n25_adj_4753)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n28323), .I0(n3102), .I1(n3116), .CO(n28324));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n27672), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n28322), .O(n23_adj_4747)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n28322), .I0(n3103), .I1(n3116), .CO(n28323));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n28321), .O(n21_adj_4764)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n28321), .I0(n3104), .I1(n3116), .CO(n28322));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n28320), .O(n19_adj_4763)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_7 (.CI(n28320), .I0(n3105), .I1(n3116), .CO(n28321));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n28319), .O(n17_adj_4756)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n28319), .I0(n3106), .I1(n3116), .CO(n28320));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n28318), .O(n15_adj_4757)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n28318), .I0(n3107), .I1(n3116), .CO(n28319));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n28317), .O(n13_adj_4762)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n28317), .I0(n3108), .I1(n3116), .CO(n28318));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n37318), 
            .I3(n28316), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_3 (.CI(n28316), .I0(n3109), .I1(n37318), .CO(n28317));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n37318), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n37318), 
            .CO(n28316));
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n28674), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29818_2_lut_4_lut (.I0(LED_c), .I1(bit_ctr[3]), .I2(bit_ctr[4]), 
            .I3(n14682), .O(n35911));   // verilog/neopixel.v(16[20:25])
    defparam i29818_2_lut_4_lut.LUT_INIT = 16'haa80;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n37538));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37538_bdd_4_lut (.I0(n37538), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n37541));
    defparam n37538_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i26804_2_lut_4_lut (.I0(bit_ctr[28]), .I1(n7966), .I2(n608), 
            .I3(bit_ctr[29]), .O(n33188));
    defparam i26804_2_lut_4_lut.LUT_INIT = 16'h02a8;
    SB_LUT4 i3896_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n7966));   // verilog/neopixel.v(22[26:36])
    defparam i3896_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i30903_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37298));
    defparam i30903_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1607 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4824));
    defparam i6_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1608 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4825));
    defparam i1_3_lut_adj_1608.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1609 (.I0(n9_adj_4825), .I1(n14_adj_4824), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i29748_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n739), .I2(bit_ctr[27]), 
            .I3(n838), .O(n18398));
    defparam i29748_3_lut_4_lut.LUT_INIT = 16'h9969;
    SB_LUT4 bit_ctr_0__bdd_4_lut_31104 (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n37478));
    defparam bit_ctr_0__bdd_4_lut_31104.LUT_INIT = 16'he4aa;
    SB_LUT4 n37478_bdd_4_lut (.I0(n37478), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n35154));
    defparam n37478_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_31054 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n37472));
    defparam bit_ctr_0__bdd_4_lut_31054.LUT_INIT = 16'he4aa;
    SB_LUT4 n37472_bdd_4_lut (.I0(n37472), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n35157));
    defparam n37472_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(n26386), 
            .I3(\neo_pixel_transmitter.done ), .O(n34915));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 bit_ctr_0__bdd_4_lut_31049 (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n37460));
    defparam bit_ctr_0__bdd_4_lut_31049.LUT_INIT = 16'he4aa;
    SB_LUT4 n37460_bdd_4_lut (.I0(n37460), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n35163));
    defparam n37460_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n27666));
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n27696), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n27695), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_32 (.CI(n27695), .I0(bit_ctr[30]), .I1(GND_net), .CO(n27696));
    SB_LUT4 bit_ctr_0__bdd_4_lut_31039 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n37424));
    defparam bit_ctr_0__bdd_4_lut_31039.LUT_INIT = 16'he4aa;
    SB_LUT4 n37424_bdd_4_lut (.I0(n37424), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n37427));
    defparam n37424_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n27694), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_18 (.CI(n28674), .I0(n2094), .I1(n2126), .CO(n28675));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n28673), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_31 (.CI(n27694), .I0(bit_ctr[29]), .I1(GND_net), .CO(n27695));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n27693), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n27693), .I0(bit_ctr[28]), .I1(GND_net), .CO(n27694));
    SB_CARRY mod_5_add_1473_17 (.CI(n28673), .I0(n2095), .I1(n2126), .CO(n28674));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n27692), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n27692), .I0(bit_ctr[27]), .I1(GND_net), .CO(n27693));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n28672), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n28672), .I0(n2096), .I1(n2126), .CO(n28673));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n28671), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n28671), .I0(n2097), .I1(n2126), .CO(n28672));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n28670), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n27691), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_28 (.CI(n27691), .I0(bit_ctr[26]), .I1(GND_net), .CO(n27692));
    SB_CARRY mod_5_add_1473_14 (.CI(n28670), .I0(n2098), .I1(n2126), .CO(n28671));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n27671), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n28669), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n28669), .I0(n2099), .I1(n2126), .CO(n28670));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n27690), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_27 (.CI(n27690), .I0(bit_ctr[25]), .I1(GND_net), .CO(n27691));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n27689), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n28668), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_26 (.CI(n27689), .I0(bit_ctr[24]), .I1(GND_net), .CO(n27690));
    SB_CARRY mod_5_add_1473_12 (.CI(n28668), .I0(n2100), .I1(n2126), .CO(n28669));
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n27688), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n28667), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_25 (.CI(n27688), .I0(bit_ctr[23]), .I1(GND_net), .CO(n27689));
    SB_CARRY mod_5_add_1473_11 (.CI(n28667), .I0(n2101), .I1(n2126), .CO(n28668));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n28666), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n27687), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_10 (.CI(n28666), .I0(n2102), .I1(n2126), .CO(n28667));
    SB_CARRY add_21_24 (.CI(n27687), .I0(bit_ctr[22]), .I1(GND_net), .CO(n27688));
    SB_CARRY add_21_11 (.CI(n27674), .I0(bit_ctr[9]), .I1(GND_net), .CO(n27675));
    SB_LUT4 i7_3_lut_adj_1610 (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), 
            .I3(GND_net), .O(n27_adj_4826));
    defparam i7_3_lut_adj_1610.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1611 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4827));
    defparam i13_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n28665), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n7_adj_4770), 
            .D(state_3__N_365[0]), .S(n26337));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1473_9 (.CI(n28665), .I0(n2103), .I1(n2126), .CO(n28666));
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n27686), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n27686), .I0(bit_ctr[21]), .I1(GND_net), .CO(n27687));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n28664), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n28664), .I0(n2104), .I1(n2126), .CO(n28665));
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n27685), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n28663), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_22 (.CI(n27685), .I0(bit_ctr[20]), .I1(GND_net), .CO(n27686));
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n27684), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_7 (.CI(n28663), .I0(n2105), .I1(n2126), .CO(n28664));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n28662), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n28662), .I0(n2106), .I1(n2126), .CO(n28663));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n28661), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n18162), 
            .D(n255[0]), .R(n18520));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE start_103 (.Q(start), .C(clk32MHz), .E(VCC_net), .D(n31374));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n19149));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n19148));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n19147));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n19146));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n19145));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n19144));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n19143));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n19142));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n19141));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n19140));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n19139));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n19138));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n19137));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n19136));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n19135));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n19134));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n19133));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n19132));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n19131));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n19130));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n19129));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n19128));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n19127));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n19126));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n19125));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n19124));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n19123));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n19122));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n19121));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n19120));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n19119));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1473_5 (.CI(n28661), .I0(n2107), .I1(n2126), .CO(n28662));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n28660), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n28660), .I0(n2108), .I1(n2126), .CO(n28661));
    SB_LUT4 i12_4_lut_adj_1612 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4830));
    defparam i12_4_lut_adj_1612.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1613 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4831));
    defparam i11_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1614 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4832));
    defparam i15_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1615 (.I0(n33_adj_4827), .I1(n27_adj_4826), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4833));
    defparam i17_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1616 (.I0(n37_adj_4833), .I1(n35_adj_4832), .I2(n31_adj_4831), 
            .I3(n32_adj_4830), .O(n2423));
    defparam i19_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n37319), 
            .I3(n28659), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_516[25]), .I1(timer[31]), 
            .I2(n56[31]), .I3(n27877), .O(n22_adj_4733)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1473_3 (.CI(n28659), .I0(n2109), .I1(n37319), .CO(n28660));
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_516[24]), .I1(timer[30]), 
            .I2(n56[30]), .I3(n27876), .O(n23_adj_4732)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n37319), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_32 (.CI(n27876), .I0(timer[30]), .I1(n56[30]), 
            .CO(n27877));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_516[19]), .I1(timer[29]), 
            .I2(n56[29]), .I3(n27875), .O(n28_adj_4736)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n27875), .I0(timer[29]), .I1(n56[29]), 
            .CO(n27876));
    SB_CARRY add_21_21 (.CI(n27684), .I0(bit_ctr[19]), .I1(GND_net), .CO(n27685));
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n37319), 
            .CO(n28659));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_516[26]), .I1(timer[28]), 
            .I2(n56[28]), .I3(n27874), .O(n26_adj_4735)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n27683), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n28658), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n28657), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_30 (.CI(n27874), .I0(timer[28]), .I1(n56[28]), 
            .CO(n27875));
    SB_CARRY mod_5_add_1540_19 (.CI(n28657), .I0(n2193), .I1(n2225), .CO(n28658));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_516[18]), .I1(timer[27]), 
            .I2(n56[27]), .I3(n27873), .O(n21_adj_4731)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_20 (.CI(n27683), .I0(bit_ctr[18]), .I1(GND_net), .CO(n27684));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n27682), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n28656), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n28656), .I0(n2194), .I1(n2225), .CO(n28657));
    SB_CARRY sub_14_add_2_29 (.CI(n27873), .I0(timer[27]), .I1(n56[27]), 
            .CO(n27874));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n56[26]), 
            .I3(n27872), .O(one_wire_N_516[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_28 (.CI(n27872), .I0(timer[26]), .I1(n56[26]), 
            .CO(n27873));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n28655), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n33275), .D(\neo_pixel_transmitter.done_N_579 ), 
            .R(n34915));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_19 (.CI(n27682), .I0(bit_ctr[17]), .I1(GND_net), .CO(n27683));
    SB_CARRY mod_5_add_1540_17 (.CI(n28655), .I0(n2195), .I1(n2225), .CO(n28656));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n56[25]), 
            .I3(n27871), .O(one_wire_N_516[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n27681), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n28654), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_18 (.CI(n27681), .I0(bit_ctr[16]), .I1(GND_net), .CO(n27682));
    SB_CARRY sub_14_add_2_27 (.CI(n27871), .I0(timer[25]), .I1(n56[25]), 
            .CO(n27872));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n56[24]), 
            .I3(n27870), .O(one_wire_N_516[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_16 (.CI(n28654), .I0(n2196), .I1(n2225), .CO(n28655));
    SB_CARRY sub_14_add_2_26 (.CI(n27870), .I0(timer[24]), .I1(n56[24]), 
            .CO(n27871));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n28653), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_516[16]), .I1(timer[23]), 
            .I2(n56[23]), .I3(n27869), .O(n30_adj_4738)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n27680), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_25 (.CI(n27869), .I0(timer[23]), .I1(n56[23]), 
            .CO(n27870));
    SB_LUT4 i25_4_lut_adj_1617 (.I0(n26348), .I1(n26349), .I2(\state[1] ), 
            .I3(\state[0] ), .O(n11_adj_4842));   // verilog/neopixel.v(16[20:25])
    defparam i25_4_lut_adj_1617.LUT_INIT = 16'hcafa;
    SB_CARRY mod_5_add_1540_15 (.CI(n28653), .I0(n2197), .I1(n2225), .CO(n28654));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n28652), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n28652), .I0(n2198), .I1(n2225), .CO(n28653));
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n11_adj_4842));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1544__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1544__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n56[22]), 
            .I3(n27868), .O(one_wire_N_516[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n28651), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_24 (.CI(n27868), .I0(timer[22]), .I1(n56[22]), 
            .CO(n27869));
    SB_CARRY add_21_17 (.CI(n27680), .I0(bit_ctr[15]), .I1(GND_net), .CO(n27681));
    SB_LUT4 sub_14_add_2_23_lut (.I0(GND_net), .I1(timer[21]), .I2(n56[21]), 
            .I3(n27867), .O(one_wire_N_516[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28083), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28082), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28082), .I0(n1203), .I1(n1235), .CO(n28083));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28081), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n28081), .I0(n1204), .I1(n1235), .CO(n28082));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28080), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n28080), .I0(n1205), .I1(n1235), .CO(n28081));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28079), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n28079), .I0(n1206), .I1(n1235), .CO(n28080));
    SB_CARRY mod_5_add_1540_13 (.CI(n28651), .I0(n2199), .I1(n2225), .CO(n28652));
    SB_LUT4 i20_4_lut_adj_1618 (.I0(n35_adj_4823), .I1(n37_adj_4822), .I2(n36_adj_4821), 
            .I3(n38_adj_4820), .O(n2522));
    defparam i20_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28078), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n27679), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_5 (.CI(n28078), .I0(n1207), .I1(n1235), .CO(n28079));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28077), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n28650), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_23 (.CI(n27867), .I0(timer[21]), .I1(n56[21]), 
            .CO(n27868));
    SB_CARRY mod_5_add_870_4 (.CI(n28077), .I0(n1208), .I1(n1235), .CO(n28078));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n37320), 
            .I3(n28076), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n28076), .I0(n1209), .I1(n37320), .CO(n28077));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_516[15]), .I1(timer[20]), 
            .I2(n56[20]), .I3(n27866), .O(n29_adj_4737)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n37320), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n37320), 
            .CO(n28076));
    SB_CARRY mod_5_add_1540_12 (.CI(n28650), .I0(n2200), .I1(n2225), .CO(n28651));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n28649), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_22 (.CI(n27866), .I0(timer[20]), .I1(n56[20]), 
            .CO(n27867));
    SB_CARRY mod_5_add_1540_11 (.CI(n28649), .I0(n2201), .I1(n2225), .CO(n28650));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n56[19]), 
            .I3(n27865), .O(one_wire_N_516[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_21 (.CI(n27865), .I0(timer[19]), .I1(n56[19]), 
            .CO(n27866));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n28648), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n56[18]), 
            .I3(n27864), .O(one_wire_N_516[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_10 (.CI(n28648), .I0(n2202), .I1(n2225), .CO(n28649));
    SB_CARRY sub_14_add_2_20 (.CI(n27864), .I0(timer[18]), .I1(n56[18]), 
            .CO(n27865));
    SB_LUT4 sub_14_add_2_19_lut (.I0(GND_net), .I1(timer[17]), .I2(n56[17]), 
            .I3(n27863), .O(one_wire_N_516[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n28647), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2_3_lut_4_lut_adj_1619 (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(color_bit), 
            .I3(n14682), .O(state_3__N_365[0]));
    defparam i2_3_lut_4_lut_adj_1619.LUT_INIT = 16'h0070;
    SB_LUT4 i1_2_lut_3_lut_adj_1620 (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(n14682), 
            .I3(GND_net), .O(n26349));
    defparam i1_2_lut_3_lut_adj_1620.LUT_INIT = 16'hf8f8;
    SB_CARRY mod_5_add_1540_9 (.CI(n28647), .I0(n2203), .I1(n2225), .CO(n28648));
    SB_CARRY sub_14_add_2_19 (.CI(n27863), .I0(timer[17]), .I1(n56[17]), 
            .CO(n27864));
    SB_LUT4 i3_4_lut_4_lut (.I0(n33158), .I1(n15594), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n28646), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n18625));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n56[16]), 
            .I3(n27862), .O(one_wire_N_516[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n27862), .I0(timer[16]), .I1(n56[16]), 
            .CO(n27863));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n56[15]), 
            .I3(n27861), .O(one_wire_N_516[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30923_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37318));
    defparam i30923_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30052_4_lut (.I0(n26341), .I1(n33241), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n36260));
    defparam i30052_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i29780_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n36176));
    defparam i29780_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i53_4_lut (.I0(n33241), .I1(n26386), .I2(\state[1] ), .I3(start), 
            .O(n33261));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n33261), .I1(n33146), .I2(n36176), .I3(n36260), 
            .O(n33275));
    defparam i52_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 i108_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_579 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i108_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1621 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4843));
    defparam i1_2_lut_adj_1621.LUT_INIT = 16'heeee;
    SB_LUT4 i19719_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n24500));
    defparam i19719_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1622 (.I0(n2093), .I1(n2108), .I2(n2100), .I3(n18_adj_4843), 
            .O(n30_adj_4844));
    defparam i13_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1623 (.I0(n2098), .I1(n24500), .I2(n2094), .I3(n2099), 
            .O(n28_adj_4845));
    defparam i11_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1624 (.I0(n2105), .I1(n2096), .I2(n2095), .I3(n2102), 
            .O(n29_adj_4846));
    defparam i12_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1625 (.I0(n2101), .I1(n2107), .I2(n2104), .I3(n2106), 
            .O(n27_adj_4847));
    defparam i10_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1626 (.I0(n27_adj_4847), .I1(n29_adj_4846), .I2(n28_adj_4845), 
            .I3(n30_adj_4844), .O(n2126));
    defparam i16_4_lut_adj_1626.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n15594), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n33158), .O(n33247));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n56[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30924_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37319));
    defparam i30924_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_3_lut (.I0(bit_ctr[4]), .I1(n3096), .I2(n3109), .I3(GND_net), 
            .O(n37_adj_4848));
    defparam i10_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i18_4_lut_adj_1627 (.I0(n3088), .I1(n3104), .I2(n3106), .I3(n3108), 
            .O(n45_adj_4849));
    defparam i18_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1628 (.I0(n3083), .I1(n3095), .I2(n3090), .I3(n3107), 
            .O(n42_adj_4850));
    defparam i15_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut_adj_1629 (.I0(n3101), .I1(n3085), .I2(GND_net), .I3(GND_net), 
            .O(n32_adj_4851));
    defparam i5_2_lut_adj_1629.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1630 (.I0(n3093), .I1(n3084), .I2(n3100), .I3(n3103), 
            .O(n44_adj_4852));
    defparam i17_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1631 (.I0(n45_adj_4849), .I1(n37_adj_4848), .I2(n3097), 
            .I3(n3091), .O(n50));
    defparam i23_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1632 (.I0(n3089), .I1(n42_adj_4850), .I2(n3092), 
            .I3(n3099), .O(n48_adj_4853));
    defparam i21_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1633 (.I0(n3086), .I1(n44_adj_4852), .I2(n32_adj_4851), 
            .I3(n3094), .O(n49_adj_4854));
    defparam i22_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1634 (.I0(n3102), .I1(n3098), .I2(n3087), .I3(n3105), 
            .O(n47_adj_4855));
    defparam i20_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1635 (.I0(n47_adj_4855), .I1(n49_adj_4854), .I2(n48_adj_4853), 
            .I3(n50), .O(n3116));
    defparam i26_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i30921_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37316));
    defparam i30921_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30922_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37317));
    defparam i30922_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 bit_ctr_0__bdd_4_lut_31009 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n37340));
    defparam bit_ctr_0__bdd_4_lut_31009.LUT_INIT = 16'he4aa;
    SB_LUT4 n37340_bdd_4_lut (.I0(n37340), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n36546));
    defparam n37340_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n35154), .I2(n35157), 
            .I3(n38250), .O(n37334));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37334_bdd_4_lut (.I0(n37334), .I1(n36546), .I2(n35163), .I3(n38250), 
            .O(n37337));
    defparam n37334_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14_4_lut_adj_1636 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4856));
    defparam i14_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1637 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4857));
    defparam i18_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1638 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_4858));
    defparam i16_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1639 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4859));
    defparam i17_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1640 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4860));
    defparam i15_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_4861));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4856), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4862));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut_adj_1641 (.I0(n41_adj_4860), .I1(n43_adj_4859), .I2(n42_adj_4858), 
            .I3(n44_adj_4857), .O(n50_adj_4863));
    defparam i24_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4864));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut_adj_1642 (.I0(n37_adj_4864), .I1(n50_adj_4863), .I2(n46_adj_4862), 
            .I3(n38_adj_4861), .O(n3017));
    defparam i25_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i30920_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37315));
    defparam i30920_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, clk32MHz, data_o, 
            GND_net, n34883, reg_B, ENCODER1_A_c_1, VCC_net, ENCODER1_B_c_0, 
            n18645, n19185) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder1_position;
    input clk32MHz;
    output [1:0]data_o;
    input GND_net;
    output n34883;
    output [1:0]reg_B;
    input ENCODER1_A_c_1;
    input VCC_net;
    input ENCODER1_B_c_0;
    input n18645;
    input n19185;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n3074;
    
    wire count_enable, B_delayed, A_delayed, count_direction, n3063, 
        n27975, n27974, n27973, n27972, n27971, n27970, n27969, 
        n27968, n27967, n27966, n27965, n27964, n27963, n27962, 
        n27961, n27960, n27959, n27958, n27957, n27956, n27955, 
        n27954, n27953, n27952;
    
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n3074[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1170_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n3063));   // quad.v(37[5] 40[8])
    defparam i1170_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_703_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n3063), 
            .I3(n27975), .O(n3074[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_703_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n3063), 
            .I3(n27974), .O(n3074[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_24 (.CI(n27974), .I0(encoder1_position[22]), .I1(n3063), 
            .CO(n27975));
    SB_LUT4 add_703_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n3063), 
            .I3(n27973), .O(n3074[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_23 (.CI(n27973), .I0(encoder1_position[21]), .I1(n3063), 
            .CO(n27974));
    SB_LUT4 add_703_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n3063), 
            .I3(n27972), .O(n3074[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_22 (.CI(n27972), .I0(encoder1_position[20]), .I1(n3063), 
            .CO(n27973));
    SB_LUT4 add_703_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n3063), 
            .I3(n27971), .O(n3074[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_21 (.CI(n27971), .I0(encoder1_position[19]), .I1(n3063), 
            .CO(n27972));
    SB_LUT4 add_703_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n3063), 
            .I3(n27970), .O(n3074[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_20 (.CI(n27970), .I0(encoder1_position[18]), .I1(n3063), 
            .CO(n27971));
    SB_LUT4 add_703_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n3063), 
            .I3(n27969), .O(n3074[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_19 (.CI(n27969), .I0(encoder1_position[17]), .I1(n3063), 
            .CO(n27970));
    SB_LUT4 add_703_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n3063), 
            .I3(n27968), .O(n3074[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_18 (.CI(n27968), .I0(encoder1_position[16]), .I1(n3063), 
            .CO(n27969));
    SB_LUT4 add_703_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n3063), 
            .I3(n27967), .O(n3074[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_17 (.CI(n27967), .I0(encoder1_position[15]), .I1(n3063), 
            .CO(n27968));
    SB_LUT4 add_703_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n3063), 
            .I3(n27966), .O(n3074[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_16 (.CI(n27966), .I0(encoder1_position[14]), .I1(n3063), 
            .CO(n27967));
    SB_LUT4 add_703_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n3063), 
            .I3(n27965), .O(n3074[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_15 (.CI(n27965), .I0(encoder1_position[13]), .I1(n3063), 
            .CO(n27966));
    SB_LUT4 add_703_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n3063), 
            .I3(n27964), .O(n3074[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_14 (.CI(n27964), .I0(encoder1_position[12]), .I1(n3063), 
            .CO(n27965));
    SB_LUT4 add_703_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n3063), 
            .I3(n27963), .O(n3074[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_13 (.CI(n27963), .I0(encoder1_position[11]), .I1(n3063), 
            .CO(n27964));
    SB_LUT4 add_703_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n3063), 
            .I3(n27962), .O(n3074[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_12 (.CI(n27962), .I0(encoder1_position[10]), .I1(n3063), 
            .CO(n27963));
    SB_LUT4 add_703_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n3063), 
            .I3(n27961), .O(n3074[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_11 (.CI(n27961), .I0(encoder1_position[9]), .I1(n3063), 
            .CO(n27962));
    SB_LUT4 add_703_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n3063), 
            .I3(n27960), .O(n3074[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_10 (.CI(n27960), .I0(encoder1_position[8]), .I1(n3063), 
            .CO(n27961));
    SB_LUT4 add_703_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n3063), 
            .I3(n27959), .O(n3074[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_9 (.CI(n27959), .I0(encoder1_position[7]), .I1(n3063), 
            .CO(n27960));
    SB_LUT4 add_703_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n3063), 
            .I3(n27958), .O(n3074[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_8 (.CI(n27958), .I0(encoder1_position[6]), .I1(n3063), 
            .CO(n27959));
    SB_LUT4 add_703_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n3063), 
            .I3(n27957), .O(n3074[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_7 (.CI(n27957), .I0(encoder1_position[5]), .I1(n3063), 
            .CO(n27958));
    SB_LUT4 add_703_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n3063), 
            .I3(n27956), .O(n3074[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_6 (.CI(n27956), .I0(encoder1_position[4]), .I1(n3063), 
            .CO(n27957));
    SB_LUT4 add_703_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n3063), 
            .I3(n27955), .O(n3074[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_5 (.CI(n27955), .I0(encoder1_position[3]), .I1(n3063), 
            .CO(n27956));
    SB_LUT4 add_703_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n3063), 
            .I3(n27954), .O(n3074[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_4 (.CI(n27954), .I0(encoder1_position[2]), .I1(n3063), 
            .CO(n27955));
    SB_LUT4 add_703_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n3063), 
            .I3(n27953), .O(n3074[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_3 (.CI(n27953), .I0(encoder1_position[1]), .I1(n3063), 
            .CO(n27954));
    SB_LUT4 add_703_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n27952), .O(n3074[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_703_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_703_2 (.CI(n27952), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n27953));
    SB_CARRY add_703_1 (.CI(GND_net), .I0(n3063), .I1(n3063), .CO(n27952));
    \grp_debouncer(2,100)  debounce (.n34883(n34883), .reg_B({reg_B}), .GND_net(GND_net), 
            .ENCODER1_A_c_1(ENCODER1_A_c_1), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .ENCODER1_B_c_0(ENCODER1_B_c_0), .n18645(n18645), .data_o({data_o}), 
            .n19185(n19185));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (n34883, reg_B, GND_net, ENCODER1_A_c_1, 
            clk32MHz, VCC_net, ENCODER1_B_c_0, n18645, data_o, n19185);
    output n34883;
    output [1:0]reg_B;
    input GND_net;
    input ENCODER1_A_c_1;
    input clk32MHz;
    input VCC_net;
    input ENCODER1_B_c_0;
    input n18645;
    output [1:0]data_o;
    input n19185;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3693;
    wire [6:0]n33;
    
    wire n28428, n28427, n28426, n28425, n28424, n28423;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n34883));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n34883), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 cnt_reg_1551_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n28428), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1551_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1551_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n28427), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1551_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1551_add_4_7 (.CI(n28427), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n28428));
    SB_LUT4 cnt_reg_1551_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n28426), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1551_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1551_add_4_6 (.CI(n28426), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n28427));
    SB_LUT4 cnt_reg_1551_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n28425), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1551_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1551_add_4_5 (.CI(n28425), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n28426));
    SB_LUT4 cnt_reg_1551_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n28424), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1551_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1551_add_4_4 (.CI(n28424), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n28425));
    SB_LUT4 cnt_reg_1551_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n28423), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1551_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1551_add_4_3 (.CI(n28423), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n28424));
    SB_LUT4 cnt_reg_1551_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1551_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1551_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n28423));
    SB_DFFSR cnt_reg_1551__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n18645));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n19185));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1551__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1551__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1551__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1551__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1551__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1551__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3693));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Ki[8] , GND_net, IntegralLimit, \Ki[9] , \Ki[10] , 
            \Ki[11] , \Ki[12] , PWMLimit, duty, n37310, \Ki[1] , 
            \Ki[0] , \Ki[2] , \Kp[5] , \Kp[6] , \Kp[7] , \Kp[8] , 
            \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , \Kp[13] , \Kp[14] , 
            \Kp[1] , \Kp[0] , \Kp[2] , \Ki[3] , clk32MHz, \Kp[3] , 
            \Kp[4] , \Ki[4] , \Ki[5] , \Ki[6] , \Ki[7] , VCC_net, 
            \Kp[15] , \Ki[13] , \Ki[14] , \Ki[15] , setpoint, motor_state) /* synthesis syn_module_defined=1 */ ;
    input \Ki[8] ;
    input GND_net;
    input [23:0]IntegralLimit;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input [23:0]PWMLimit;
    output [23:0]duty;
    output n37310;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Ki[3] ;
    input clk32MHz;
    input \Kp[3] ;
    input \Kp[4] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input VCC_net;
    input \Kp[15] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input [23:0]setpoint;
    input [23:0]motor_state;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]\PID_CONTROLLER.integral_23__N_3509 ;
    
    wire n618;
    wire [23:0]n1;
    
    wire n691, n764, n27942;
    wire [23:0]n1_adj_4708;
    
    wire n27943, n837, n910;
    wire [23:0]duty_23__N_3609;
    wire [23:0]n257;
    
    wire n256;
    wire [23:0]duty_23__N_3584;
    
    wire duty_23__N_3608;
    wire [23:0]duty_23__N_3485;
    
    wire n110, n41, n183, n28778;
    wire [20:0]n9373;
    
    wire n734, n28779;
    wire [21:0]n9349;
    
    wire n661, n28777, n588, n28776, n515, n28775, n442, n28774, 
        n369, n28773, n27941, n296, n28772;
    wire [23:0]n28;
    
    wire n393, n466, n539, n612, n685, n758, n831, n904, \PID_CONTROLLER.integral_23__N_3557 ;
    wire [23:0]n3223;
    
    wire n977, n1050, n104, n35, n177, n223, n28771, n150, n28770, 
        n8_adj_4290, n77, n4_adj_4291;
    wire [3:0]n9925;
    
    wire n6_adj_4292;
    wire [4:0]n9918;
    
    wire n27505;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n27940, n250, n323, n396, n469, n542, n615, n688, n761, 
        n834, n256_adj_4294, n329, n402, n907, n475, n548, n621, 
        n980, n694, n767, n840, n107, n38, n113, n180, n44, 
        n27939, n186, n259, n253, n332, n405, n478, n326, n551, 
        n399, n624, n472, n545, n618_adj_4296, n691_adj_4297, n697, 
        n770, n116, n47, n189, n764_adj_4298, n837_adj_4299, n910_adj_4300, 
        n27582;
    wire [1:0]n9936;
    
    wire n4_adj_4301, n110_adj_4302, n41_adj_4303, n183_adj_4304, n262, 
        n256_adj_4305;
    wire [2:0]n9931;
    
    wire n329_adj_4306, n402_adj_4307, n475_adj_4308, n62, n131, n204, 
        n335, n4_adj_4309, n27938, n408, n548_adj_4310, n621_adj_4312, 
        n694_adj_4313, n481, n767_adj_4315, n840_adj_4316, n554, n113_adj_4317, 
        n44_adj_4318, n627, n700, n119, n50, n192, n265, n338, 
        n411, n484, n186_adj_4319, n259_adj_4320, n557, n332_adj_4321, 
        n630, n122, n405_adj_4322, n53, n195, n268_adj_4324, n478_adj_4325, 
        n341, n414, n487, n560, n27937, n125, n56, n198, n551_adj_4327, 
        n624_adj_4328, n271_adj_4329, n697_adj_4330, n344, n417, n770_adj_4331, 
        n116_adj_4332, n47_adj_4333, n189_adj_4334, n262_adj_4335, n335_adj_4336, 
        n408_adj_4337, n481_adj_4338, n554_adj_4339, n27936, n490, 
        n12_adj_4340, n8_adj_4341, n11_adj_4342, n6_adj_4343, n27607, 
        n18_adj_4344, n627_adj_4345, n700_adj_4346, n119_adj_4347, n50_adj_4348, 
        n192_adj_4349, n13_adj_4350, n34839, n265_adj_4351, n338_adj_4352, 
        n411_adj_4353, n484_adj_4354, n557_adj_4355, n27935, n27934, 
        n27933, n27932, n27931, n630_adj_4360, n122_adj_4361, n53_adj_4363, 
        n195_adj_4364, n268_adj_4365, n27930, n341_adj_4366, n414_adj_4367, 
        n487_adj_4368, n560_adj_4369, n125_adj_4370, n56_adj_4372, n198_adj_4373, 
        n271_adj_4374, n344_adj_4375, n417_adj_4376, n6_adj_4377;
    wire [3:0]n9628;
    wire [4:0]n9621;
    
    wire n27929;
    wire [1:0]n9639;
    
    wire n4_adj_4380;
    wire [2:0]n9634;
    
    wire n490_adj_4382, n12_adj_4385, n8_adj_4386, n11_adj_4387, n6_adj_4388;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3560 ;
    
    wire n27928, n27475, n18_adj_4389, n13_adj_4390, n4_adj_4391, 
        n34155, n807, n880, n77_adj_4393, n8_adj_4394, n45, n27927, 
        n43, n27926, n953, n1026, n41_adj_4395, n27925, n150_adj_4396, 
        n1099, n223_adj_4397, n296_adj_4398, n369_adj_4399, n442_adj_4401, 
        n39, n27924, n37, n27923, n35_adj_4402, n27922, n515_adj_4403, 
        n588_adj_4404, n661_adj_4405, n734_adj_4406, n807_adj_4407, 
        n880_adj_4408, n953_adj_4409, n1026_adj_4410, n1099_adj_4411, 
        n33, n27921;
    wire [47:0]n155;
    wire [47:0]n106;
    
    wire n74, n5_adj_4413, n31, n27920, n147, n220, n74_adj_4414, 
        n293, n366, n439, n512, n5_adj_4416, n585, n658, n731, 
        n804, n147_adj_4417, n877, n950, n220_adj_4418, n293_adj_4419, 
        n1023, n366_adj_4420, n439_adj_4421, n512_adj_4422, n1096;
    wire [5:0]n9910;
    
    wire n29255, n29254, n29253, n29252, n29251, n29, n27919;
    wire [6:0]n9901;
    
    wire n29250, n29249, n29248, n585_adj_4423, n658_adj_4424, n731_adj_4425, 
        n804_adj_4426, n877_adj_4427, n29247, n950_adj_4428, n29246, 
        n1023_adj_4429, n1096_adj_4430, n80, n11_adj_4433, n153, n226, 
        n299, n29245, n372, n445;
    wire [7:0]n9891;
    
    wire n29244, n518, n591, n29243, n29242, n29241, n664, n29240, 
        n29239, n29238, n737;
    wire [8:0]n9880;
    
    wire n29237, n810, n29236, n29235, n27, n27918, n883, n956, 
        n1029, n17_adj_4434, n1102, n9_adj_4435, n11_adj_4436, n29234, 
        n36171, n36168, n38226, n36534, n36428, n38208, n36426, 
        n83, n36424, n38201, n14_adj_4438, n15_adj_4439, n13_adj_4440, 
        n11_adj_4441, n36117, n21_adj_4442, n19_adj_4443, n17_adj_4444, 
        n9_adj_4445, n36123, n156, n39_adj_4446, n41_adj_4447, n45_adj_4448, 
        n43_adj_4449, n16_adj_4450, n29_adj_4452, n229, n31_adj_4453, 
        n23_adj_4454, n25_adj_4455, n37_adj_4456, n35_adj_4457, n36101, 
        n302, n375, n448, n521, n11_adj_4458, n29233, n13_adj_4459, 
        n29232, n15_adj_4460, n27_adj_4461, n29231, n33_adj_4462, 
        n9_adj_4463, n29230, n17_adj_4464, n19_adj_4465, n21_adj_4466;
    wire [9:0]n9868;
    
    wire n29229, n36088, n29228, n36082, n12_adj_4467, n29227, n10_adj_4468, 
        n29226, n30, n29225, n36099, n36362, n36358, n29224, n36657, 
        n29223, n36496, n36719, n29222, n16_adj_4469, n29221, n6_adj_4470, 
        n36633, n36634, n8_adj_4471;
    wire [10:0]n9855;
    
    wire n29220, n24_adj_4472, n29219, n36067, n36065, n36540, n36591, 
        n4_adj_4473, n29218, n36631, n36632, n36077, n36075, n36729, 
        n36593, n36780, n36781, n36760, n36069, n36691, n8_adj_4474, 
        n40, n36693, n41_adj_4475, n39_adj_4476, n23_adj_4477, n25_adj_4478, 
        n45_adj_4479, n43_adj_4480, n37_adj_4481, n29_adj_4482, n31_adj_4483, 
        n35_adj_4484, n33_adj_4485, n29217, n25_adj_4486, n27917, 
        n594, n29216, n29215, n667, n740, n813, n886, n959, 
        n1032, n11_adj_4487, n13_adj_4488, n15_adj_4489, n27_adj_4490, 
        n9_adj_4491, n17_adj_4492, n19_adj_4493, n21_adj_4494, n36051, 
        n36045, n12_adj_4495, n10_adj_4496, n30_adj_4497, n36063, 
        n36330, n36326, n36649, n36480, n36717, n16_adj_4498, n6_adj_4499, 
        n36627, n36628, n8_adj_4500, n1105, n86, n17_adj_4502, n24_adj_4503, 
        n29214, n29213, n29212, n24_adj_4504, n36029, n36027, n36542, 
        n36597, n4_adj_4505, n36625, n36626, n36041, n36039, n36731, 
        n36599, n36782, n36783, n36758, n36031, n36697, n40_adj_4506, 
        n36699, n159, n29211, n7_adj_4507, n5_adj_4508, n36134, 
        n232;
    wire [11:0]n9841;
    
    wire n29210, n36394, n305, n29209, n29208, n378, n23_adj_4509, 
        n27916, n29207, n451, n524, n29206, n545_adj_4510, n29205, 
        n472_adj_4511, n29204, n399_adj_4512, n29203, n326_adj_4513, 
        n29202, n253_adj_4514, n29201, n180_adj_4515, n29200, n597, 
        n38_adj_4516, n107_adj_4517;
    wire [12:0]n9826;
    
    wire n980_adj_4518, n29199, n907_adj_4519, n29198, n670, n834_adj_4520, 
        n29197, n27915, n36390, n743, n761_adj_4522, n29196, n27914, 
        n688_adj_4524, n29195, n615_adj_4525, n29194, n27913, n542_adj_4527, 
        n29193, n816, n469_adj_4528, n29192, n27912, n396_adj_4530, 
        n29191, n323_adj_4531, n29190, n8_adj_4532, n27911, n889, 
        n250_adj_4534, n29189;
    wire [0:0]n8060;
    wire [0:0]n8064;
    
    wire n27779, n177_adj_4535, n29188, n35_adj_4536, n104_adj_4537;
    wire [13:0]n9810;
    
    wire n1050_adj_4538, n29187, n36665, n977_adj_4539, n29186, n27910, 
        n27909, n27778, n36512, n27908, n904_adj_4543, n29185, n962, 
        n831_adj_4544, n29184, n758_adj_4545, n29183, n685_adj_4546, 
        n29182, n1035, n36721, n612_adj_4547, n29181, n539_adj_4548, 
        n29180, n466_adj_4549, n29179, n393_adj_4550, n29178, n320, 
        n29177, n247, n29176, n27777, n174, n29175, n32, n101;
    wire [14:0]n9793;
    
    wire n1120, n29174, n1047, n29173, n36430, n38195, n974, n29172, 
        n36418, n1108, n901, n29171, n38189, n828, n29170, n755, 
        n29169, n682, n29168, n609, n29167, n536, n29166, n463, 
        n29165, n390, n29164, n12_adj_4551, n36147, n317, n29163, 
        n244, n29162, n171, n29161, n38213, n29_adj_4552, n98, 
        n10_adj_4553;
    wire [15:0]n9775;
    
    wire n29160, n30_adj_4554, n1117, n29159, n1044, n29158, n36576, 
        n971, n29157, n898, n29156, n825, n29155, n752, n29154, 
        n679, n29153, n606, n29152, n27907, n36156, n27776, n533, 
        n29151, n460, n29150, n38193, n36528, n38219, n36671, 
        n387, n29149, n3_adj_4557, n27906, n38184, n89, n314, 
        n29148, n241, n29147, n168, n29146, n20_adj_4560, n36743, 
        n26_adj_4561, n95;
    wire [16:0]n9756;
    
    wire n29145, n29144, n38181, n16_adj_4562, n162, n1114, n29143, 
        n1041, n29142, n36136, n968, n29141, n895, n29140, n822, 
        n29139, n235, n749, n29138, n676, n29137, n24_adj_4563, 
        n603, n29136, n530, n29135, n457, n29134, n6_adj_4564, 
        n384, n29133, n311, n29132, n36675, n238, n29131, n165, 
        n29130, n23_adj_4565, n92;
    wire [17:0]n9736;
    
    wire n29129, n29128, n29127, n1111, n29126, n1038, n29125, 
        n36676, n308, n36138, n38179, n36536, n965, n29124, n892, 
        n29123, n36579, n4_adj_4566, n381, n36643, n454, n36644, 
        n12_adj_4567, n819, n29122, n36111, n527, n746, n29121, 
        n10_adj_4568, n30_adj_4570, n600, n673, n36113, n746_adj_4571, 
        n673_adj_4572, n29120, n819_adj_4573, n600_adj_4574, n29119, 
        n527_adj_4575, n29118, n454_adj_4576, n29117, n892_adj_4577, 
        n381_adj_4578, n29116, n308_adj_4579, n29115, n235_adj_4580, 
        n29114, n162_adj_4581, n29113, n20_adj_4582, n89_adj_4583;
    wire [18:0]n9715;
    
    wire n29112, n29111, n29110, n29109, n1108_adj_4584, n29108, 
        n1035_adj_4585, n29107, n962_adj_4586, n29106, n889_adj_4587, 
        n29105, n816_adj_4588, n29104, n743_adj_4589, n29103, n36727, 
        n670_adj_4590, n29102, n597_adj_4591, n29101, n524_adj_4592, 
        n29100, n36587, n451_adj_4593, n29099, n378_adj_4594, n29098, 
        n305_adj_4595, n29097, n232_adj_4596, n29096, n965_adj_4597, 
        n36778, n36779, n36762, n6_adj_4598, n159_adj_4599, n29095, 
        n1038_adj_4600, n17_adj_4601, n86_adj_4602;
    wire [19:0]n9693;
    
    wire n29094, n29093, n29092, n29091, n29090, n36651, n36652, 
        n36103, n36538, n36585, n1111_adj_4603, n36105, n36685, 
        n1105_adj_4604, n29089, n1032_adj_4605, n29088, n27775, n40_adj_4606, 
        n36687, n959_adj_4607, n29087, n886_adj_4608, n29086, n4_adj_4609, 
        n813_adj_4610, n29085, n36667, n36668, n36149, n36725, n740_adj_4611, 
        n29084, n27774, n36581, n667_adj_4612, n29083, n36776, n36777, 
        n36764, n27773, n594_adj_4614, n29082, n521_adj_4615, n29081, 
        n448_adj_4616, n29080, n375_adj_4617, n29079, n302_adj_4618, 
        n29078, n229_adj_4619, n29077, n156_adj_4620, n29076, n14_adj_4621, 
        n83_adj_4622;
    wire [20:0]n9670;
    
    wire n29075, n29074, n29073, n29072, n29071, n29070, n1102_adj_4623, 
        n29069, n1029_adj_4624, n29068, n956_adj_4625, n29067, n883_adj_4626, 
        n29066, n27900, n810_adj_4627, n29065, n27772, n737_adj_4628, 
        n29064, n27899, n664_adj_4629, n29063, n591_adj_4630, n29062, 
        n518_adj_4631, n29061, n445_adj_4632, n29060, n372_adj_4633, 
        n29059, n299_adj_4634, n29058, n226_adj_4635, n29057, n153_adj_4636, 
        n29056, n11_adj_4637, n80_adj_4638, n27898, n36140;
    wire [21:0]n9646;
    
    wire n29055, n29054, n36679, n29053, n40_adj_4639, \PID_CONTROLLER.integral_23__N_3559 , 
        n29052, n27897, n92_adj_4640, n36681, n29051, n23_adj_4642, 
        n29050, n27771, n27896, n27822, n27821, n27895, n27894, 
        n165_adj_4643, n27770, n27820, n27893, n27892, n29049, n29048, 
        n29047, n29046, n27769, n29045, n29044, n29043, n29042, 
        n29041, n29040, n27891, n27819, n29039, n29038, n27818, 
        n29037, n29036, n29035, n27890, n29034, n27817, n29033, 
        n29032, n29031, n29030, n29029, n29028, n29027, n29026, 
        n29025, n29024, n29023, n29022, n29021, n29020, n29019, 
        n29018, n27889, n29017, n29016, n29015, n29014, n27816, 
        n29013, n27888;
    wire [5:0]n9613;
    
    wire n29012, n29011, n29010, n29009, n29008;
    wire [6:0]n9604;
    
    wire n29007, n29006, n29005, n29004, n29003, n238_adj_4649, 
        n29002, n27815, n27887;
    wire [7:0]n9594;
    
    wire n29001, n29000, n28999, n28998, n28997, n311_adj_4650, 
        n28996, n28995;
    wire [8:0]n9583;
    
    wire n28994, n28993, n28992, n28991, n28990, n28989, n27886, 
        n28988, n28987, n384_adj_4651;
    wire [9:0]n9571;
    
    wire n28986, n28985, n28984, n28983, n28982, n27814, n28981, 
        n28980, n28979, n28978, n27885, n27768;
    wire [10:0]n9558;
    
    wire n28977, n28976, n28975, n28974, n27813, n28973, n457_adj_4653, 
        n27884, n28972, n28971, n28970, n28969, n28968;
    wire [11:0]n9544;
    
    wire n28967, n28966, n28965, n28964, n27767, n28963, n28962, 
        n28961, n28960, n28959, n28958, n28957, n27883;
    wire [12:0]n9529;
    
    wire n28956, n28955, n28954, n27812, n28953, n28952, n28951, 
        n28950, n28949, n28948, n28947, n28946, n530_adj_4654, n603_adj_4655, 
        n676_adj_4656, n749_adj_4657, n822_adj_4658, n895_adj_4659, 
        n968_adj_4660, n27882, n27766, n1041_adj_4661, n1114_adj_4662, 
        n27811, n27765, n27810, n28945;
    wire [13:0]n9513;
    
    wire n28944, n28943, n27881, n27764, n27880, n27809, n27763, 
        n27808, n28942, n28941, n28940, n28939, n28938, n28937, 
        n27879, n27878, n95_adj_4664, n28936, n27762, n28935, n26_adj_4665, 
        n168_adj_4666, n241_adj_4667, n314_adj_4668, n387_adj_4669, 
        n460_adj_4670, n533_adj_4671, n606_adj_4672, n679_adj_4673, 
        n752_adj_4674, n825_adj_4675, n320_adj_4676, n28934, n247_adj_4677, 
        n28933, n27761, n27807, n174_adj_4678, n28932, n27806, n27805, 
        n32_adj_4679, n101_adj_4680, n27804, n27760;
    wire [14:0]n9496;
    
    wire n1120_adj_4682, n28931, n1047_adj_4683, n28930, n27803, n27759, 
        n974_adj_4684, n28929, n27951, n27950, n27802, n27949, n27758, 
        n901_adj_4688, n28928, n27801, n828_adj_4689, n28927, n755_adj_4690, 
        n28926, n682_adj_4691, n28925, n609_adj_4692, n28924, n536_adj_4693, 
        n28923, n27757, n463_adj_4695, n28922, n390_adj_4696, n28921, 
        n317_adj_4697, n28920, n244_adj_4698, n28919, n171_adj_4699, 
        n28918, n27948, n29_adj_4701, n98_adj_4702;
    wire [15:0]n9478;
    
    wire n28917, n1117_adj_4703, n28916, n1044_adj_4704, n28915, n971_adj_4705, 
        n28914, n898_adj_4706, n28913, n28912, n28911, n28910, n27800, 
        n28909, n28908, n28907, n28906, n28905, n28904, n28903;
    wire [16:0]n9459;
    
    wire n28902, n28901, n28900, n28899, n28898, n28897, n28896, 
        n28895, n28894, n28893, n28892, n28891, n28890, n28889, 
        n28888, n27947, n28887;
    wire [17:0]n9439;
    
    wire n28886, n28885, n28884, n28883, n28882, n28881, n28880, 
        n28879, n28878, n28877, n28876, n28875, n28874, n28873, 
        n28872, n28871, n28870;
    wire [18:0]n9418;
    
    wire n28869, n28868, n28867, n28866, n28865, n28864, n28863, 
        n28862, n28861, n28860, n28859, n28858, n28857, n28856, 
        n28855, n28854, n28853, n28852;
    wire [19:0]n9396;
    
    wire n28851, n28850, n28849, n28848, n28847, n28846, n28845, 
        n28844, n28843, n28842, n28841, n28840, n28839, n28838, 
        n28837, n28836, n28835, n28834, n27946, n28833, n28832, 
        n28831, n28830, n28829, n28828, n28827, n28826, n28825, 
        n28824, n28823, n28822, n28821, n28820, n28819, n28818, 
        n28817, n28816, n28815, n28814, n28813, n28812, n28811, 
        n28810, n28809, n28808, n28807, n28806, n28805, n28804, 
        n28803, n28802, n28801, n28800, n28799, n28798, n28797, 
        n28796, n28795, n27945, n28794, n28793, n28792, n28791, 
        n27450, n27944, n28790, n28789, n28788, n28787, n28786, 
        n28785, n28784, n28783, n28782, n28781, n28780, n27416, 
        n4_adj_4707, n27373;
    
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n27942), .I0(GND_net), .I1(n1_adj_4708[14]), 
            .CO(n27943));
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3609[1]), .I1(n257[1]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3584[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30915_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n37310));   // verilog/motorControl.v(29[14] 48[8])
    defparam i30915_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5203_11 (.CI(n28778), .I0(n9373[8]), .I1(n734), .CO(n28779));
    SB_LUT4 add_5203_10_lut (.I0(GND_net), .I1(n9373[7]), .I2(n661), .I3(n28777), 
            .O(n9349[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_10 (.CI(n28777), .I0(n9373[7]), .I1(n661), .CO(n28778));
    SB_LUT4 add_5203_9_lut (.I0(GND_net), .I1(n9373[6]), .I2(n588), .I3(n28776), 
            .O(n9349[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_9 (.CI(n28776), .I0(n9373[6]), .I1(n588), .CO(n28777));
    SB_LUT4 add_5203_8_lut (.I0(GND_net), .I1(n9373[5]), .I2(n515), .I3(n28775), 
            .O(n9349[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_8 (.CI(n28775), .I0(n9373[5]), .I1(n515), .CO(n28776));
    SB_LUT4 add_5203_7_lut (.I0(GND_net), .I1(n9373[4]), .I2(n442), .I3(n28774), 
            .O(n9349[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_7 (.CI(n28774), .I0(n9373[4]), .I1(n442), .CO(n28775));
    SB_LUT4 add_5203_6_lut (.I0(GND_net), .I1(n9373[3]), .I2(n369), .I3(n28773), 
            .O(n9349[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_6 (.CI(n28773), .I0(n9373[3]), .I1(n369), .CO(n28774));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[13]), 
            .I3(n27941), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5203_5_lut (.I0(GND_net), .I1(n9373[2]), .I2(n296), .I3(n28772), 
            .O(n9349[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19385_2_lut (.I0(n28[9]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19385_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19386_2_lut (.I0(n28[10]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19386_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n27941), .I0(GND_net), .I1(n1_adj_4708[13]), 
            .CO(n27942));
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19387_2_lut (.I0(n28[11]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19387_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5203_5 (.CI(n28772), .I0(n9373[2]), .I1(n296), .CO(n28773));
    SB_LUT4 add_5203_4_lut (.I0(GND_net), .I1(n9373[1]), .I2(n223), .I3(n28771), 
            .O(n9349[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19388_2_lut (.I0(n28[12]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19388_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5203_4 (.CI(n28771), .I0(n9373[1]), .I1(n223), .CO(n28772));
    SB_LUT4 add_5203_3_lut (.I0(GND_net), .I1(n9373[0]), .I2(n150), .I3(n28770), 
            .O(n9349[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_3 (.CI(n28770), .I0(n9373[0]), .I1(n150), .CO(n28771));
    SB_LUT4 add_5203_2_lut (.I0(GND_net), .I1(n8_adj_4290), .I2(n77), 
            .I3(GND_net), .O(n9349[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22776_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [18]), 
            .I2(n4_adj_4291), .I3(n9925[1]), .O(n6_adj_4292));   // verilog/motorControl.v(34[25:36])
    defparam i22776_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [18]), 
            .I2(n9925[1]), .I3(n4_adj_4291), .O(n9918[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1497 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [18]), 
            .I2(n9925[0]), .I3(n27505), .O(n9918[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1497.LUT_INIT = 16'h8778;
    SB_LUT4 i22768_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [18]), 
            .I2(n27505), .I3(n9925[0]), .O(n4_adj_4291));   // verilog/motorControl.v(34[25:36])
    defparam i22768_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_5203_2 (.CI(GND_net), .I0(n8_adj_4290), .I1(n77), .CO(n28770));
    SB_LUT4 i22757_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3509 [18]), .I3(\Ki[1] ), 
            .O(n27505));   // verilog/motorControl.v(34[25:36])
    defparam i22757_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3485[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i22755_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3509 [18]), .I3(\Ki[1] ), 
            .O(n9918[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22755_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[12]), 
            .I3(n27940), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n27940), .I0(GND_net), .I1(n1_adj_4708[12]), 
            .CO(n27941));
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19389_2_lut (.I0(n28[13]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19389_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4294));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[11]), 
            .I3(n27939), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4297));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4298));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4300));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22838_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [20]), 
            .I2(n27582), .I3(n9936[0]), .O(n4_adj_4301));   // verilog/motorControl.v(34[25:36])
    defparam i22838_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n27939), .I0(GND_net), .I1(n1_adj_4708[11]), 
            .CO(n27940));
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4303));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4304));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1498 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [20]), 
            .I2(n9936[0]), .I3(n27582), .O(n9931[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1498.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4306));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4307));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1499 (.I0(n62), .I1(n131), .I2(n9931[0]), 
            .I3(n204), .O(n9925[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1499.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22807_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n9931[0]), 
            .O(n4_adj_4309));   // verilog/motorControl.v(34[25:36])
    defparam i22807_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[10]), 
            .I3(n27938), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22825_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3509 [20]), .I3(\Ki[1] ), 
            .O(n9931[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22825_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n27938), .I0(GND_net), .I1(n1_adj_4708[10]), 
            .CO(n27939));
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4310));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19390_2_lut (.I0(n28[14]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19390_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4312));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22827_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3509 [20]), .I3(\Ki[1] ), 
            .O(n27582));   // verilog/motorControl.v(34[25:36])
    defparam i22827_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4313));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4315));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4316));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4317));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4318));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4319));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4320));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4321));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4322));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19391_2_lut (.I0(n28[15]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19391_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4324));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4325));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[9]), 
            .I3(n27937), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4327));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4328));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4330));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4292), .I1(\Ki[4] ), .I2(n9925[2]), .I3(\PID_CONTROLLER.integral_23__N_3509 [18]), 
            .O(n9918[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4331));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4333));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4334));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22848_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3509 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [21]), .O(n9936[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22848_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4336));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4337));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4339));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1500 (.I0(n4_adj_4309), .I1(\Ki[3] ), .I2(n9931[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [19]), .O(n9925[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1500.LUT_INIT = 16'h965a;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n27937), .I0(GND_net), .I1(n1_adj_4708[9]), 
            .CO(n27938));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[8]), 
            .I3(n27936), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1501 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3509 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [20]), .O(n12_adj_4340));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1501.LUT_INIT = 16'h9c50;
    SB_LUT4 i22784_4_lut (.I0(n9925[2]), .I1(\Ki[4] ), .I2(n6_adj_4292), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [18]), .O(n8_adj_4341));   // verilog/motorControl.v(34[25:36])
    defparam i22784_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3509 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [21]), .O(n11_adj_4342));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22815_4_lut (.I0(n9931[1]), .I1(\Ki[3] ), .I2(n4_adj_4309), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [19]), .O(n6_adj_4343));   // verilog/motorControl.v(34[25:36])
    defparam i22815_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i22850_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3509 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [21]), .O(n27607));   // verilog/motorControl.v(34[25:36])
    defparam i22850_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4343), .I1(n11_adj_4342), .I2(n8_adj_4341), 
            .I3(n12_adj_4340), .O(n18_adj_4344));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4345));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4346));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4347));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4348));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4349));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3509 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3509 [22]), .O(n13_adj_4350));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4350), .I1(n18_adj_4344), .I2(n27607), 
            .I3(n4_adj_4301), .O(n34839));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4351));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4352));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n27936), .I0(GND_net), .I1(n1_adj_4708[8]), 
            .CO(n27937));
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4353));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4354));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4355));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[7]), 
            .I3(n27935), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n27935), .I0(GND_net), .I1(n1_adj_4708[7]), 
            .CO(n27936));
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3609[23]), .I1(n257[23]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3584[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[6]), 
            .I3(n27934), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3609[22]), .I1(n257[22]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3584[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3609[21]), .I1(n257[21]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3584[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3609[20]), .I1(n257[20]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3584[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3609[19]), .I1(n257[19]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3584[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n27934), .I0(GND_net), .I1(n1_adj_4708[6]), 
            .CO(n27935));
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3609[18]), .I1(n257[18]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3584[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3609[17]), .I1(n257[17]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3584[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3609[16]), .I1(n257[16]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3584[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[5]), 
            .I3(n27933), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3609[15]), .I1(n257[15]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n27933), .I0(GND_net), .I1(n1_adj_4708[5]), 
            .CO(n27934));
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3584[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[4]), 
            .I3(n27932), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3609[14]), .I1(n257[14]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3584[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n27932), .I0(GND_net), .I1(n1_adj_4708[4]), 
            .CO(n27933));
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3609[13]), .I1(n257[13]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[3]), 
            .I3(n27931), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3584[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3609[12]), .I1(n257[12]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3584[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3609[11]), .I1(n257[11]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3584[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3609[10]), .I1(n257[10]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3584[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3609[9]), .I1(n257[9]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3584[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3609[8]), .I1(n257[8]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3584[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3609[7]), .I1(n257[7]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3584[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3609[6]), .I1(n257[6]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3584[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n27931), .I0(GND_net), .I1(n1_adj_4708[3]), 
            .CO(n27932));
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3609[5]), .I1(n257[5]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3584[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3609[4]), .I1(n257[4]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3584[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3609[3]), .I1(n257[3]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3584[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4360));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4361));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4363));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19392_2_lut (.I0(n28[16]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3609[2]), .I1(n257[2]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3584[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4364));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4365));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[2]), 
            .I3(n27930), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4367));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4368));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4370));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n28[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4373));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4374));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4375));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4376));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1502 (.I0(n6_adj_4377), .I1(\Kp[4] ), .I2(n9628[2]), 
            .I3(n28[18]), .O(n9621[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1502.LUT_INIT = 16'h965a;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n27930), .I0(GND_net), .I1(n1_adj_4708[2]), 
            .CO(n27931));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[1]), 
            .I3(n27929), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22726_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n9639[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22726_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i2_4_lut_adj_1503 (.I0(n4_adj_4380), .I1(\Kp[3] ), .I2(n9634[1]), 
            .I3(n28[19]), .O(n9628[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1503.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4382));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1504 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n28[23]), 
            .I3(n28[20]), .O(n12_adj_4385));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1504.LUT_INIT = 16'h9c50;
    SB_LUT4 i22662_4_lut (.I0(n9628[2]), .I1(\Kp[4] ), .I2(n6_adj_4377), 
            .I3(n28[18]), .O(n8_adj_4386));   // verilog/motorControl.v(34[16:22])
    defparam i22662_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1505 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n28[19]), 
            .I3(n28[21]), .O(n11_adj_4387));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut_adj_1505.LUT_INIT = 16'h6ca0;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n27929), .I0(GND_net), .I1(n1_adj_4708[1]), 
            .CO(n27930));
    SB_LUT4 i22693_4_lut (.I0(n9634[1]), .I1(\Kp[3] ), .I2(n4_adj_4380), 
            .I3(n28[19]), .O(n6_adj_4388));   // verilog/motorControl.v(34[16:22])
    defparam i22693_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4708[0]), 
            .CO(n27929));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n27928), .O(\PID_CONTROLLER.integral_23__N_3560 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22728_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n27475));   // verilog/motorControl.v(34[16:22])
    defparam i22728_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1506 (.I0(n6_adj_4388), .I1(n11_adj_4387), .I2(n8_adj_4386), 
            .I3(n12_adj_4385), .O(n18_adj_4389));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut_adj_1506.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1507 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n28[18]), 
            .I3(n28[22]), .O(n13_adj_4390));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut_adj_1507.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1508 (.I0(n13_adj_4390), .I1(n18_adj_4389), .I2(n27475), 
            .I3(n4_adj_4391), .O(n34155));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1508.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4394));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1[22]), .I3(n27927), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n27927), .I0(GND_net), .I1(n1[22]), 
            .CO(n27928));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1[21]), .I3(n27926), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n27926), .I0(GND_net), .I1(n1[21]), 
            .CO(n27927));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1[20]), .I3(n27925), .O(n41_adj_4395)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19393_2_lut (.I0(n28[17]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19393_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4397));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4398));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4399));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4401));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n27925), .I0(GND_net), .I1(n1[20]), 
            .CO(n27926));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1[19]), .I3(n27924), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n27924), .I0(GND_net), .I1(n1[19]), 
            .CO(n27925));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1[18]), .I3(n27923), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n27923), .I0(GND_net), .I1(n1[18]), 
            .CO(n27924));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1[17]), .I3(n27922), .O(n35_adj_4402)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n27922), .I0(GND_net), .I1(n1[17]), 
            .CO(n27923));
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4403));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4404));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4406));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4407));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4409));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4410));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1[16]), .I3(n27921), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4413));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n27921), .I0(GND_net), .I1(n1[16]), 
            .CO(n27922));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1[15]), .I3(n27920), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4414));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4416));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19394_2_lut (.I0(n28[18]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4418));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4419));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4420));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19395_2_lut (.I0(n28[19]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19395_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4421));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4422));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19396_2_lut (.I0(n28[20]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n27920), .I0(GND_net), .I1(n1[15]), 
            .CO(n27921));
    SB_LUT4 add_5241_7_lut (.I0(GND_net), .I1(n34839), .I2(n490), .I3(n29255), 
            .O(n9910[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5241_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5241_6_lut (.I0(GND_net), .I1(n9918[3]), .I2(n417), .I3(n29254), 
            .O(n9910[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5241_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5241_6 (.CI(n29254), .I0(n9918[3]), .I1(n417), .CO(n29255));
    SB_LUT4 add_5241_5_lut (.I0(GND_net), .I1(n9918[2]), .I2(n344), .I3(n29253), 
            .O(n9910[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5241_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5241_5 (.CI(n29253), .I0(n9918[2]), .I1(n344), .CO(n29254));
    SB_LUT4 add_5241_4_lut (.I0(GND_net), .I1(n9918[1]), .I2(n271_adj_4329), 
            .I3(n29252), .O(n9910[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5241_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5241_4 (.CI(n29252), .I0(n9918[1]), .I1(n271_adj_4329), 
            .CO(n29253));
    SB_LUT4 add_5241_3_lut (.I0(GND_net), .I1(n9918[0]), .I2(n198), .I3(n29251), 
            .O(n9910[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5241_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1[14]), .I3(n27919), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5241_3 (.CI(n29251), .I0(n9918[0]), .I1(n198), .CO(n29252));
    SB_LUT4 add_5241_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n9910[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5241_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5241_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n29251));
    SB_LUT4 add_5240_8_lut (.I0(GND_net), .I1(n9910[5]), .I2(n560), .I3(n29250), 
            .O(n9901[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5240_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5240_7_lut (.I0(GND_net), .I1(n9910[4]), .I2(n487), .I3(n29249), 
            .O(n9901[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5240_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5240_7 (.CI(n29249), .I0(n9910[4]), .I1(n487), .CO(n29250));
    SB_LUT4 add_5240_6_lut (.I0(GND_net), .I1(n9910[3]), .I2(n414), .I3(n29248), 
            .O(n9901[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5240_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5240_6 (.CI(n29248), .I0(n9910[3]), .I1(n414), .CO(n29249));
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4423));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4424));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4425));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4426));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4427));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5240_5_lut (.I0(GND_net), .I1(n9910[2]), .I2(n341), .I3(n29247), 
            .O(n9901[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5240_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5240_5 (.CI(n29247), .I0(n9910[2]), .I1(n341), .CO(n29248));
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4428));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5240_4_lut (.I0(GND_net), .I1(n9910[1]), .I2(n268_adj_4324), 
            .I3(n29246), .O(n9901[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5240_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5240_4 (.CI(n29246), .I0(n9910[1]), .I1(n268_adj_4324), 
            .CO(n29247));
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4429));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4430));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4433));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5240_3_lut (.I0(GND_net), .I1(n9910[0]), .I2(n195), .I3(n29245), 
            .O(n9901[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5240_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5240_3 (.CI(n29245), .I0(n9910[0]), .I1(n195), .CO(n29246));
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5240_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n9901[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5240_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5240_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n29245));
    SB_LUT4 add_5239_9_lut (.I0(GND_net), .I1(n9901[6]), .I2(n630), .I3(n29244), 
            .O(n9891[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19397_2_lut (.I0(n28[21]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19397_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5239_8_lut (.I0(GND_net), .I1(n9901[5]), .I2(n557), .I3(n29243), 
            .O(n9891[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5239_8 (.CI(n29243), .I0(n9901[5]), .I1(n557), .CO(n29244));
    SB_LUT4 add_5239_7_lut (.I0(GND_net), .I1(n9901[4]), .I2(n484), .I3(n29242), 
            .O(n9891[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5239_7 (.CI(n29242), .I0(n9901[4]), .I1(n484), .CO(n29243));
    SB_LUT4 add_5239_6_lut (.I0(GND_net), .I1(n9901[3]), .I2(n411), .I3(n29241), 
            .O(n9891[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n27919), .I0(GND_net), .I1(n1[14]), 
            .CO(n27920));
    SB_CARRY add_5239_6 (.CI(n29241), .I0(n9901[3]), .I1(n411), .CO(n29242));
    SB_LUT4 add_5239_5_lut (.I0(GND_net), .I1(n9901[2]), .I2(n338), .I3(n29240), 
            .O(n9891[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5239_5 (.CI(n29240), .I0(n9901[2]), .I1(n338), .CO(n29241));
    SB_LUT4 add_5239_4_lut (.I0(GND_net), .I1(n9901[1]), .I2(n265), .I3(n29239), 
            .O(n9891[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5239_4 (.CI(n29239), .I0(n9901[1]), .I1(n265), .CO(n29240));
    SB_LUT4 add_5239_3_lut (.I0(GND_net), .I1(n9901[0]), .I2(n192), .I3(n29238), 
            .O(n9891[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5239_3 (.CI(n29238), .I0(n9901[0]), .I1(n192), .CO(n29239));
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5239_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n9891[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5239_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5239_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n29238));
    SB_LUT4 add_5238_10_lut (.I0(GND_net), .I1(n9891[7]), .I2(n700), .I3(n29237), 
            .O(n9880[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5238_9_lut (.I0(GND_net), .I1(n9891[6]), .I2(n627), .I3(n29236), 
            .O(n9880[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5238_9 (.CI(n29236), .I0(n9891[6]), .I1(n627), .CO(n29237));
    SB_LUT4 add_5238_8_lut (.I0(GND_net), .I1(n9891[5]), .I2(n554), .I3(n29235), 
            .O(n9880[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5238_8 (.CI(n29235), .I0(n9891[5]), .I1(n554), .CO(n29236));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1[13]), .I3(n27918), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n27918), .I0(GND_net), .I1(n1[13]), 
            .CO(n27919));
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19398_2_lut (.I0(n28[22]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4434));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4435));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4436));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5238_7_lut (.I0(GND_net), .I1(n9891[4]), .I2(n481), .I3(n29234), 
            .O(n9880[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29775_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n36171));
    defparam i29775_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i29772_3_lut (.I0(n11_adj_4436), .I1(n9_adj_4435), .I2(n36171), 
            .I3(GND_net), .O(n36168));
    defparam i29772_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_264_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n38226));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_264_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30137_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n38226), 
            .I2(IntegralLimit[7]), .I3(n36168), .O(n36534));
    defparam i30137_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i30031_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4434), 
            .I2(IntegralLimit[9]), .I3(n36534), .O(n36428));
    defparam i30031_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_246_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n38208));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_246_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30029_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4434), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4435), .O(n36426));
    defparam i30029_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30027_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n38208), 
            .I2(IntegralLimit[11]), .I3(n36426), .O(n36424));
    defparam i30027_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_239_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n38201));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_239_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4438));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29721_4_lut (.I0(n27), .I1(n15_adj_4439), .I2(n13_adj_4440), 
            .I3(n11_adj_4441), .O(n36117));
    defparam i29721_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29727_4_lut (.I0(n21_adj_4442), .I1(n19_adj_4443), .I2(n17_adj_4444), 
            .I3(n9_adj_4445), .O(n36123));
    defparam i29727_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_831_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3609[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4446));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3609[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4447));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3609[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4448));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3609[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4449));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4450));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 duty_23__I_831_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3609[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4452));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_831_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3609[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4453));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3609[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4454));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3609[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4455));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3609[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4456));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3609[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4457));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29705_2_lut (.I0(n43), .I1(n19_adj_4443), .I2(GND_net), .I3(GND_net), 
            .O(n36101));
    defparam i29705_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5238_7 (.CI(n29234), .I0(n9891[4]), .I1(n481), .CO(n29235));
    SB_LUT4 duty_23__I_831_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3609[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4458));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5238_6_lut (.I0(GND_net), .I1(n9891[3]), .I2(n408), .I3(n29233), 
            .O(n9880[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5238_6 (.CI(n29233), .I0(n9891[3]), .I1(n408), .CO(n29234));
    SB_LUT4 duty_23__I_831_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3609[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4459));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5238_5_lut (.I0(GND_net), .I1(n9891[2]), .I2(n335), .I3(n29232), 
            .O(n9880[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3609[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4460));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5238_5 (.CI(n29232), .I0(n9891[2]), .I1(n335), .CO(n29233));
    SB_LUT4 duty_23__I_831_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3609[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4461));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5238_4_lut (.I0(GND_net), .I1(n9891[1]), .I2(n262), .I3(n29231), 
            .O(n9880[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3609[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4462));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i33_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5238_4 (.CI(n29231), .I0(n9891[1]), .I1(n262), .CO(n29232));
    SB_LUT4 duty_23__I_831_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3609[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4463));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5238_3_lut (.I0(GND_net), .I1(n9891[0]), .I2(n189), .I3(n29230), 
            .O(n9880[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3609[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4464));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5238_3 (.CI(n29230), .I0(n9891[0]), .I1(n189), .CO(n29231));
    SB_LUT4 duty_23__I_831_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3609[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4465));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5238_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n9880[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5238_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3609[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4466));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i21_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5238_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n29230));
    SB_LUT4 add_5237_11_lut (.I0(GND_net), .I1(n9880[8]), .I2(n770), .I3(n29229), 
            .O(n9868[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29692_4_lut (.I0(n21_adj_4466), .I1(n19_adj_4465), .I2(n17_adj_4464), 
            .I3(n9_adj_4463), .O(n36088));
    defparam i29692_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5237_10_lut (.I0(GND_net), .I1(n9880[7]), .I2(n697), .I3(n29228), 
            .O(n9868[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29686_4_lut (.I0(n27_adj_4461), .I1(n15_adj_4460), .I2(n13_adj_4459), 
            .I3(n11_adj_4458), .O(n36082));
    defparam i29686_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5237_10 (.CI(n29228), .I0(n9880[7]), .I1(n697), .CO(n29229));
    SB_LUT4 duty_23__I_831_i12_3_lut (.I0(duty_23__N_3609[7]), .I1(duty_23__N_3609[16]), 
            .I2(n33_adj_4462), .I3(GND_net), .O(n12_adj_4467));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5237_9_lut (.I0(GND_net), .I1(n9880[6]), .I2(n624), .I3(n29227), 
            .O(n9868[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_9 (.CI(n29227), .I0(n9880[6]), .I1(n624), .CO(n29228));
    SB_LUT4 duty_23__I_831_i10_3_lut (.I0(duty_23__N_3609[5]), .I1(duty_23__N_3609[6]), 
            .I2(n13_adj_4459), .I3(GND_net), .O(n10_adj_4468));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5237_8_lut (.I0(GND_net), .I1(n9880[5]), .I2(n551), .I3(n29226), 
            .O(n9868[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i30_3_lut (.I0(n12_adj_4467), .I1(duty_23__N_3609[17]), 
            .I2(n35_adj_4457), .I3(GND_net), .O(n30));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5237_8 (.CI(n29226), .I0(n9880[5]), .I1(n551), .CO(n29227));
    SB_LUT4 add_5237_7_lut (.I0(GND_net), .I1(n9880[4]), .I2(n478), .I3(n29225), 
            .O(n9868[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29965_4_lut (.I0(n13_adj_4459), .I1(n11_adj_4458), .I2(n9_adj_4463), 
            .I3(n36099), .O(n36362));
    defparam i29965_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5237_7 (.CI(n29225), .I0(n9880[4]), .I1(n478), .CO(n29226));
    SB_LUT4 i29961_4_lut (.I0(n19_adj_4465), .I1(n17_adj_4464), .I2(n15_adj_4460), 
            .I3(n36362), .O(n36358));
    defparam i29961_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_5237_6_lut (.I0(GND_net), .I1(n9880[3]), .I2(n405), .I3(n29224), 
            .O(n9868[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30260_4_lut (.I0(n25_adj_4455), .I1(n23_adj_4454), .I2(n21_adj_4466), 
            .I3(n36358), .O(n36657));
    defparam i30260_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_5237_6 (.CI(n29224), .I0(n9880[3]), .I1(n405), .CO(n29225));
    SB_LUT4 add_5237_5_lut (.I0(GND_net), .I1(n9880[2]), .I2(n332), .I3(n29223), 
            .O(n9868[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30099_4_lut (.I0(n31_adj_4453), .I1(n29_adj_4452), .I2(n27_adj_4461), 
            .I3(n36657), .O(n36496));
    defparam i30099_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_5237_5 (.CI(n29223), .I0(n9880[2]), .I1(n332), .CO(n29224));
    SB_LUT4 i30322_4_lut (.I0(n37_adj_4456), .I1(n35_adj_4457), .I2(n33_adj_4462), 
            .I3(n36496), .O(n36719));
    defparam i30322_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5237_4_lut (.I0(GND_net), .I1(n9880[1]), .I2(n259), .I3(n29222), 
            .O(n9868[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i16_3_lut (.I0(duty_23__N_3609[9]), .I1(duty_23__N_3609[21]), 
            .I2(n43_adj_4449), .I3(GND_net), .O(n16_adj_4469));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5237_4 (.CI(n29222), .I0(n9880[1]), .I1(n259), .CO(n29223));
    SB_LUT4 add_5237_3_lut (.I0(GND_net), .I1(n9880[0]), .I2(n186), .I3(n29221), 
            .O(n9868[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30236_3_lut (.I0(n6_adj_4470), .I1(duty_23__N_3609[10]), .I2(n21_adj_4466), 
            .I3(GND_net), .O(n36633));   // verilog/motorControl.v(36[10:25])
    defparam i30236_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5237_3 (.CI(n29221), .I0(n9880[0]), .I1(n186), .CO(n29222));
    SB_LUT4 i30237_3_lut (.I0(n36633), .I1(duty_23__N_3609[11]), .I2(n23_adj_4454), 
            .I3(GND_net), .O(n36634));   // verilog/motorControl.v(36[10:25])
    defparam i30237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5237_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n9868[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5237_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5237_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n29221));
    SB_LUT4 duty_23__I_831_i8_3_lut (.I0(duty_23__N_3609[4]), .I1(duty_23__N_3609[8]), 
            .I2(n17_adj_4464), .I3(GND_net), .O(n8_adj_4471));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5236_12_lut (.I0(GND_net), .I1(n9868[9]), .I2(n840), .I3(n29220), 
            .O(n9855[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i24_3_lut (.I0(n16_adj_4469), .I1(duty_23__N_3609[22]), 
            .I2(n45_adj_4448), .I3(GND_net), .O(n24_adj_4472));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5236_11_lut (.I0(GND_net), .I1(n9868[8]), .I2(n767), .I3(n29219), 
            .O(n9855[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29671_4_lut (.I0(n43_adj_4449), .I1(n25_adj_4455), .I2(n23_adj_4454), 
            .I3(n36088), .O(n36067));
    defparam i29671_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30143_4_lut (.I0(n24_adj_4472), .I1(n8_adj_4471), .I2(n45_adj_4448), 
            .I3(n36065), .O(n36540));   // verilog/motorControl.v(36[10:25])
    defparam i30143_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5236_11 (.CI(n29219), .I0(n9868[8]), .I1(n767), .CO(n29220));
    SB_LUT4 i30194_3_lut (.I0(n36634), .I1(duty_23__N_3609[12]), .I2(n25_adj_4455), 
            .I3(GND_net), .O(n36591));   // verilog/motorControl.v(36[10:25])
    defparam i30194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i4_4_lut (.I0(duty_23__N_3609[0]), .I1(duty_23__N_3609[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4473));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 add_5236_10_lut (.I0(GND_net), .I1(n9868[7]), .I2(n694), .I3(n29218), 
            .O(n9855[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30234_3_lut (.I0(n4_adj_4473), .I1(duty_23__N_3609[13]), .I2(n27_adj_4461), 
            .I3(GND_net), .O(n36631));   // verilog/motorControl.v(36[10:25])
    defparam i30234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30235_3_lut (.I0(n36631), .I1(duty_23__N_3609[14]), .I2(n29_adj_4452), 
            .I3(GND_net), .O(n36632));   // verilog/motorControl.v(36[10:25])
    defparam i30235_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5236_10 (.CI(n29218), .I0(n9868[7]), .I1(n694), .CO(n29219));
    SB_LUT4 i29681_4_lut (.I0(n33_adj_4462), .I1(n31_adj_4453), .I2(n29_adj_4452), 
            .I3(n36082), .O(n36077));
    defparam i29681_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30332_4_lut (.I0(n30), .I1(n10_adj_4468), .I2(n35_adj_4457), 
            .I3(n36075), .O(n36729));   // verilog/motorControl.v(36[10:25])
    defparam i30332_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30196_3_lut (.I0(n36632), .I1(duty_23__N_3609[15]), .I2(n31_adj_4453), 
            .I3(GND_net), .O(n36593));   // verilog/motorControl.v(36[10:25])
    defparam i30196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30383_4_lut (.I0(n36593), .I1(n36729), .I2(n35_adj_4457), 
            .I3(n36077), .O(n36780));   // verilog/motorControl.v(36[10:25])
    defparam i30383_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30384_3_lut (.I0(n36780), .I1(duty_23__N_3609[18]), .I2(n37_adj_4456), 
            .I3(GND_net), .O(n36781));   // verilog/motorControl.v(36[10:25])
    defparam i30384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30363_3_lut (.I0(n36781), .I1(duty_23__N_3609[19]), .I2(n39_adj_4446), 
            .I3(GND_net), .O(n36760));   // verilog/motorControl.v(36[10:25])
    defparam i30363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29673_4_lut (.I0(n43_adj_4449), .I1(n41_adj_4447), .I2(n39_adj_4446), 
            .I3(n36719), .O(n36069));
    defparam i29673_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30294_4_lut (.I0(n36591), .I1(n36540), .I2(n45_adj_4448), 
            .I3(n36067), .O(n36691));   // verilog/motorControl.v(36[10:25])
    defparam i30294_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4444), .I3(GND_net), 
            .O(n8_adj_4474));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i30353_3_lut (.I0(n36760), .I1(duty_23__N_3609[20]), .I2(n41_adj_4447), 
            .I3(GND_net), .O(n40));   // verilog/motorControl.v(36[10:25])
    defparam i30353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30296_4_lut (.I0(n40), .I1(n36691), .I2(n45_adj_4448), .I3(n36069), 
            .O(n36693));   // verilog/motorControl.v(36[10:25])
    defparam i30296_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30297_3_lut (.I0(n36693), .I1(PWMLimit[23]), .I2(duty_23__N_3609[23]), 
            .I3(GND_net), .O(duty_23__N_3608));   // verilog/motorControl.v(36[10:25])
    defparam i30297_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3609[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4475));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3609[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4476));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3609[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4477));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3609[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4478));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3609[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4479));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3609[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4480));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3609[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4481));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3609[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4482));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3609[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4483));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3609[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4484));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3609[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4485));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5236_9_lut (.I0(GND_net), .I1(n9868[6]), .I2(n621), .I3(n29217), 
            .O(n9855[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_9 (.CI(n29217), .I0(n9868[6]), .I1(n621), .CO(n29218));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1[12]), .I3(n27917), .O(n25_adj_4486)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5236_8_lut (.I0(GND_net), .I1(n9868[5]), .I2(n548), .I3(n29216), 
            .O(n9855[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_8 (.CI(n29216), .I0(n9868[5]), .I1(n548), .CO(n29217));
    SB_LUT4 add_5236_7_lut (.I0(GND_net), .I1(n9868[4]), .I2(n475), .I3(n29215), 
            .O(n9855[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3609[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4487));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3609[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4488));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3609[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4489));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3609[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4490));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3609[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4491));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3609[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4492));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3609[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4493));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3609[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4494));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29655_4_lut (.I0(n21_adj_4494), .I1(n19_adj_4493), .I2(n17_adj_4492), 
            .I3(n9_adj_4491), .O(n36051));
    defparam i29655_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29649_4_lut (.I0(n27_adj_4490), .I1(n15_adj_4489), .I2(n13_adj_4488), 
            .I3(n11_adj_4487), .O(n36045));
    defparam i29649_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4485), 
            .I3(GND_net), .O(n12_adj_4495));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4488), 
            .I3(GND_net), .O(n10_adj_4496));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4495), .I1(n257[17]), .I2(n35_adj_4484), 
            .I3(GND_net), .O(n30_adj_4497));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29933_4_lut (.I0(n13_adj_4488), .I1(n11_adj_4487), .I2(n9_adj_4491), 
            .I3(n36063), .O(n36330));
    defparam i29933_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29929_4_lut (.I0(n19_adj_4493), .I1(n17_adj_4492), .I2(n15_adj_4489), 
            .I3(n36330), .O(n36326));
    defparam i29929_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i30252_4_lut (.I0(n25_adj_4478), .I1(n23_adj_4477), .I2(n21_adj_4494), 
            .I3(n36326), .O(n36649));
    defparam i30252_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30083_4_lut (.I0(n31_adj_4483), .I1(n29_adj_4482), .I2(n27_adj_4490), 
            .I3(n36649), .O(n36480));
    defparam i30083_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30320_4_lut (.I0(n37_adj_4481), .I1(n35_adj_4484), .I2(n33_adj_4485), 
            .I3(n36480), .O(n36717));
    defparam i30320_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4480), 
            .I3(GND_net), .O(n16_adj_4498));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30230_3_lut (.I0(n6_adj_4499), .I1(n257[10]), .I2(n21_adj_4494), 
            .I3(GND_net), .O(n36627));   // verilog/motorControl.v(38[19:35])
    defparam i30230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30231_3_lut (.I0(n36627), .I1(n257[11]), .I2(n23_adj_4477), 
            .I3(GND_net), .O(n36628));   // verilog/motorControl.v(38[19:35])
    defparam i30231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4492), 
            .I3(GND_net), .O(n8_adj_4500));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18936_2_lut (.I0(n28[0]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i18936_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4502));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5236_7 (.CI(n29215), .I0(n9868[4]), .I1(n475), .CO(n29216));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4450), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4503));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_5236_6_lut (.I0(GND_net), .I1(n9868[3]), .I2(n402), .I3(n29214), 
            .O(n9855[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_6 (.CI(n29214), .I0(n9868[3]), .I1(n402), .CO(n29215));
    SB_LUT4 add_5236_5_lut (.I0(GND_net), .I1(n9868[2]), .I2(n329), .I3(n29213), 
            .O(n9855[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_5 (.CI(n29213), .I0(n9868[2]), .I1(n329), .CO(n29214));
    SB_LUT4 add_5236_4_lut (.I0(GND_net), .I1(n9868[1]), .I2(n256_adj_4294), 
            .I3(n29212), .O(n9855[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4498), .I1(n257[22]), .I2(n45_adj_4479), 
            .I3(GND_net), .O(n24_adj_4504));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29633_4_lut (.I0(n43_adj_4480), .I1(n25_adj_4478), .I2(n23_adj_4477), 
            .I3(n36051), .O(n36029));
    defparam i29633_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30145_4_lut (.I0(n24_adj_4504), .I1(n8_adj_4500), .I2(n45_adj_4479), 
            .I3(n36027), .O(n36542));   // verilog/motorControl.v(38[19:35])
    defparam i30145_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30200_3_lut (.I0(n36628), .I1(n257[12]), .I2(n25_adj_4478), 
            .I3(GND_net), .O(n36597));   // verilog/motorControl.v(38[19:35])
    defparam i30200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3609[0]), .I1(n257[1]), 
            .I2(duty_23__N_3609[1]), .I3(n257[0]), .O(n4_adj_4505));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i30228_3_lut (.I0(n4_adj_4505), .I1(n257[13]), .I2(n27_adj_4490), 
            .I3(GND_net), .O(n36625));   // verilog/motorControl.v(38[19:35])
    defparam i30228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30229_3_lut (.I0(n36625), .I1(n257[14]), .I2(n29_adj_4482), 
            .I3(GND_net), .O(n36626));   // verilog/motorControl.v(38[19:35])
    defparam i30229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29645_4_lut (.I0(n33_adj_4485), .I1(n31_adj_4483), .I2(n29_adj_4482), 
            .I3(n36045), .O(n36041));
    defparam i29645_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30334_4_lut (.I0(n30_adj_4497), .I1(n10_adj_4496), .I2(n35_adj_4484), 
            .I3(n36039), .O(n36731));   // verilog/motorControl.v(38[19:35])
    defparam i30334_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30202_3_lut (.I0(n36626), .I1(n257[15]), .I2(n31_adj_4483), 
            .I3(GND_net), .O(n36599));   // verilog/motorControl.v(38[19:35])
    defparam i30202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30385_4_lut (.I0(n36599), .I1(n36731), .I2(n35_adj_4484), 
            .I3(n36041), .O(n36782));   // verilog/motorControl.v(38[19:35])
    defparam i30385_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30386_3_lut (.I0(n36782), .I1(n257[18]), .I2(n37_adj_4481), 
            .I3(GND_net), .O(n36783));   // verilog/motorControl.v(38[19:35])
    defparam i30386_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30361_3_lut (.I0(n36783), .I1(n257[19]), .I2(n39_adj_4476), 
            .I3(GND_net), .O(n36758));   // verilog/motorControl.v(38[19:35])
    defparam i30361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29635_4_lut (.I0(n43_adj_4480), .I1(n41_adj_4475), .I2(n39_adj_4476), 
            .I3(n36717), .O(n36031));
    defparam i29635_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30300_4_lut (.I0(n36597), .I1(n36542), .I2(n45_adj_4479), 
            .I3(n36029), .O(n36697));   // verilog/motorControl.v(38[19:35])
    defparam i30300_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30355_3_lut (.I0(n36758), .I1(n257[20]), .I2(n41_adj_4475), 
            .I3(GND_net), .O(n40_adj_4506));   // verilog/motorControl.v(38[19:35])
    defparam i30355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30302_4_lut (.I0(n40_adj_4506), .I1(n36697), .I2(n45_adj_4479), 
            .I3(n36031), .O(n36699));   // verilog/motorControl.v(38[19:35])
    defparam i30302_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30303_3_lut (.I0(n36699), .I1(duty_23__N_3609[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(38[19:35])
    defparam i30303_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3609[0]), .I1(n257[0]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3584[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3584[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3608), .I3(GND_net), .O(duty_23__N_3485[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5236_4 (.CI(n29212), .I0(n9868[1]), .I1(n256_adj_4294), 
            .CO(n29213));
    SB_LUT4 add_5236_3_lut (.I0(GND_net), .I1(n9868[0]), .I2(n183), .I3(n29211), 
            .O(n9855[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29738_2_lut (.I0(n7_adj_4507), .I1(n5_adj_4508), .I2(GND_net), 
            .I3(GND_net), .O(n36134));
    defparam i29738_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_5236_3 (.CI(n29211), .I0(n9868[0]), .I1(n183), .CO(n29212));
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5236_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n9855[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5236_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5236_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n29211));
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3485[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5235_13_lut (.I0(GND_net), .I1(n9855[10]), .I2(n910), 
            .I3(n29210), .O(n9841[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29997_4_lut (.I0(n13_adj_4440), .I1(n11_adj_4441), .I2(n9_adj_4445), 
            .I3(n36134), .O(n36394));
    defparam i29997_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5235_12_lut (.I0(GND_net), .I1(n9855[9]), .I2(n837), .I3(n29209), 
            .O(n9841[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n27917), .I0(GND_net), .I1(n1[12]), 
            .CO(n27918));
    SB_CARRY add_5235_12 (.CI(n29209), .I0(n9855[9]), .I1(n837), .CO(n29210));
    SB_LUT4 add_5235_11_lut (.I0(GND_net), .I1(n9855[8]), .I2(n764), .I3(n29208), 
            .O(n9841[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5235_11 (.CI(n29208), .I0(n9855[8]), .I1(n764), .CO(n29209));
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1[11]), .I3(n27916), .O(n23_adj_4509)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5235_10_lut (.I0(GND_net), .I1(n9855[7]), .I2(n691), .I3(n29207), 
            .O(n9841[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_10 (.CI(n29207), .I0(n9855[7]), .I1(n691), .CO(n29208));
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5235_9_lut (.I0(GND_net), .I1(n9855[6]), .I2(n618), .I3(n29206), 
            .O(n9841[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_9 (.CI(n29206), .I0(n9855[6]), .I1(n618), .CO(n29207));
    SB_LUT4 add_5235_8_lut (.I0(GND_net), .I1(n9855[5]), .I2(n545_adj_4510), 
            .I3(n29205), .O(n9841[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_8 (.CI(n29205), .I0(n9855[5]), .I1(n545_adj_4510), 
            .CO(n29206));
    SB_LUT4 add_5235_7_lut (.I0(GND_net), .I1(n9855[4]), .I2(n472_adj_4511), 
            .I3(n29204), .O(n9841[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_7 (.CI(n29204), .I0(n9855[4]), .I1(n472_adj_4511), 
            .CO(n29205));
    SB_LUT4 add_5235_6_lut (.I0(GND_net), .I1(n9855[3]), .I2(n399_adj_4512), 
            .I3(n29203), .O(n9841[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_6 (.CI(n29203), .I0(n9855[3]), .I1(n399_adj_4512), 
            .CO(n29204));
    SB_LUT4 add_5235_5_lut (.I0(GND_net), .I1(n9855[2]), .I2(n326_adj_4513), 
            .I3(n29202), .O(n9841[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_5 (.CI(n29202), .I0(n9855[2]), .I1(n326_adj_4513), 
            .CO(n29203));
    SB_LUT4 add_5235_4_lut (.I0(GND_net), .I1(n9855[1]), .I2(n253_adj_4514), 
            .I3(n29201), .O(n9841[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_4 (.CI(n29201), .I0(n9855[1]), .I1(n253_adj_4514), 
            .CO(n29202));
    SB_LUT4 add_5235_3_lut (.I0(GND_net), .I1(n9855[0]), .I2(n180_adj_4515), 
            .I3(n29200), .O(n9841[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5235_3 (.CI(n29200), .I0(n9855[0]), .I1(n180_adj_4515), 
            .CO(n29201));
    SB_CARRY unary_minus_5_add_3_13 (.CI(n27916), .I0(GND_net), .I1(n1[11]), 
            .CO(n27917));
    SB_LUT4 add_5235_2_lut (.I0(GND_net), .I1(n38_adj_4516), .I2(n107_adj_4517), 
            .I3(GND_net), .O(n9841[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5235_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5235_2 (.CI(GND_net), .I0(n38_adj_4516), .I1(n107_adj_4517), 
            .CO(n29200));
    SB_LUT4 add_5234_14_lut (.I0(GND_net), .I1(n9841[11]), .I2(n980_adj_4518), 
            .I3(n29199), .O(n9826[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5234_13_lut (.I0(GND_net), .I1(n9841[10]), .I2(n907_adj_4519), 
            .I3(n29198), .O(n9826[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_13 (.CI(n29198), .I0(n9841[10]), .I1(n907_adj_4519), 
            .CO(n29199));
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5234_12_lut (.I0(GND_net), .I1(n9841[9]), .I2(n834_adj_4520), 
            .I3(n29197), .O(n9826[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1[10]), .I3(n27915), .O(n21_adj_4442)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29993_4_lut (.I0(n19_adj_4443), .I1(n17_adj_4444), .I2(n15_adj_4439), 
            .I3(n36394), .O(n36390));
    defparam i29993_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n27915), .I0(GND_net), .I1(n1[10]), 
            .CO(n27916));
    SB_CARRY add_5234_12 (.CI(n29197), .I0(n9841[9]), .I1(n834_adj_4520), 
            .CO(n29198));
    SB_LUT4 add_5234_11_lut (.I0(GND_net), .I1(n9841[8]), .I2(n761_adj_4522), 
            .I3(n29196), .O(n9826[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1[9]), .I3(n27914), .O(n19_adj_4443)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4290));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5234_11 (.CI(n29196), .I0(n9841[8]), .I1(n761_adj_4522), 
            .CO(n29197));
    SB_LUT4 add_5234_10_lut (.I0(GND_net), .I1(n9841[7]), .I2(n688_adj_4524), 
            .I3(n29195), .O(n9826[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_10 (.CI(n29195), .I0(n9841[7]), .I1(n688_adj_4524), 
            .CO(n29196));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n27914), .I0(GND_net), .I1(n1[9]), 
            .CO(n27915));
    SB_LUT4 add_5234_9_lut (.I0(GND_net), .I1(n9841[6]), .I2(n615_adj_4525), 
            .I3(n29194), .O(n9826[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_9 (.CI(n29194), .I0(n9841[6]), .I1(n615_adj_4525), 
            .CO(n29195));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1[8]), .I3(n27913), .O(n17_adj_4444)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5234_8_lut (.I0(GND_net), .I1(n9841[5]), .I2(n542_adj_4527), 
            .I3(n29193), .O(n9826[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_8 (.CI(n29193), .I0(n9841[5]), .I1(n542_adj_4527), 
            .CO(n29194));
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n27913), .I0(GND_net), .I1(n1[8]), 
            .CO(n27914));
    SB_LUT4 add_5234_7_lut (.I0(GND_net), .I1(n9841[4]), .I2(n469_adj_4528), 
            .I3(n29192), .O(n9826[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1[7]), .I3(n27912), .O(n15_adj_4439)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5234_7 (.CI(n29192), .I0(n9841[4]), .I1(n469_adj_4528), 
            .CO(n29193));
    SB_LUT4 add_5234_6_lut (.I0(GND_net), .I1(n9841[3]), .I2(n396_adj_4530), 
            .I3(n29191), .O(n9826[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_6 (.CI(n29191), .I0(n9841[3]), .I1(n396_adj_4530), 
            .CO(n29192));
    SB_LUT4 add_5234_5_lut (.I0(GND_net), .I1(n9841[2]), .I2(n323_adj_4531), 
            .I3(n29190), .O(n9826[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n27912), .I0(GND_net), .I1(n1[7]), 
            .CO(n27913));
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4532));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5234_5 (.CI(n29190), .I0(n9841[2]), .I1(n323_adj_4531), 
            .CO(n29191));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1[6]), .I3(n27911), .O(n13_adj_4440)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5234_4_lut (.I0(GND_net), .I1(n9841[1]), .I2(n250_adj_4534), 
            .I3(n29189), .O(n9826[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n8060[0]), .I2(n8064[0]), 
            .I3(n27779), .O(duty_23__N_3609[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_4 (.CI(n29189), .I0(n9841[1]), .I1(n250_adj_4534), 
            .CO(n29190));
    SB_LUT4 add_5234_3_lut (.I0(GND_net), .I1(n9841[0]), .I2(n177_adj_4535), 
            .I3(n29188), .O(n9826[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_3 (.CI(n29188), .I0(n9841[0]), .I1(n177_adj_4535), 
            .CO(n29189));
    SB_LUT4 add_5234_2_lut (.I0(GND_net), .I1(n35_adj_4536), .I2(n104_adj_4537), 
            .I3(GND_net), .O(n9826[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n27911), .I0(GND_net), .I1(n1[6]), 
            .CO(n27912));
    SB_CARRY add_5234_2 (.CI(GND_net), .I0(n35_adj_4536), .I1(n104_adj_4537), 
            .CO(n29188));
    SB_LUT4 add_5233_15_lut (.I0(GND_net), .I1(n9826[12]), .I2(n1050_adj_4538), 
            .I3(n29187), .O(n9810[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30268_4_lut (.I0(n25_adj_4486), .I1(n23_adj_4509), .I2(n21_adj_4442), 
            .I3(n36390), .O(n36665));
    defparam i30268_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5233_14_lut (.I0(GND_net), .I1(n9826[11]), .I2(n977_adj_4539), 
            .I3(n29186), .O(n9810[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1[5]), .I3(n27910), .O(n11_adj_4441)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n27910), .I0(GND_net), .I1(n1[5]), 
            .CO(n27911));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1[4]), .I3(n27909), .O(n9_adj_4445)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n27778), .O(duty_23__N_3609[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30115_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n36665), 
            .O(n36512));
    defparam i30115_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY add_12_24 (.CI(n27778), .I0(n106[22]), .I1(n155[22]), .CO(n27779));
    SB_CARRY unary_minus_5_add_3_6 (.CI(n27909), .I0(GND_net), .I1(n1[4]), 
            .CO(n27910));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1[3]), .I3(n27908), .O(n7_adj_4507)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n27908), .I0(GND_net), .I1(n1[3]), 
            .CO(n27909));
    SB_CARRY add_5233_14 (.CI(n29186), .I0(n9826[11]), .I1(n977_adj_4539), 
            .CO(n29187));
    SB_LUT4 add_5233_13_lut (.I0(GND_net), .I1(n9826[10]), .I2(n904_adj_4543), 
            .I3(n29185), .O(n9810[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_13 (.CI(n29185), .I0(n9826[10]), .I1(n904_adj_4543), 
            .CO(n29186));
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5233_12_lut (.I0(GND_net), .I1(n9826[9]), .I2(n831_adj_4544), 
            .I3(n29184), .O(n9810[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_12 (.CI(n29184), .I0(n9826[9]), .I1(n831_adj_4544), 
            .CO(n29185));
    SB_LUT4 add_5233_11_lut (.I0(GND_net), .I1(n9826[8]), .I2(n758_adj_4545), 
            .I3(n29183), .O(n9810[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_11 (.CI(n29183), .I0(n9826[8]), .I1(n758_adj_4545), 
            .CO(n29184));
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5233_10_lut (.I0(GND_net), .I1(n9826[7]), .I2(n685_adj_4546), 
            .I3(n29182), .O(n9810[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5233_10 (.CI(n29182), .I0(n9826[7]), .I1(n685_adj_4546), 
            .CO(n29183));
    SB_LUT4 i30324_4_lut (.I0(n37), .I1(n35_adj_4402), .I2(n33), .I3(n36512), 
            .O(n36721));
    defparam i30324_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_5233_9_lut (.I0(GND_net), .I1(n9826[6]), .I2(n612_adj_4547), 
            .I3(n29181), .O(n9810[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_9 (.CI(n29181), .I0(n9826[6]), .I1(n612_adj_4547), 
            .CO(n29182));
    SB_LUT4 add_5233_8_lut (.I0(GND_net), .I1(n9826[5]), .I2(n539_adj_4548), 
            .I3(n29180), .O(n9810[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_8 (.CI(n29180), .I0(n9826[5]), .I1(n539_adj_4548), 
            .CO(n29181));
    SB_LUT4 add_5233_7_lut (.I0(GND_net), .I1(n9826[4]), .I2(n466_adj_4549), 
            .I3(n29179), .O(n9810[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_7 (.CI(n29179), .I0(n9826[4]), .I1(n466_adj_4549), 
            .CO(n29180));
    SB_LUT4 add_5233_6_lut (.I0(GND_net), .I1(n9826[3]), .I2(n393_adj_4550), 
            .I3(n29178), .O(n9810[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_6 (.CI(n29178), .I0(n9826[3]), .I1(n393_adj_4550), 
            .CO(n29179));
    SB_LUT4 add_5233_5_lut (.I0(GND_net), .I1(n9826[2]), .I2(n320), .I3(n29177), 
            .O(n9810[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_5 (.CI(n29177), .I0(n9826[2]), .I1(n320), .CO(n29178));
    SB_LUT4 add_5233_4_lut (.I0(GND_net), .I1(n9826[1]), .I2(n247), .I3(n29176), 
            .O(n9810[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_4 (.CI(n29176), .I0(n9826[1]), .I1(n247), .CO(n29177));
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n27777), .O(duty_23__N_3609[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5233_3_lut (.I0(GND_net), .I1(n9826[0]), .I2(n174), .I3(n29175), 
            .O(n9810[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_3 (.CI(n29175), .I0(n9826[0]), .I1(n174), .CO(n29176));
    SB_LUT4 add_5233_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n9810[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5233_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5233_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n29175));
    SB_LUT4 add_5232_16_lut (.I0(GND_net), .I1(n9810[13]), .I2(n1120), 
            .I3(n29174), .O(n9793[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5232_15_lut (.I0(GND_net), .I1(n9810[12]), .I2(n1047), 
            .I3(n29173), .O(n9793[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_15 (.CI(n29173), .I0(n9810[12]), .I1(n1047), .CO(n29174));
    SB_LUT4 i30033_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n38226), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4436), .O(n36430));
    defparam i30033_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_233_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n38195));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_233_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29631_2_lut_4_lut (.I0(duty_23__N_3609[21]), .I1(n257[21]), 
            .I2(duty_23__N_3609[9]), .I3(n257[9]), .O(n36027));
    defparam i29631_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5232_14_lut (.I0(GND_net), .I1(n9810[11]), .I2(n974), 
            .I3(n29172), .O(n9793[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_14 (.CI(n29172), .I0(n9810[11]), .I1(n974), .CO(n29173));
    SB_LUT4 i30021_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n38195), 
            .I2(IntegralLimit[14]), .I3(n36430), .O(n36418));
    defparam i30021_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5232_13_lut (.I0(GND_net), .I1(n9810[10]), .I2(n901), 
            .I3(n29171), .O(n9793[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29643_2_lut_4_lut (.I0(duty_23__N_3609[16]), .I1(n257[16]), 
            .I2(duty_23__N_3609[7]), .I3(n257[7]), .O(n36039));
    defparam i29643_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5232_13 (.CI(n29171), .I0(n9810[10]), .I1(n901), .CO(n29172));
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_227_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n38189));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_227_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5232_12_lut (.I0(GND_net), .I1(n9810[9]), .I2(n828), .I3(n29170), 
            .O(n9793[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_12 (.CI(n29170), .I0(n9810[9]), .I1(n828), .CO(n29171));
    SB_LUT4 i29669_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3609[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3609[9]), .O(n36065));
    defparam i29669_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5232_11_lut (.I0(GND_net), .I1(n9810[8]), .I2(n755), .I3(n29169), 
            .O(n9793[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_11 (.CI(n29169), .I0(n9810[8]), .I1(n755), .CO(n29170));
    SB_LUT4 add_5232_10_lut (.I0(GND_net), .I1(n9810[7]), .I2(n682), .I3(n29168), 
            .O(n9793[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_10 (.CI(n29168), .I0(n9810[7]), .I1(n682), .CO(n29169));
    SB_LUT4 add_5232_9_lut (.I0(GND_net), .I1(n9810[6]), .I2(n609), .I3(n29167), 
            .O(n9793[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_9 (.CI(n29167), .I0(n9810[6]), .I1(n609), .CO(n29168));
    SB_LUT4 add_5232_8_lut (.I0(GND_net), .I1(n9810[5]), .I2(n536), .I3(n29166), 
            .O(n9793[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_8 (.CI(n29166), .I0(n9810[5]), .I1(n536), .CO(n29167));
    SB_LUT4 add_5232_7_lut (.I0(GND_net), .I1(n9810[4]), .I2(n463), .I3(n29165), 
            .O(n9793[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_7 (.CI(n29165), .I0(n9810[4]), .I1(n463), .CO(n29166));
    SB_LUT4 add_5232_6_lut (.I0(GND_net), .I1(n9810[3]), .I2(n390), .I3(n29164), 
            .O(n9793[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4551));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29751_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n36147));
    defparam i29751_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_5232_6 (.CI(n29164), .I0(n9810[3]), .I1(n390), .CO(n29165));
    SB_LUT4 add_5232_5_lut (.I0(GND_net), .I1(n9810[2]), .I2(n317), .I3(n29163), 
            .O(n9793[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29679_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3609[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3609[7]), .O(n36075));
    defparam i29679_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5232_5 (.CI(n29163), .I0(n9810[2]), .I1(n317), .CO(n29164));
    SB_LUT4 add_5232_4_lut (.I0(GND_net), .I1(n9810[1]), .I2(n244), .I3(n29162), 
            .O(n9793[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_4 (.CI(n29162), .I0(n9810[1]), .I1(n244), .CO(n29163));
    SB_LUT4 add_5232_3_lut (.I0(GND_net), .I1(n9810[0]), .I2(n171), .I3(n29161), 
            .O(n9793[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5232_3 (.CI(n29161), .I0(n9810[0]), .I1(n171), .CO(n29162));
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_251_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n38213));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_251_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5232_2_lut (.I0(GND_net), .I1(n29_adj_4552), .I2(n98), 
            .I3(GND_net), .O(n9793[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5232_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4553));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5232_2 (.CI(GND_net), .I0(n29_adj_4552), .I1(n98), .CO(n29161));
    SB_LUT4 add_5231_17_lut (.I0(GND_net), .I1(n9793[14]), .I2(GND_net), 
            .I3(n29160), .O(n9775[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4551), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_4554));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5231_16_lut (.I0(GND_net), .I1(n9793[13]), .I2(n1117), 
            .I3(n29159), .O(n9775[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_16 (.CI(n29159), .I0(n9793[13]), .I1(n1117), .CO(n29160));
    SB_LUT4 add_5231_15_lut (.I0(GND_net), .I1(n9793[12]), .I2(n1044), 
            .I3(n29158), .O(n9775[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_15 (.CI(n29158), .I0(n9793[12]), .I1(n1044), .CO(n29159));
    SB_LUT4 i30179_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n38208), 
            .I2(IntegralLimit[11]), .I3(n36428), .O(n36576));
    defparam i30179_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_5231_14_lut (.I0(GND_net), .I1(n9793[11]), .I2(n971), 
            .I3(n29157), .O(n9775[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_14 (.CI(n29157), .I0(n9793[11]), .I1(n971), .CO(n29158));
    SB_LUT4 add_5231_13_lut (.I0(GND_net), .I1(n9793[10]), .I2(n898), 
            .I3(n29156), .O(n9775[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_13 (.CI(n29156), .I0(n9793[10]), .I1(n898), .CO(n29157));
    SB_LUT4 add_5231_12_lut (.I0(GND_net), .I1(n9793[9]), .I2(n825), .I3(n29155), 
            .O(n9775[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_12 (.CI(n29155), .I0(n9793[9]), .I1(n825), .CO(n29156));
    SB_LUT4 add_5231_11_lut (.I0(GND_net), .I1(n9793[8]), .I2(n752), .I3(n29154), 
            .O(n9775[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_11 (.CI(n29154), .I0(n9793[8]), .I1(n752), .CO(n29155));
    SB_LUT4 add_5231_10_lut (.I0(GND_net), .I1(n9793[7]), .I2(n679), .I3(n29153), 
            .O(n9775[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_10 (.CI(n29153), .I0(n9793[7]), .I1(n679), .CO(n29154));
    SB_LUT4 add_5231_9_lut (.I0(GND_net), .I1(n9793[6]), .I2(n606), .I3(n29152), 
            .O(n9775[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_23 (.CI(n27777), .I0(n106[21]), .I1(n155[21]), .CO(n27778));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1[2]), .I3(n27907), .O(n5_adj_4508)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29760_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n38201), 
            .I2(IntegralLimit[13]), .I3(n36576), .O(n36156));
    defparam i29760_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n27776), .O(duty_23__N_3609[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_9 (.CI(n29152), .I0(n9793[6]), .I1(n606), .CO(n29153));
    SB_LUT4 add_5231_8_lut (.I0(GND_net), .I1(n9793[5]), .I2(n533), .I3(n29151), 
            .O(n9775[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_8 (.CI(n29151), .I0(n9793[5]), .I1(n533), .CO(n29152));
    SB_LUT4 add_5231_7_lut (.I0(GND_net), .I1(n9793[4]), .I2(n460), .I3(n29150), 
            .O(n9775[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_231_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n38193));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_231_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30131_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n38193), 
            .I2(IntegralLimit[15]), .I3(n36156), .O(n36528));
    defparam i30131_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_257_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n38219));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_257_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i30274_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n38219), 
            .I2(IntegralLimit[17]), .I3(n36528), .O(n36671));
    defparam i30274_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_5231_7 (.CI(n29150), .I0(n9793[4]), .I1(n460), .CO(n29151));
    SB_LUT4 add_5231_6_lut (.I0(GND_net), .I1(n9793[3]), .I2(n387), .I3(n29149), 
            .O(n9775[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n27907), .I0(GND_net), .I1(n1[2]), 
            .CO(n27908));
    SB_CARRY add_5231_6 (.CI(n29149), .I0(n9793[3]), .I1(n387), .CO(n29150));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1[1]), .I3(n27906), .O(n3_adj_4557)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_222_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n38184));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_222_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n27906), .I0(GND_net), .I1(n1[1]), 
            .CO(n27907));
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5231_5_lut (.I0(GND_net), .I1(n9793[2]), .I2(n314), .I3(n29148), 
            .O(n9775[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_5 (.CI(n29148), .I0(n9793[2]), .I1(n314), .CO(n29149));
    SB_LUT4 add_5231_4_lut (.I0(GND_net), .I1(n9793[1]), .I2(n241), .I3(n29147), 
            .O(n9775[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_4 (.CI(n29147), .I0(n9793[1]), .I1(n241), .CO(n29148));
    SB_LUT4 add_5231_3_lut (.I0(GND_net), .I1(n9793[0]), .I2(n168), .I3(n29146), 
            .O(n9775[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5231_3 (.CI(n29146), .I0(n9793[0]), .I1(n168), .CO(n29147));
    SB_LUT4 i30346_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n38184), 
            .I2(IntegralLimit[19]), .I3(n36671), .O(n36743));
    defparam i30346_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 add_5231_2_lut (.I0(GND_net), .I1(n26_adj_4561), .I2(n95), 
            .I3(GND_net), .O(n9775[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5231_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5231_2 (.CI(GND_net), .I0(n26_adj_4561), .I1(n95), .CO(n29146));
    SB_LUT4 add_5230_18_lut (.I0(GND_net), .I1(n9775[15]), .I2(GND_net), 
            .I3(n29145), .O(n9756[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5230_17_lut (.I0(GND_net), .I1(n9775[14]), .I2(GND_net), 
            .I3(n29144), .O(n9756[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_17 (.CI(n29144), .I0(n9775[14]), .I1(GND_net), .CO(n29145));
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_219_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n38181));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_219_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4562));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5230_16_lut (.I0(GND_net), .I1(n9775[13]), .I2(n1114), 
            .I3(n29143), .O(n9756[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n27776), .I0(n106[20]), .I1(n155[20]), .CO(n27777));
    SB_CARRY add_5230_16 (.CI(n29143), .I0(n9775[13]), .I1(n1114), .CO(n29144));
    SB_LUT4 add_5230_15_lut (.I0(GND_net), .I1(n9775[12]), .I2(n1041), 
            .I3(n29142), .O(n9756[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29740_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n36136));
    defparam i29740_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_5230_15 (.CI(n29142), .I0(n9775[12]), .I1(n1041), .CO(n29143));
    SB_LUT4 add_5230_14_lut (.I0(GND_net), .I1(n9775[11]), .I2(n968), 
            .I3(n29141), .O(n9756[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_14 (.CI(n29141), .I0(n9775[11]), .I1(n968), .CO(n29142));
    SB_LUT4 add_5230_13_lut (.I0(GND_net), .I1(n9775[10]), .I2(n895), 
            .I3(n29140), .O(n9756[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_13 (.CI(n29140), .I0(n9775[10]), .I1(n895), .CO(n29141));
    SB_LUT4 add_5230_12_lut (.I0(GND_net), .I1(n9775[9]), .I2(n822), .I3(n29139), 
            .O(n9756[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5230_12 (.CI(n29139), .I0(n9775[9]), .I1(n822), .CO(n29140));
    SB_LUT4 add_5230_11_lut (.I0(GND_net), .I1(n9775[8]), .I2(n749), .I3(n29138), 
            .O(n9756[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_11 (.CI(n29138), .I0(n9775[8]), .I1(n749), .CO(n29139));
    SB_LUT4 add_5230_10_lut (.I0(GND_net), .I1(n9775[7]), .I2(n676), .I3(n29137), 
            .O(n9756[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_10 (.CI(n29137), .I0(n9775[7]), .I1(n676), .CO(n29138));
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4562), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4563));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5230_9_lut (.I0(GND_net), .I1(n9775[6]), .I2(n603), .I3(n29136), 
            .O(n9756[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_9 (.CI(n29136), .I0(n9775[6]), .I1(n603), .CO(n29137));
    SB_LUT4 add_5230_8_lut (.I0(GND_net), .I1(n9775[5]), .I2(n530), .I3(n29135), 
            .O(n9756[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_8 (.CI(n29135), .I0(n9775[5]), .I1(n530), .CO(n29136));
    SB_LUT4 add_5230_7_lut (.I0(GND_net), .I1(n9775[4]), .I2(n457), .I3(n29134), 
            .O(n9756[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4564));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5230_7 (.CI(n29134), .I0(n9775[4]), .I1(n457), .CO(n29135));
    SB_LUT4 add_5230_6_lut (.I0(GND_net), .I1(n9775[3]), .I2(n384), .I3(n29133), 
            .O(n9756[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_6 (.CI(n29133), .I0(n9775[3]), .I1(n384), .CO(n29134));
    SB_LUT4 add_5230_5_lut (.I0(GND_net), .I1(n9775[2]), .I2(n311), .I3(n29132), 
            .O(n9756[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30278_3_lut (.I0(n6_adj_4564), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n36675));   // verilog/motorControl.v(31[10:34])
    defparam i30278_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5230_5 (.CI(n29132), .I0(n9775[2]), .I1(n311), .CO(n29133));
    SB_LUT4 add_5230_4_lut (.I0(GND_net), .I1(n9775[1]), .I2(n238), .I3(n29131), 
            .O(n9756[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_4 (.CI(n29131), .I0(n9775[1]), .I1(n238), .CO(n29132));
    SB_LUT4 add_5230_3_lut (.I0(GND_net), .I1(n9775[0]), .I2(n165), .I3(n29130), 
            .O(n9756[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_3 (.CI(n29130), .I0(n9775[0]), .I1(n165), .CO(n29131));
    SB_LUT4 add_5230_2_lut (.I0(GND_net), .I1(n23_adj_4565), .I2(n92), 
            .I3(GND_net), .O(n9756[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5230_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5230_2 (.CI(GND_net), .I0(n23_adj_4565), .I1(n92), .CO(n29130));
    SB_LUT4 add_5229_19_lut (.I0(GND_net), .I1(n9756[16]), .I2(GND_net), 
            .I3(n29129), .O(n9736[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5229_18_lut (.I0(GND_net), .I1(n9756[15]), .I2(GND_net), 
            .I3(n29128), .O(n9736[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_18 (.CI(n29128), .I0(n9756[15]), .I1(GND_net), .CO(n29129));
    SB_LUT4 add_5229_17_lut (.I0(GND_net), .I1(n9756[14]), .I2(GND_net), 
            .I3(n29127), .O(n9736[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_17 (.CI(n29127), .I0(n9756[14]), .I1(GND_net), .CO(n29128));
    SB_LUT4 add_5229_16_lut (.I0(GND_net), .I1(n9756[13]), .I2(n1111), 
            .I3(n29126), .O(n9736[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_16 (.CI(n29126), .I0(n9756[13]), .I1(n1111), .CO(n29127));
    SB_LUT4 add_5229_15_lut (.I0(GND_net), .I1(n9756[12]), .I2(n1038), 
            .I3(n29125), .O(n9736[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30279_3_lut (.I0(n36675), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n36676));   // verilog/motorControl.v(31[10:34])
    defparam i30279_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29742_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n38201), 
            .I2(IntegralLimit[21]), .I3(n36424), .O(n36138));
    defparam i29742_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i30139_4_lut (.I0(n24_adj_4563), .I1(n8_adj_4532), .I2(n38179), 
            .I3(n36136), .O(n36536));   // verilog/motorControl.v(31[10:34])
    defparam i30139_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5229_15 (.CI(n29125), .I0(n9756[12]), .I1(n1038), .CO(n29126));
    SB_LUT4 add_5229_14_lut (.I0(GND_net), .I1(n9756[11]), .I2(n965), 
            .I3(n29124), .O(n9736[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_14 (.CI(n29124), .I0(n9756[11]), .I1(n965), .CO(n29125));
    SB_LUT4 add_5229_13_lut (.I0(GND_net), .I1(n9756[10]), .I2(n892), 
            .I3(n29123), .O(n9736[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30182_3_lut (.I0(n36676), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n36579));   // verilog/motorControl.v(31[10:34])
    defparam i30182_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3560 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4557), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4566));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30246_3_lut (.I0(n4_adj_4566), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n36643));   // verilog/motorControl.v(31[38:63])
    defparam i30246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22794_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3509 [19]), 
            .O(n9925[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22794_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30247_3_lut (.I0(n36643), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n36644));   // verilog/motorControl.v(31[38:63])
    defparam i30247_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5229_13 (.CI(n29123), .I0(n9756[10]), .I1(n892), .CO(n29124));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4567));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_5229_12_lut (.I0(GND_net), .I1(n9756[9]), .I2(n819), .I3(n29122), 
            .O(n9736[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29715_2_lut (.I0(n33), .I1(n15_adj_4439), .I2(GND_net), .I3(GND_net), 
            .O(n36111));
    defparam i29715_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_5229_12 (.CI(n29122), .I0(n9756[9]), .I1(n819), .CO(n29123));
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5229_11_lut (.I0(GND_net), .I1(n9756[8]), .I2(n746), .I3(n29121), 
            .O(n9736[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4440), .I3(GND_net), 
            .O(n10_adj_4568));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3560 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4567), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4402), .I3(GND_net), 
            .O(n30_adj_4570));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29717_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n36117), 
            .O(n36113));
    defparam i29717_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746_adj_4571));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n27906));
    SB_CARRY add_5229_11 (.CI(n29121), .I0(n9756[8]), .I1(n746), .CO(n29122));
    SB_LUT4 add_5229_10_lut (.I0(GND_net), .I1(n9756[7]), .I2(n673_adj_4572), 
            .I3(n29120), .O(n9736[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819_adj_4573));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5229_10 (.CI(n29120), .I0(n9756[7]), .I1(n673_adj_4572), 
            .CO(n29121));
    SB_LUT4 add_5229_9_lut (.I0(GND_net), .I1(n9756[6]), .I2(n600_adj_4574), 
            .I3(n29119), .O(n9736[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_9 (.CI(n29119), .I0(n9756[6]), .I1(n600_adj_4574), 
            .CO(n29120));
    SB_LUT4 add_5229_8_lut (.I0(GND_net), .I1(n9756[5]), .I2(n527_adj_4575), 
            .I3(n29118), .O(n9736[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_8 (.CI(n29118), .I0(n9756[5]), .I1(n527_adj_4575), 
            .CO(n29119));
    SB_LUT4 add_5229_7_lut (.I0(GND_net), .I1(n9756[4]), .I2(n454_adj_4576), 
            .I3(n29117), .O(n9736[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892_adj_4577));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5229_7 (.CI(n29117), .I0(n9756[4]), .I1(n454_adj_4576), 
            .CO(n29118));
    SB_LUT4 add_5229_6_lut (.I0(GND_net), .I1(n9756[3]), .I2(n381_adj_4578), 
            .I3(n29116), .O(n9736[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_6 (.CI(n29116), .I0(n9756[3]), .I1(n381_adj_4578), 
            .CO(n29117));
    SB_LUT4 add_5229_5_lut (.I0(GND_net), .I1(n9756[2]), .I2(n308_adj_4579), 
            .I3(n29115), .O(n9736[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_5 (.CI(n29115), .I0(n9756[2]), .I1(n308_adj_4579), 
            .CO(n29116));
    SB_LUT4 add_5229_4_lut (.I0(GND_net), .I1(n9756[1]), .I2(n235_adj_4580), 
            .I3(n29114), .O(n9736[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_4 (.CI(n29114), .I0(n9756[1]), .I1(n235_adj_4580), 
            .CO(n29115));
    SB_LUT4 add_5229_3_lut (.I0(GND_net), .I1(n9756[0]), .I2(n162_adj_4581), 
            .I3(n29113), .O(n9736[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_3 (.CI(n29113), .I0(n9756[0]), .I1(n162_adj_4581), 
            .CO(n29114));
    SB_LUT4 add_5229_2_lut (.I0(GND_net), .I1(n20_adj_4582), .I2(n89_adj_4583), 
            .I3(GND_net), .O(n9736[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5229_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5229_2 (.CI(GND_net), .I0(n20_adj_4582), .I1(n89_adj_4583), 
            .CO(n29113));
    SB_LUT4 add_5228_20_lut (.I0(GND_net), .I1(n9736[17]), .I2(GND_net), 
            .I3(n29112), .O(n9715[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5228_19_lut (.I0(GND_net), .I1(n9736[16]), .I2(GND_net), 
            .I3(n29111), .O(n9715[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_19 (.CI(n29111), .I0(n9736[16]), .I1(GND_net), .CO(n29112));
    SB_LUT4 add_5228_18_lut (.I0(GND_net), .I1(n9736[15]), .I2(GND_net), 
            .I3(n29110), .O(n9715[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_18 (.CI(n29110), .I0(n9736[15]), .I1(GND_net), .CO(n29111));
    SB_LUT4 add_5228_17_lut (.I0(GND_net), .I1(n9736[14]), .I2(GND_net), 
            .I3(n29109), .O(n9715[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_17 (.CI(n29109), .I0(n9736[14]), .I1(GND_net), .CO(n29110));
    SB_LUT4 add_5228_16_lut (.I0(GND_net), .I1(n9736[13]), .I2(n1108_adj_4584), 
            .I3(n29108), .O(n9715[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_16 (.CI(n29108), .I0(n9736[13]), .I1(n1108_adj_4584), 
            .CO(n29109));
    SB_LUT4 add_5228_15_lut (.I0(GND_net), .I1(n9736[12]), .I2(n1035_adj_4585), 
            .I3(n29107), .O(n9715[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_15 (.CI(n29107), .I0(n9736[12]), .I1(n1035_adj_4585), 
            .CO(n29108));
    SB_LUT4 add_5228_14_lut (.I0(GND_net), .I1(n9736[11]), .I2(n962_adj_4586), 
            .I3(n29106), .O(n9715[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_14 (.CI(n29106), .I0(n9736[11]), .I1(n962_adj_4586), 
            .CO(n29107));
    SB_LUT4 add_5228_13_lut (.I0(GND_net), .I1(n9736[10]), .I2(n889_adj_4587), 
            .I3(n29105), .O(n9715[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_13 (.CI(n29105), .I0(n9736[10]), .I1(n889_adj_4587), 
            .CO(n29106));
    SB_LUT4 add_5228_12_lut (.I0(GND_net), .I1(n9736[9]), .I2(n816_adj_4588), 
            .I3(n29104), .O(n9715[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_12 (.CI(n29104), .I0(n9736[9]), .I1(n816_adj_4588), 
            .CO(n29105));
    SB_LUT4 add_5228_11_lut (.I0(GND_net), .I1(n9736[8]), .I2(n743_adj_4589), 
            .I3(n29103), .O(n9715[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30330_4_lut (.I0(n30_adj_4570), .I1(n10_adj_4568), .I2(n35_adj_4402), 
            .I3(n36111), .O(n36727));   // verilog/motorControl.v(31[38:63])
    defparam i30330_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5228_11 (.CI(n29103), .I0(n9736[8]), .I1(n743_adj_4589), 
            .CO(n29104));
    SB_LUT4 add_5228_10_lut (.I0(GND_net), .I1(n9736[7]), .I2(n670_adj_4590), 
            .I3(n29102), .O(n9715[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_10 (.CI(n29102), .I0(n9736[7]), .I1(n670_adj_4590), 
            .CO(n29103));
    SB_LUT4 add_5228_9_lut (.I0(GND_net), .I1(n9736[6]), .I2(n597_adj_4591), 
            .I3(n29101), .O(n9715[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_9 (.CI(n29101), .I0(n9736[6]), .I1(n597_adj_4591), 
            .CO(n29102));
    SB_LUT4 add_5228_8_lut (.I0(GND_net), .I1(n9736[5]), .I2(n524_adj_4592), 
            .I3(n29100), .O(n9715[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30190_3_lut (.I0(n36644), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n36587));   // verilog/motorControl.v(31[38:63])
    defparam i30190_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5228_8 (.CI(n29100), .I0(n9736[5]), .I1(n524_adj_4592), 
            .CO(n29101));
    SB_LUT4 add_5228_7_lut (.I0(GND_net), .I1(n9736[4]), .I2(n451_adj_4593), 
            .I3(n29099), .O(n9715[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_7 (.CI(n29099), .I0(n9736[4]), .I1(n451_adj_4593), 
            .CO(n29100));
    SB_LUT4 add_5228_6_lut (.I0(GND_net), .I1(n9736[3]), .I2(n378_adj_4594), 
            .I3(n29098), .O(n9715[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_6 (.CI(n29098), .I0(n9736[3]), .I1(n378_adj_4594), 
            .CO(n29099));
    SB_LUT4 add_5228_5_lut (.I0(GND_net), .I1(n9736[2]), .I2(n305_adj_4595), 
            .I3(n29097), .O(n9715[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_5 (.CI(n29097), .I0(n9736[2]), .I1(n305_adj_4595), 
            .CO(n29098));
    SB_LUT4 add_5228_4_lut (.I0(GND_net), .I1(n9736[1]), .I2(n232_adj_4596), 
            .I3(n29096), .O(n9715[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_4 (.CI(n29096), .I0(n9736[1]), .I1(n232_adj_4596), 
            .CO(n29097));
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965_adj_4597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30381_4_lut (.I0(n36587), .I1(n36727), .I2(n35_adj_4402), 
            .I3(n36113), .O(n36778));   // verilog/motorControl.v(31[38:63])
    defparam i30381_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30382_3_lut (.I0(n36778), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n36779));   // verilog/motorControl.v(31[38:63])
    defparam i30382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30365_3_lut (.I0(n36779), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n36762));   // verilog/motorControl.v(31[38:63])
    defparam i30365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4507), .I3(GND_net), 
            .O(n6_adj_4598));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_5228_3_lut (.I0(GND_net), .I1(n9736[0]), .I2(n159_adj_4599), 
            .I3(n29095), .O(n9715[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038_adj_4600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5228_3 (.CI(n29095), .I0(n9736[0]), .I1(n159_adj_4599), 
            .CO(n29096));
    SB_LUT4 add_5228_2_lut (.I0(GND_net), .I1(n17_adj_4601), .I2(n86_adj_4602), 
            .I3(GND_net), .O(n9715[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5228_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5228_2 (.CI(GND_net), .I0(n17_adj_4601), .I1(n86_adj_4602), 
            .CO(n29095));
    SB_LUT4 add_5227_21_lut (.I0(GND_net), .I1(n9715[18]), .I2(GND_net), 
            .I3(n29094), .O(n9693[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5227_20_lut (.I0(GND_net), .I1(n9715[17]), .I2(GND_net), 
            .I3(n29093), .O(n9693[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_20 (.CI(n29093), .I0(n9715[17]), .I1(GND_net), .CO(n29094));
    SB_LUT4 add_5227_19_lut (.I0(GND_net), .I1(n9715[16]), .I2(GND_net), 
            .I3(n29092), .O(n9693[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_19 (.CI(n29092), .I0(n9715[16]), .I1(GND_net), .CO(n29093));
    SB_LUT4 add_5227_18_lut (.I0(GND_net), .I1(n9715[15]), .I2(GND_net), 
            .I3(n29091), .O(n9693[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_18 (.CI(n29091), .I0(n9715[15]), .I1(GND_net), .CO(n29092));
    SB_LUT4 add_5227_17_lut (.I0(GND_net), .I1(n9715[14]), .I2(GND_net), 
            .I3(n29090), .O(n9693[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30254_3_lut (.I0(n6_adj_4598), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4442), .I3(GND_net), .O(n36651));   // verilog/motorControl.v(31[38:63])
    defparam i30254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30255_3_lut (.I0(n36651), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4509), .I3(GND_net), .O(n36652));   // verilog/motorControl.v(31[38:63])
    defparam i30255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29707_4_lut (.I0(n43), .I1(n25_adj_4486), .I2(n23_adj_4509), 
            .I3(n36123), .O(n36103));
    defparam i29707_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30141_4_lut (.I0(n24_adj_4503), .I1(n8_adj_4474), .I2(n45), 
            .I3(n36101), .O(n36538));   // verilog/motorControl.v(31[38:63])
    defparam i30141_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30188_3_lut (.I0(n36652), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4486), .I3(GND_net), .O(n36585));   // verilog/motorControl.v(31[38:63])
    defparam i30188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111_adj_4603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29709_4_lut (.I0(n43), .I1(n41_adj_4395), .I2(n39), .I3(n36721), 
            .O(n36105));
    defparam i29709_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30288_4_lut (.I0(n36585), .I1(n36538), .I2(n45), .I3(n36103), 
            .O(n36685));   // verilog/motorControl.v(31[38:63])
    defparam i30288_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5227_17 (.CI(n29090), .I0(n9715[14]), .I1(GND_net), .CO(n29091));
    SB_LUT4 add_5227_16_lut (.I0(GND_net), .I1(n9715[13]), .I2(n1105_adj_4604), 
            .I3(n29089), .O(n9693[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_16 (.CI(n29089), .I0(n9715[13]), .I1(n1105_adj_4604), 
            .CO(n29090));
    SB_LUT4 add_5227_15_lut (.I0(GND_net), .I1(n9715[12]), .I2(n1032_adj_4605), 
            .I3(n29088), .O(n9693[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_15 (.CI(n29088), .I0(n9715[12]), .I1(n1032_adj_4605), 
            .CO(n29089));
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n27775), .O(duty_23__N_3609[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30351_3_lut (.I0(n36762), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4395), .I3(GND_net), .O(n40_adj_4606));   // verilog/motorControl.v(31[38:63])
    defparam i30351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30290_4_lut (.I0(n40_adj_4606), .I1(n36685), .I2(n45), .I3(n36105), 
            .O(n36687));   // verilog/motorControl.v(31[38:63])
    defparam i30290_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5227_14_lut (.I0(GND_net), .I1(n9715[11]), .I2(n959_adj_4607), 
            .I3(n29087), .O(n9693[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_14 (.CI(n29087), .I0(n9715[11]), .I1(n959_adj_4607), 
            .CO(n29088));
    SB_CARRY add_12_21 (.CI(n27775), .I0(n106[19]), .I1(n155[19]), .CO(n27776));
    SB_LUT4 add_5227_13_lut (.I0(GND_net), .I1(n9715[10]), .I2(n886_adj_4608), 
            .I3(n29086), .O(n9693[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_13 (.CI(n29086), .I0(n9715[10]), .I1(n886_adj_4608), 
            .CO(n29087));
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4609));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 add_5227_12_lut (.I0(GND_net), .I1(n9715[9]), .I2(n813_adj_4610), 
            .I3(n29085), .O(n9693[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30270_3_lut (.I0(n4_adj_4609), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n36667));   // verilog/motorControl.v(31[10:34])
    defparam i30270_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5227_12 (.CI(n29085), .I0(n9715[9]), .I1(n813_adj_4610), 
            .CO(n29086));
    SB_LUT4 i30271_3_lut (.I0(n36667), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n36668));   // verilog/motorControl.v(31[10:34])
    defparam i30271_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29753_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n38189), 
            .I2(IntegralLimit[16]), .I3(n36418), .O(n36149));
    defparam i29753_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i30328_4_lut (.I0(n30_adj_4554), .I1(n10_adj_4553), .I2(n38213), 
            .I3(n36147), .O(n36725));   // verilog/motorControl.v(31[10:34])
    defparam i30328_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_5227_11_lut (.I0(GND_net), .I1(n9715[8]), .I2(n740_adj_4611), 
            .I3(n29084), .O(n9693[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n27774), .O(duty_23__N_3609[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30184_3_lut (.I0(n36668), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n36581));   // verilog/motorControl.v(31[10:34])
    defparam i30184_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5227_11 (.CI(n29084), .I0(n9715[8]), .I1(n740_adj_4611), 
            .CO(n29085));
    SB_LUT4 add_5227_10_lut (.I0(GND_net), .I1(n9715[7]), .I2(n667_adj_4612), 
            .I3(n29083), .O(n9693[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_20 (.CI(n27774), .I0(n106[18]), .I1(n155[18]), .CO(n27775));
    SB_LUT4 i30379_4_lut (.I0(n36581), .I1(n36725), .I2(n38213), .I3(n36149), 
            .O(n36776));   // verilog/motorControl.v(31[10:34])
    defparam i30379_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30380_3_lut (.I0(n36776), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n36777));   // verilog/motorControl.v(31[10:34])
    defparam i30380_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5227_10 (.CI(n29083), .I0(n9715[7]), .I1(n667_adj_4612), 
            .CO(n29084));
    SB_LUT4 i30367_3_lut (.I0(n36777), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n36764));   // verilog/motorControl.v(31[10:34])
    defparam i30367_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n27773), .O(duty_23__N_3609[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5227_9_lut (.I0(GND_net), .I1(n9715[6]), .I2(n594_adj_4614), 
            .I3(n29082), .O(n9693[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_9 (.CI(n29082), .I0(n9715[6]), .I1(n594_adj_4614), 
            .CO(n29083));
    SB_LUT4 add_5227_8_lut (.I0(GND_net), .I1(n9715[5]), .I2(n521_adj_4615), 
            .I3(n29081), .O(n9693[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n27773), .I0(n106[17]), .I1(n155[17]), .CO(n27774));
    SB_CARRY add_5227_8 (.CI(n29081), .I0(n9715[5]), .I1(n521_adj_4615), 
            .CO(n29082));
    SB_LUT4 add_5227_7_lut (.I0(GND_net), .I1(n9715[4]), .I2(n448_adj_4616), 
            .I3(n29080), .O(n9693[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_7 (.CI(n29080), .I0(n9715[4]), .I1(n448_adj_4616), 
            .CO(n29081));
    SB_LUT4 add_5227_6_lut (.I0(GND_net), .I1(n9715[3]), .I2(n375_adj_4617), 
            .I3(n29079), .O(n9693[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_6 (.CI(n29079), .I0(n9715[3]), .I1(n375_adj_4617), 
            .CO(n29080));
    SB_LUT4 add_5227_5_lut (.I0(GND_net), .I1(n9715[2]), .I2(n302_adj_4618), 
            .I3(n29078), .O(n9693[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_5 (.CI(n29078), .I0(n9715[2]), .I1(n302_adj_4618), 
            .CO(n29079));
    SB_LUT4 add_5227_4_lut (.I0(GND_net), .I1(n9715[1]), .I2(n229_adj_4619), 
            .I3(n29077), .O(n9693[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_4 (.CI(n29077), .I0(n9715[1]), .I1(n229_adj_4619), 
            .CO(n29078));
    SB_LUT4 add_5227_3_lut (.I0(GND_net), .I1(n9715[0]), .I2(n156_adj_4620), 
            .I3(n29076), .O(n9693[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_3 (.CI(n29076), .I0(n9715[0]), .I1(n156_adj_4620), 
            .CO(n29077));
    SB_LUT4 add_5227_2_lut (.I0(GND_net), .I1(n14_adj_4621), .I2(n83_adj_4622), 
            .I3(GND_net), .O(n9693[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5227_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5227_2 (.CI(GND_net), .I0(n14_adj_4621), .I1(n83_adj_4622), 
            .CO(n29076));
    SB_LUT4 add_5226_22_lut (.I0(GND_net), .I1(n9693[19]), .I2(GND_net), 
            .I3(n29075), .O(n9670[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5226_21_lut (.I0(GND_net), .I1(n9693[18]), .I2(GND_net), 
            .I3(n29074), .O(n9670[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_21 (.CI(n29074), .I0(n9693[18]), .I1(GND_net), .CO(n29075));
    SB_LUT4 add_5226_20_lut (.I0(GND_net), .I1(n9693[17]), .I2(GND_net), 
            .I3(n29073), .O(n9670[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_20 (.CI(n29073), .I0(n9693[17]), .I1(GND_net), .CO(n29074));
    SB_LUT4 add_5226_19_lut (.I0(GND_net), .I1(n9693[16]), .I2(GND_net), 
            .I3(n29072), .O(n9670[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_19 (.CI(n29072), .I0(n9693[16]), .I1(GND_net), .CO(n29073));
    SB_LUT4 add_5226_18_lut (.I0(GND_net), .I1(n9693[15]), .I2(GND_net), 
            .I3(n29071), .O(n9670[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_18 (.CI(n29071), .I0(n9693[15]), .I1(GND_net), .CO(n29072));
    SB_LUT4 add_5226_17_lut (.I0(GND_net), .I1(n9693[14]), .I2(GND_net), 
            .I3(n29070), .O(n9670[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_17 (.CI(n29070), .I0(n9693[14]), .I1(GND_net), .CO(n29071));
    SB_LUT4 add_5226_16_lut (.I0(GND_net), .I1(n9693[13]), .I2(n1102_adj_4623), 
            .I3(n29069), .O(n9670[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_16 (.CI(n29069), .I0(n9693[13]), .I1(n1102_adj_4623), 
            .CO(n29070));
    SB_LUT4 add_5226_15_lut (.I0(GND_net), .I1(n9693[12]), .I2(n1029_adj_4624), 
            .I3(n29068), .O(n9670[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_15 (.CI(n29068), .I0(n9693[12]), .I1(n1029_adj_4624), 
            .CO(n29069));
    SB_LUT4 add_5226_14_lut (.I0(GND_net), .I1(n9693[11]), .I2(n956_adj_4625), 
            .I3(n29067), .O(n9670[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_14 (.CI(n29067), .I0(n9693[11]), .I1(n956_adj_4625), 
            .CO(n29068));
    SB_LUT4 add_5226_13_lut (.I0(GND_net), .I1(n9693[10]), .I2(n883_adj_4626), 
            .I3(n29066), .O(n9670[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n27900), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_13 (.CI(n29066), .I0(n9693[10]), .I1(n883_adj_4626), 
            .CO(n29067));
    SB_LUT4 add_5226_12_lut (.I0(GND_net), .I1(n9693[9]), .I2(n810_adj_4627), 
            .I3(n29065), .O(n9670[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_12 (.CI(n29065), .I0(n9693[9]), .I1(n810_adj_4627), 
            .CO(n29066));
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n27772), .O(duty_23__N_3609[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5226_11_lut (.I0(GND_net), .I1(n9693[8]), .I2(n737_adj_4628), 
            .I3(n29064), .O(n9670[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_11 (.CI(n29064), .I0(n9693[8]), .I1(n737_adj_4628), 
            .CO(n29065));
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n27899), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5226_10_lut (.I0(GND_net), .I1(n9693[7]), .I2(n664_adj_4629), 
            .I3(n29063), .O(n9670[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_10 (.CI(n29063), .I0(n9693[7]), .I1(n664_adj_4629), 
            .CO(n29064));
    SB_LUT4 add_5226_9_lut (.I0(GND_net), .I1(n9693[6]), .I2(n591_adj_4630), 
            .I3(n29062), .O(n9670[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_9 (.CI(n29062), .I0(n9693[6]), .I1(n591_adj_4630), 
            .CO(n29063));
    SB_LUT4 add_5226_8_lut (.I0(GND_net), .I1(n9693[5]), .I2(n518_adj_4631), 
            .I3(n29061), .O(n9670[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_8 (.CI(n29061), .I0(n9693[5]), .I1(n518_adj_4631), 
            .CO(n29062));
    SB_LUT4 add_5226_7_lut (.I0(GND_net), .I1(n9693[4]), .I2(n445_adj_4632), 
            .I3(n29060), .O(n9670[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_7 (.CI(n29060), .I0(n9693[4]), .I1(n445_adj_4632), 
            .CO(n29061));
    SB_LUT4 add_5226_6_lut (.I0(GND_net), .I1(n9693[3]), .I2(n372_adj_4633), 
            .I3(n29059), .O(n9670[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_6 (.CI(n29059), .I0(n9693[3]), .I1(n372_adj_4633), 
            .CO(n29060));
    SB_LUT4 add_5226_5_lut (.I0(GND_net), .I1(n9693[2]), .I2(n299_adj_4634), 
            .I3(n29058), .O(n9670[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_5 (.CI(n29058), .I0(n9693[2]), .I1(n299_adj_4634), 
            .CO(n29059));
    SB_LUT4 add_5226_4_lut (.I0(GND_net), .I1(n9693[1]), .I2(n226_adj_4635), 
            .I3(n29057), .O(n9670[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_4 (.CI(n29057), .I0(n9693[1]), .I1(n226_adj_4635), 
            .CO(n29058));
    SB_LUT4 add_5226_3_lut (.I0(GND_net), .I1(n9693[0]), .I2(n153_adj_4636), 
            .I3(n29056), .O(n9670[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_3 (.CI(n29056), .I0(n9693[0]), .I1(n153_adj_4636), 
            .CO(n29057));
    SB_LUT4 add_5226_2_lut (.I0(GND_net), .I1(n11_adj_4637), .I2(n80_adj_4638), 
            .I3(GND_net), .O(n9670[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5226_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n27899), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n27900));
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n27898), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5226_2 (.CI(GND_net), .I0(n11_adj_4637), .I1(n80_adj_4638), 
            .CO(n29056));
    SB_LUT4 i29744_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n38181), 
            .I2(IntegralLimit[21]), .I3(n36743), .O(n36140));
    defparam i29744_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3509 [23]), 
            .I1(n9646[21]), .I2(GND_net), .I3(n29055), .O(n8064[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_217_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n38179));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_217_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n9646[20]), .I2(GND_net), 
            .I3(n29054), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n29054), .I0(n9646[20]), .I1(GND_net), 
            .CO(n29055));
    SB_LUT4 i30282_4_lut (.I0(n36579), .I1(n36536), .I2(n38179), .I3(n36138), 
            .O(n36679));   // verilog/motorControl.v(31[10:34])
    defparam i30282_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n9646[19]), .I2(GND_net), 
            .I3(n29053), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30349_3_lut (.I0(n36764), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n40_adj_4639));   // verilog/motorControl.v(31[10:34])
    defparam i30349_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30291_3_lut (.I0(n36687), .I1(\PID_CONTROLLER.integral_23__N_3560 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3559 ));   // verilog/motorControl.v(31[38:63])
    defparam i30291_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY mult_11_add_1225_22 (.CI(n29053), .I0(n9646[19]), .I1(GND_net), 
            .CO(n29054));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n9646[18]), .I2(GND_net), 
            .I3(n29052), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_23 (.CI(n27898), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n27899));
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n27897), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n29052), .I0(n9646[18]), .I1(GND_net), 
            .CO(n29053));
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4640));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30284_4_lut (.I0(n40_adj_4639), .I1(n36679), .I2(n38179), 
            .I3(n36140), .O(n36681));   // verilog/motorControl.v(31[10:34])
    defparam i30284_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n9646[17]), .I2(GND_net), 
            .I3(n29051), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4642));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_20 (.CI(n29051), .I0(n9646[17]), .I1(GND_net), 
            .CO(n29052));
    SB_CARRY add_12_18 (.CI(n27772), .I0(n106[16]), .I1(n155[16]), .CO(n27773));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n9646[16]), .I2(GND_net), 
            .I3(n29050), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_830_4_lut  (.I0(n36681), .I1(\PID_CONTROLLER.integral_23__N_3559 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3557 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_830_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n27771), .O(duty_23__N_3609[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n29050), .I0(n9646[16]), .I1(GND_net), 
            .CO(n29051));
    SB_CARRY add_12_17 (.CI(n27771), .I0(n106[15]), .I1(n155[15]), .CO(n27772));
    SB_CARRY sub_3_add_2_22 (.CI(n27897), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n27898));
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n27896), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n27896), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n27897));
    SB_LUT4 add_739_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n3223[23]), .I3(n27822), .O(\PID_CONTROLLER.integral_23__N_3509 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n3223[22]), .I3(n27821), .O(\PID_CONTROLLER.integral_23__N_3509 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n27895), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n27895), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n27896));
    SB_CARRY add_739_24 (.CI(n27821), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n3223[22]), .CO(n27822));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n27894), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4643));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n27770), .O(duty_23__N_3609[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n27894), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n27895));
    SB_LUT4 add_739_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n3223[21]), .I3(n27820), .O(\PID_CONTROLLER.integral_23__N_3509 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_16 (.CI(n27770), .I0(n106[14]), .I1(n155[14]), .CO(n27771));
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n27893), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n27893), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n27894));
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n27892), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n9646[15]), .I2(GND_net), 
            .I3(n29049), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_23 (.CI(n27820), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n3223[21]), .CO(n27821));
    SB_CARRY mult_11_add_1225_18 (.CI(n29049), .I0(n9646[15]), .I1(GND_net), 
            .CO(n29050));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n9646[14]), .I2(GND_net), 
            .I3(n29048), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n29048), .I0(n9646[14]), .I1(GND_net), 
            .CO(n29049));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n9646[13]), .I2(n1096_adj_4430), 
            .I3(n29047), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n29047), .I0(n9646[13]), .I1(n1096_adj_4430), 
            .CO(n29048));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n9646[12]), .I2(n1023_adj_4429), 
            .I3(n29046), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n27769), .O(duty_23__N_3609[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n29046), .I0(n9646[12]), .I1(n1023_adj_4429), 
            .CO(n29047));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n9646[11]), .I2(n950_adj_4428), 
            .I3(n29045), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n29045), .I0(n9646[11]), .I1(n950_adj_4428), 
            .CO(n29046));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n9646[10]), .I2(n877_adj_4427), 
            .I3(n29044), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_17 (.CI(n27892), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n27893));
    SB_CARRY mult_11_add_1225_13 (.CI(n29044), .I0(n9646[10]), .I1(n877_adj_4427), 
            .CO(n29045));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n9646[9]), .I2(n804_adj_4426), 
            .I3(n29043), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n29043), .I0(n9646[9]), .I1(n804_adj_4426), 
            .CO(n29044));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n9646[8]), .I2(n731_adj_4425), 
            .I3(n29042), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n29042), .I0(n9646[8]), .I1(n731_adj_4425), 
            .CO(n29043));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n9646[7]), .I2(n658_adj_4424), 
            .I3(n29041), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n29041), .I0(n9646[7]), .I1(n658_adj_4424), 
            .CO(n29042));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n9646[6]), .I2(n585_adj_4423), 
            .I3(n29040), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n27891), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n29040), .I0(n9646[6]), .I1(n585_adj_4423), 
            .CO(n29041));
    SB_LUT4 add_739_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n3223[20]), .I3(n27819), .O(\PID_CONTROLLER.integral_23__N_3509 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n9646[5]), .I2(n512_adj_4422), 
            .I3(n29039), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n29039), .I0(n9646[5]), .I1(n512_adj_4422), 
            .CO(n29040));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n9646[4]), .I2(n439_adj_4421), 
            .I3(n29038), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_22 (.CI(n27819), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n3223[20]), .CO(n27820));
    SB_CARRY mult_11_add_1225_7 (.CI(n29038), .I0(n9646[4]), .I1(n439_adj_4421), 
            .CO(n29039));
    SB_LUT4 add_739_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n3223[19]), .I3(n27818), .O(\PID_CONTROLLER.integral_23__N_3509 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n27891), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n27892));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n9646[3]), .I2(n366_adj_4420), 
            .I3(n29037), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n29037), .I0(n9646[3]), .I1(n366_adj_4420), 
            .CO(n29038));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n9646[2]), .I2(n293_adj_4419), 
            .I3(n29036), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n29036), .I0(n9646[2]), .I1(n293_adj_4419), 
            .CO(n29037));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n9646[1]), .I2(n220_adj_4418), 
            .I3(n29035), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n29035), .I0(n9646[1]), .I1(n220_adj_4418), 
            .CO(n29036));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n27890), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_21 (.CI(n27818), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n3223[19]), .CO(n27819));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n9646[0]), .I2(n147_adj_4417), 
            .I3(n29034), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n27890), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n27891));
    SB_LUT4 add_739_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n3223[18]), .I3(n27817), .O(\PID_CONTROLLER.integral_23__N_3509 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n29034), .I0(n9646[0]), .I1(n147_adj_4417), 
            .CO(n29035));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4416), .I2(n74_adj_4414), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4416), .I1(n74_adj_4414), 
            .CO(n29034));
    SB_LUT4 add_5225_23_lut (.I0(GND_net), .I1(n9670[20]), .I2(GND_net), 
            .I3(n29033), .O(n9646[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5225_22_lut (.I0(GND_net), .I1(n9670[19]), .I2(GND_net), 
            .I3(n29032), .O(n9646[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_22 (.CI(n29032), .I0(n9670[19]), .I1(GND_net), .CO(n29033));
    SB_LUT4 add_5225_21_lut (.I0(GND_net), .I1(n9670[18]), .I2(GND_net), 
            .I3(n29031), .O(n9646[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_20 (.CI(n27817), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n3223[18]), .CO(n27818));
    SB_CARRY add_5225_21 (.CI(n29031), .I0(n9670[18]), .I1(GND_net), .CO(n29032));
    SB_LUT4 add_5225_20_lut (.I0(GND_net), .I1(n9670[17]), .I2(GND_net), 
            .I3(n29030), .O(n9646[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_20 (.CI(n29030), .I0(n9670[17]), .I1(GND_net), .CO(n29031));
    SB_CARRY add_12_15 (.CI(n27769), .I0(n106[13]), .I1(n155[13]), .CO(n27770));
    SB_LUT4 add_5225_19_lut (.I0(GND_net), .I1(n9670[16]), .I2(GND_net), 
            .I3(n29029), .O(n9646[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_19 (.CI(n29029), .I0(n9670[16]), .I1(GND_net), .CO(n29030));
    SB_LUT4 add_5225_18_lut (.I0(GND_net), .I1(n9670[15]), .I2(GND_net), 
            .I3(n29028), .O(n9646[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_18 (.CI(n29028), .I0(n9670[15]), .I1(GND_net), .CO(n29029));
    SB_LUT4 add_5225_17_lut (.I0(GND_net), .I1(n9670[14]), .I2(GND_net), 
            .I3(n29027), .O(n9646[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_17 (.CI(n29027), .I0(n9670[14]), .I1(GND_net), .CO(n29028));
    SB_LUT4 add_5225_16_lut (.I0(GND_net), .I1(n9670[13]), .I2(n1099_adj_4411), 
            .I3(n29026), .O(n9646[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_16 (.CI(n29026), .I0(n9670[13]), .I1(n1099_adj_4411), 
            .CO(n29027));
    SB_LUT4 add_5225_15_lut (.I0(GND_net), .I1(n9670[12]), .I2(n1026_adj_4410), 
            .I3(n29025), .O(n9646[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_15 (.CI(n29025), .I0(n9670[12]), .I1(n1026_adj_4410), 
            .CO(n29026));
    SB_LUT4 add_5225_14_lut (.I0(GND_net), .I1(n9670[11]), .I2(n953_adj_4409), 
            .I3(n29024), .O(n9646[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_14 (.CI(n29024), .I0(n9670[11]), .I1(n953_adj_4409), 
            .CO(n29025));
    SB_LUT4 add_5225_13_lut (.I0(GND_net), .I1(n9670[10]), .I2(n880_adj_4408), 
            .I3(n29023), .O(n9646[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_13 (.CI(n29023), .I0(n9670[10]), .I1(n880_adj_4408), 
            .CO(n29024));
    SB_LUT4 add_5225_12_lut (.I0(GND_net), .I1(n9670[9]), .I2(n807_adj_4407), 
            .I3(n29022), .O(n9646[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_12 (.CI(n29022), .I0(n9670[9]), .I1(n807_adj_4407), 
            .CO(n29023));
    SB_LUT4 add_5225_11_lut (.I0(GND_net), .I1(n9670[8]), .I2(n734_adj_4406), 
            .I3(n29021), .O(n9646[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_11 (.CI(n29021), .I0(n9670[8]), .I1(n734_adj_4406), 
            .CO(n29022));
    SB_LUT4 add_5225_10_lut (.I0(GND_net), .I1(n9670[7]), .I2(n661_adj_4405), 
            .I3(n29020), .O(n9646[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_10 (.CI(n29020), .I0(n9670[7]), .I1(n661_adj_4405), 
            .CO(n29021));
    SB_LUT4 add_5225_9_lut (.I0(GND_net), .I1(n9670[6]), .I2(n588_adj_4404), 
            .I3(n29019), .O(n9646[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_9 (.CI(n29019), .I0(n9670[6]), .I1(n588_adj_4404), 
            .CO(n29020));
    SB_LUT4 add_5225_8_lut (.I0(GND_net), .I1(n9670[5]), .I2(n515_adj_4403), 
            .I3(n29018), .O(n9646[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n27889), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_8 (.CI(n29018), .I0(n9670[5]), .I1(n515_adj_4403), 
            .CO(n29019));
    SB_LUT4 add_5225_7_lut (.I0(GND_net), .I1(n9670[4]), .I2(n442_adj_4401), 
            .I3(n29017), .O(n9646[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_7 (.CI(n29017), .I0(n9670[4]), .I1(n442_adj_4401), 
            .CO(n29018));
    SB_LUT4 add_5225_6_lut (.I0(GND_net), .I1(n9670[3]), .I2(n369_adj_4399), 
            .I3(n29016), .O(n9646[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_6 (.CI(n29016), .I0(n9670[3]), .I1(n369_adj_4399), 
            .CO(n29017));
    SB_LUT4 add_5225_5_lut (.I0(GND_net), .I1(n9670[2]), .I2(n296_adj_4398), 
            .I3(n29015), .O(n9646[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_5 (.CI(n29015), .I0(n9670[2]), .I1(n296_adj_4398), 
            .CO(n29016));
    SB_LUT4 add_5225_4_lut (.I0(GND_net), .I1(n9670[1]), .I2(n223_adj_4397), 
            .I3(n29014), .O(n9646[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n3223[17]), .I3(n27816), .O(\PID_CONTROLLER.integral_23__N_3509 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_4 (.CI(n29014), .I0(n9670[1]), .I1(n223_adj_4397), 
            .CO(n29015));
    SB_CARRY sub_3_add_2_14 (.CI(n27889), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n27890));
    SB_LUT4 add_5225_3_lut (.I0(GND_net), .I1(n9670[0]), .I2(n150_adj_4396), 
            .I3(n29013), .O(n9646[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n27888), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_3 (.CI(n29013), .I0(n9670[0]), .I1(n150_adj_4396), 
            .CO(n29014));
    SB_LUT4 add_5225_2_lut (.I0(GND_net), .I1(n8_adj_4394), .I2(n77_adj_4393), 
            .I3(GND_net), .O(n9646[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5225_2 (.CI(GND_net), .I0(n8_adj_4394), .I1(n77_adj_4393), 
            .CO(n29013));
    SB_LUT4 add_5219_7_lut (.I0(GND_net), .I1(n34155), .I2(n490_adj_4382), 
            .I3(n29012), .O(n9613[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5219_6_lut (.I0(GND_net), .I1(n9621[3]), .I2(n417_adj_4376), 
            .I3(n29011), .O(n9613[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_6 (.CI(n29011), .I0(n9621[3]), .I1(n417_adj_4376), 
            .CO(n29012));
    SB_LUT4 add_5219_5_lut (.I0(GND_net), .I1(n9621[2]), .I2(n344_adj_4375), 
            .I3(n29010), .O(n9613[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_5 (.CI(n29010), .I0(n9621[2]), .I1(n344_adj_4375), 
            .CO(n29011));
    SB_LUT4 add_5219_4_lut (.I0(GND_net), .I1(n9621[1]), .I2(n271_adj_4374), 
            .I3(n29009), .O(n9613[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_4 (.CI(n29009), .I0(n9621[1]), .I1(n271_adj_4374), 
            .CO(n29010));
    SB_LUT4 add_5219_3_lut (.I0(GND_net), .I1(n9621[0]), .I2(n198_adj_4373), 
            .I3(n29008), .O(n9613[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_13 (.CI(n27888), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n27889));
    SB_CARRY add_5219_3 (.CI(n29008), .I0(n9621[0]), .I1(n198_adj_4373), 
            .CO(n29009));
    SB_LUT4 add_5219_2_lut (.I0(GND_net), .I1(n56_adj_4372), .I2(n125_adj_4370), 
            .I3(GND_net), .O(n9613[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5219_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5219_2 (.CI(GND_net), .I0(n56_adj_4372), .I1(n125_adj_4370), 
            .CO(n29008));
    SB_LUT4 add_5218_8_lut (.I0(GND_net), .I1(n9613[5]), .I2(n560_adj_4369), 
            .I3(n29007), .O(n9604[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_19 (.CI(n27816), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n3223[17]), .CO(n27817));
    SB_LUT4 add_5218_7_lut (.I0(GND_net), .I1(n9613[4]), .I2(n487_adj_4368), 
            .I3(n29006), .O(n9604[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5218_7 (.CI(n29006), .I0(n9613[4]), .I1(n487_adj_4368), 
            .CO(n29007));
    SB_LUT4 add_5218_6_lut (.I0(GND_net), .I1(n9613[3]), .I2(n414_adj_4367), 
            .I3(n29005), .O(n9604[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_6 (.CI(n29005), .I0(n9613[3]), .I1(n414_adj_4367), 
            .CO(n29006));
    SB_LUT4 add_5218_5_lut (.I0(GND_net), .I1(n9613[2]), .I2(n341_adj_4366), 
            .I3(n29004), .O(n9604[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_5 (.CI(n29004), .I0(n9613[2]), .I1(n341_adj_4366), 
            .CO(n29005));
    SB_LUT4 add_5218_4_lut (.I0(GND_net), .I1(n9613[1]), .I2(n268_adj_4365), 
            .I3(n29003), .O(n9604[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_4 (.CI(n29003), .I0(n9613[1]), .I1(n268_adj_4365), 
            .CO(n29004));
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4649));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5218_3_lut (.I0(GND_net), .I1(n9613[0]), .I2(n195_adj_4364), 
            .I3(n29002), .O(n9604[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3485[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5218_3 (.CI(n29002), .I0(n9613[0]), .I1(n195_adj_4364), 
            .CO(n29003));
    SB_LUT4 add_739_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n3223[16]), .I3(n27815), .O(\PID_CONTROLLER.integral_23__N_3509 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5218_2_lut (.I0(GND_net), .I1(n53_adj_4363), .I2(n122_adj_4361), 
            .I3(GND_net), .O(n9604[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5218_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5218_2 (.CI(GND_net), .I0(n53_adj_4363), .I1(n122_adj_4361), 
            .CO(n29002));
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n27887), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5217_9_lut (.I0(GND_net), .I1(n9604[6]), .I2(n630_adj_4360), 
            .I3(n29001), .O(n9594[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3485[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3485[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3485[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3485[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3485[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3485[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3485[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3485[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3485[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3485[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3485[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3485[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3485[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3485[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3485[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3485[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3485[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3485[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3485[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3485[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3485[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3509 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5217_8_lut (.I0(GND_net), .I1(n9604[5]), .I2(n557_adj_4355), 
            .I3(n29000), .O(n9594[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_8 (.CI(n29000), .I0(n9604[5]), .I1(n557_adj_4355), 
            .CO(n29001));
    SB_LUT4 add_5217_7_lut (.I0(GND_net), .I1(n9604[4]), .I2(n484_adj_4354), 
            .I3(n28999), .O(n9594[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_7 (.CI(n28999), .I0(n9604[4]), .I1(n484_adj_4354), 
            .CO(n29000));
    SB_LUT4 add_5217_6_lut (.I0(GND_net), .I1(n9604[3]), .I2(n411_adj_4353), 
            .I3(n28998), .O(n9594[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_6 (.CI(n28998), .I0(n9604[3]), .I1(n411_adj_4353), 
            .CO(n28999));
    SB_LUT4 add_5217_5_lut (.I0(GND_net), .I1(n9604[2]), .I2(n338_adj_4352), 
            .I3(n28997), .O(n9594[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4650));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5217_5 (.CI(n28997), .I0(n9604[2]), .I1(n338_adj_4352), 
            .CO(n28998));
    SB_LUT4 add_5217_4_lut (.I0(GND_net), .I1(n9604[1]), .I2(n265_adj_4351), 
            .I3(n28996), .O(n9594[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_4 (.CI(n28996), .I0(n9604[1]), .I1(n265_adj_4351), 
            .CO(n28997));
    SB_LUT4 add_5217_3_lut (.I0(GND_net), .I1(n9604[0]), .I2(n192_adj_4349), 
            .I3(n28995), .O(n9594[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_3 (.CI(n28995), .I0(n9604[0]), .I1(n192_adj_4349), 
            .CO(n28996));
    SB_LUT4 add_5217_2_lut (.I0(GND_net), .I1(n50_adj_4348), .I2(n119_adj_4347), 
            .I3(GND_net), .O(n9594[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5217_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5217_2 (.CI(GND_net), .I0(n50_adj_4348), .I1(n119_adj_4347), 
            .CO(n28995));
    SB_LUT4 add_5216_10_lut (.I0(GND_net), .I1(n9594[7]), .I2(n700_adj_4346), 
            .I3(n28994), .O(n9583[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5216_9_lut (.I0(GND_net), .I1(n9594[6]), .I2(n627_adj_4345), 
            .I3(n28993), .O(n9583[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_9 (.CI(n28993), .I0(n9594[6]), .I1(n627_adj_4345), 
            .CO(n28994));
    SB_LUT4 add_5216_8_lut (.I0(GND_net), .I1(n9594[5]), .I2(n554_adj_4339), 
            .I3(n28992), .O(n9583[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_8 (.CI(n28992), .I0(n9594[5]), .I1(n554_adj_4339), 
            .CO(n28993));
    SB_LUT4 add_5216_7_lut (.I0(GND_net), .I1(n9594[4]), .I2(n481_adj_4338), 
            .I3(n28991), .O(n9583[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_7 (.CI(n28991), .I0(n9594[4]), .I1(n481_adj_4338), 
            .CO(n28992));
    SB_LUT4 add_5216_6_lut (.I0(GND_net), .I1(n9594[3]), .I2(n408_adj_4337), 
            .I3(n28990), .O(n9583[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_6 (.CI(n28990), .I0(n9594[3]), .I1(n408_adj_4337), 
            .CO(n28991));
    SB_LUT4 add_5216_5_lut (.I0(GND_net), .I1(n9594[2]), .I2(n335_adj_4336), 
            .I3(n28989), .O(n9583[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_18 (.CI(n27815), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n3223[16]), .CO(n27816));
    SB_CARRY sub_3_add_2_12 (.CI(n27887), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n27888));
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n27886), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_5 (.CI(n28989), .I0(n9594[2]), .I1(n335_adj_4336), 
            .CO(n28990));
    SB_LUT4 add_5216_4_lut (.I0(GND_net), .I1(n9594[1]), .I2(n262_adj_4335), 
            .I3(n28988), .O(n9583[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_4 (.CI(n28988), .I0(n9594[1]), .I1(n262_adj_4335), 
            .CO(n28989));
    SB_LUT4 add_5216_3_lut (.I0(GND_net), .I1(n9594[0]), .I2(n189_adj_4334), 
            .I3(n28987), .O(n9583[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4651));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5216_3 (.CI(n28987), .I0(n9594[0]), .I1(n189_adj_4334), 
            .CO(n28988));
    SB_LUT4 add_5216_2_lut (.I0(GND_net), .I1(n47_adj_4333), .I2(n116_adj_4332), 
            .I3(GND_net), .O(n9583[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5216_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5216_2 (.CI(GND_net), .I0(n47_adj_4333), .I1(n116_adj_4332), 
            .CO(n28987));
    SB_LUT4 add_5215_11_lut (.I0(GND_net), .I1(n9583[8]), .I2(n770_adj_4331), 
            .I3(n28986), .O(n9571[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5215_10_lut (.I0(GND_net), .I1(n9583[7]), .I2(n697_adj_4330), 
            .I3(n28985), .O(n9571[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_10 (.CI(n28985), .I0(n9583[7]), .I1(n697_adj_4330), 
            .CO(n28986));
    SB_LUT4 add_5215_9_lut (.I0(GND_net), .I1(n9583[6]), .I2(n624_adj_4328), 
            .I3(n28984), .O(n9571[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_9 (.CI(n28984), .I0(n9583[6]), .I1(n624_adj_4328), 
            .CO(n28985));
    SB_LUT4 add_5215_8_lut (.I0(GND_net), .I1(n9583[5]), .I2(n551_adj_4327), 
            .I3(n28983), .O(n9571[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_8 (.CI(n28983), .I0(n9583[5]), .I1(n551_adj_4327), 
            .CO(n28984));
    SB_LUT4 add_5215_7_lut (.I0(GND_net), .I1(n9583[4]), .I2(n478_adj_4325), 
            .I3(n28982), .O(n9571[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n3223[15]), .I3(n27814), .O(\PID_CONTROLLER.integral_23__N_3509 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_7 (.CI(n28982), .I0(n9583[4]), .I1(n478_adj_4325), 
            .CO(n28983));
    SB_LUT4 add_5215_6_lut (.I0(GND_net), .I1(n9583[3]), .I2(n405_adj_4322), 
            .I3(n28981), .O(n9571[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_17 (.CI(n27814), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n3223[15]), .CO(n27815));
    SB_CARRY add_5215_6 (.CI(n28981), .I0(n9583[3]), .I1(n405_adj_4322), 
            .CO(n28982));
    SB_CARRY sub_3_add_2_11 (.CI(n27886), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n27887));
    SB_LUT4 add_5215_5_lut (.I0(GND_net), .I1(n9583[2]), .I2(n332_adj_4321), 
            .I3(n28980), .O(n9571[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_5 (.CI(n28980), .I0(n9583[2]), .I1(n332_adj_4321), 
            .CO(n28981));
    SB_LUT4 add_5215_4_lut (.I0(GND_net), .I1(n9583[1]), .I2(n259_adj_4320), 
            .I3(n28979), .O(n9571[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_4 (.CI(n28979), .I0(n9583[1]), .I1(n259_adj_4320), 
            .CO(n28980));
    SB_LUT4 add_5215_3_lut (.I0(GND_net), .I1(n9583[0]), .I2(n186_adj_4319), 
            .I3(n28978), .O(n9571[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n27885), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_3 (.CI(n28978), .I0(n9583[0]), .I1(n186_adj_4319), 
            .CO(n28979));
    SB_CARRY sub_3_add_2_10 (.CI(n27885), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n27886));
    SB_LUT4 add_5215_2_lut (.I0(GND_net), .I1(n44_adj_4318), .I2(n113_adj_4317), 
            .I3(GND_net), .O(n9571[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_2 (.CI(GND_net), .I0(n44_adj_4318), .I1(n113_adj_4317), 
            .CO(n28978));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n27768), .O(duty_23__N_3609[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_12_lut (.I0(GND_net), .I1(n9571[9]), .I2(n840_adj_4316), 
            .I3(n28977), .O(n9558[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n27768), .I0(n106[12]), .I1(n155[12]), .CO(n27769));
    SB_LUT4 add_5214_11_lut (.I0(GND_net), .I1(n9571[8]), .I2(n767_adj_4315), 
            .I3(n28976), .O(n9558[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_11 (.CI(n28976), .I0(n9571[8]), .I1(n767_adj_4315), 
            .CO(n28977));
    SB_LUT4 add_5214_10_lut (.I0(GND_net), .I1(n9571[7]), .I2(n694_adj_4313), 
            .I3(n28975), .O(n9558[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_10 (.CI(n28975), .I0(n9571[7]), .I1(n694_adj_4313), 
            .CO(n28976));
    SB_LUT4 add_5214_9_lut (.I0(GND_net), .I1(n9571[6]), .I2(n621_adj_4312), 
            .I3(n28974), .O(n9558[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n3223[14]), .I3(n27813), .O(\PID_CONTROLLER.integral_23__N_3509 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_9 (.CI(n28974), .I0(n9571[6]), .I1(n621_adj_4312), 
            .CO(n28975));
    SB_LUT4 add_5214_8_lut (.I0(GND_net), .I1(n9571[5]), .I2(n548_adj_4310), 
            .I3(n28973), .O(n9558[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_8 (.CI(n28973), .I0(n9571[5]), .I1(n548_adj_4310), 
            .CO(n28974));
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4653));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n27884), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5214_7_lut (.I0(GND_net), .I1(n9571[4]), .I2(n475_adj_4308), 
            .I3(n28972), .O(n9558[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_7 (.CI(n28972), .I0(n9571[4]), .I1(n475_adj_4308), 
            .CO(n28973));
    SB_LUT4 add_5214_6_lut (.I0(GND_net), .I1(n9571[3]), .I2(n402_adj_4307), 
            .I3(n28971), .O(n9558[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_6 (.CI(n28971), .I0(n9571[3]), .I1(n402_adj_4307), 
            .CO(n28972));
    SB_LUT4 add_5214_5_lut (.I0(GND_net), .I1(n9571[2]), .I2(n329_adj_4306), 
            .I3(n28970), .O(n9558[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_5 (.CI(n28970), .I0(n9571[2]), .I1(n329_adj_4306), 
            .CO(n28971));
    SB_LUT4 add_5214_4_lut (.I0(GND_net), .I1(n9571[1]), .I2(n256_adj_4305), 
            .I3(n28969), .O(n9558[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_9 (.CI(n27884), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n27885));
    SB_CARRY add_5214_4 (.CI(n28969), .I0(n9571[1]), .I1(n256_adj_4305), 
            .CO(n28970));
    SB_LUT4 add_5214_3_lut (.I0(GND_net), .I1(n9571[0]), .I2(n183_adj_4304), 
            .I3(n28968), .O(n9558[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_3 (.CI(n28968), .I0(n9571[0]), .I1(n183_adj_4304), 
            .CO(n28969));
    SB_LUT4 add_5214_2_lut (.I0(GND_net), .I1(n41_adj_4303), .I2(n110_adj_4302), 
            .I3(GND_net), .O(n9558[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5214_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5214_2 (.CI(GND_net), .I0(n41_adj_4303), .I1(n110_adj_4302), 
            .CO(n28968));
    SB_LUT4 add_5213_13_lut (.I0(GND_net), .I1(n9558[10]), .I2(n910_adj_4300), 
            .I3(n28967), .O(n9544[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5213_12_lut (.I0(GND_net), .I1(n9558[9]), .I2(n837_adj_4299), 
            .I3(n28966), .O(n9544[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_12 (.CI(n28966), .I0(n9558[9]), .I1(n837_adj_4299), 
            .CO(n28967));
    SB_LUT4 add_5213_11_lut (.I0(GND_net), .I1(n9558[8]), .I2(n764_adj_4298), 
            .I3(n28965), .O(n9544[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_11 (.CI(n28965), .I0(n9558[8]), .I1(n764_adj_4298), 
            .CO(n28966));
    SB_LUT4 add_5213_10_lut (.I0(GND_net), .I1(n9558[7]), .I2(n691_adj_4297), 
            .I3(n28964), .O(n9544[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n27767), .O(duty_23__N_3609[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_10 (.CI(n28964), .I0(n9558[7]), .I1(n691_adj_4297), 
            .CO(n28965));
    SB_LUT4 add_5213_9_lut (.I0(GND_net), .I1(n9558[6]), .I2(n618_adj_4296), 
            .I3(n28963), .O(n9544[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_9 (.CI(n28963), .I0(n9558[6]), .I1(n618_adj_4296), 
            .CO(n28964));
    SB_LUT4 add_5213_8_lut (.I0(GND_net), .I1(n9558[5]), .I2(n545), .I3(n28962), 
            .O(n9544[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_8 (.CI(n28962), .I0(n9558[5]), .I1(n545), .CO(n28963));
    SB_LUT4 add_5213_7_lut (.I0(GND_net), .I1(n9558[4]), .I2(n472), .I3(n28961), 
            .O(n9544[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_7 (.CI(n28961), .I0(n9558[4]), .I1(n472), .CO(n28962));
    SB_LUT4 add_5213_6_lut (.I0(GND_net), .I1(n9558[3]), .I2(n399), .I3(n28960), 
            .O(n9544[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_6 (.CI(n28960), .I0(n9558[3]), .I1(n399), .CO(n28961));
    SB_LUT4 add_5213_5_lut (.I0(GND_net), .I1(n9558[2]), .I2(n326), .I3(n28959), 
            .O(n9544[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_5 (.CI(n28959), .I0(n9558[2]), .I1(n326), .CO(n28960));
    SB_CARRY add_12_13 (.CI(n27767), .I0(n106[11]), .I1(n155[11]), .CO(n27768));
    SB_LUT4 add_5213_4_lut (.I0(GND_net), .I1(n9558[1]), .I2(n253), .I3(n28958), 
            .O(n9544[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_4 (.CI(n28958), .I0(n9558[1]), .I1(n253), .CO(n28959));
    SB_LUT4 add_5213_3_lut (.I0(GND_net), .I1(n9558[0]), .I2(n180), .I3(n28957), 
            .O(n9544[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_3 (.CI(n28957), .I0(n9558[0]), .I1(n180), .CO(n28958));
    SB_LUT4 add_5213_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n9544[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5213_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n27883), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5213_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n28957));
    SB_LUT4 add_5212_14_lut (.I0(GND_net), .I1(n9544[11]), .I2(n980), 
            .I3(n28956), .O(n9529[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5212_13_lut (.I0(GND_net), .I1(n9544[10]), .I2(n907), 
            .I3(n28955), .O(n9529[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_13 (.CI(n28955), .I0(n9544[10]), .I1(n907), .CO(n28956));
    SB_CARRY add_739_16 (.CI(n27813), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n3223[14]), .CO(n27814));
    SB_LUT4 add_5212_12_lut (.I0(GND_net), .I1(n9544[9]), .I2(n834), .I3(n28954), 
            .O(n9529[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_12 (.CI(n28954), .I0(n9544[9]), .I1(n834), .CO(n28955));
    SB_LUT4 add_739_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n3223[13]), .I3(n27812), .O(\PID_CONTROLLER.integral_23__N_3509 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5212_11_lut (.I0(GND_net), .I1(n9544[8]), .I2(n761), .I3(n28953), 
            .O(n9529[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_11 (.CI(n28953), .I0(n9544[8]), .I1(n761), .CO(n28954));
    SB_LUT4 add_5212_10_lut (.I0(GND_net), .I1(n9544[7]), .I2(n688), .I3(n28952), 
            .O(n9529[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_10 (.CI(n28952), .I0(n9544[7]), .I1(n688), .CO(n28953));
    SB_LUT4 add_5212_9_lut (.I0(GND_net), .I1(n9544[6]), .I2(n615), .I3(n28951), 
            .O(n9529[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_9 (.CI(n28951), .I0(n9544[6]), .I1(n615), .CO(n28952));
    SB_CARRY add_739_15 (.CI(n27812), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n3223[13]), .CO(n27813));
    SB_LUT4 add_5212_8_lut (.I0(GND_net), .I1(n9544[5]), .I2(n542), .I3(n28950), 
            .O(n9529[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_8 (.CI(n28950), .I0(n9544[5]), .I1(n542), .CO(n28951));
    SB_LUT4 add_5212_7_lut (.I0(GND_net), .I1(n9544[4]), .I2(n469), .I3(n28949), 
            .O(n9529[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_7 (.CI(n28949), .I0(n9544[4]), .I1(n469), .CO(n28950));
    SB_LUT4 add_5212_6_lut (.I0(GND_net), .I1(n9544[3]), .I2(n396), .I3(n28948), 
            .O(n9529[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_6 (.CI(n28948), .I0(n9544[3]), .I1(n396), .CO(n28949));
    SB_LUT4 add_5212_5_lut (.I0(GND_net), .I1(n9544[2]), .I2(n323), .I3(n28947), 
            .O(n9529[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_5 (.CI(n28947), .I0(n9544[2]), .I1(n323), .CO(n28948));
    SB_LUT4 add_5212_4_lut (.I0(GND_net), .I1(n9544[1]), .I2(n250), .I3(n28946), 
            .O(n9529[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4654));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4655));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4656));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4657));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4659));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19399_2_lut (.I0(n28[23]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19399_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968_adj_4660));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_8 (.CI(n27883), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n27884));
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n27882), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n27766), .O(duty_23__N_3609[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041_adj_4661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114_adj_4662));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_739_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n3223[12]), .I3(n27811), .O(\PID_CONTROLLER.integral_23__N_3509 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n27766), .I0(n106[10]), .I1(n155[10]), .CO(n27767));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n27765), 
            .O(duty_23__N_3609[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_14 (.CI(n27811), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n3223[12]), .CO(n27812));
    SB_LUT4 add_739_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n3223[11]), .I3(n27810), .O(\PID_CONTROLLER.integral_23__N_3509 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_4 (.CI(n28946), .I0(n9544[1]), .I1(n250), .CO(n28947));
    SB_LUT4 add_5212_3_lut (.I0(GND_net), .I1(n9544[0]), .I2(n177), .I3(n28945), 
            .O(n9529[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5212_3 (.CI(n28945), .I0(n9544[0]), .I1(n177), .CO(n28946));
    SB_LUT4 add_5212_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n9529[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5212_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n27765), .I0(n106[9]), .I1(n155[9]), .CO(n27766));
    SB_CARRY add_5212_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n28945));
    SB_LUT4 add_5211_15_lut (.I0(GND_net), .I1(n9529[12]), .I2(n1050), 
            .I3(n28944), .O(n9513[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5211_14_lut (.I0(GND_net), .I1(n9529[11]), .I2(n977), 
            .I3(n28943), .O(n9513[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_14 (.CI(n28943), .I0(n9529[11]), .I1(n977), .CO(n28944));
    SB_CARRY sub_3_add_2_7 (.CI(n27882), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n27883));
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n27881), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n27764), 
            .O(duty_23__N_3609[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n27764), .I0(n106[8]), .I1(n155[8]), .CO(n27765));
    SB_CARRY add_739_13 (.CI(n27810), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n3223[11]), .CO(n27811));
    SB_CARRY sub_3_add_2_6 (.CI(n27881), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n27882));
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4638));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n27880), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4637));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_739_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n3223[10]), .I3(n27809), .O(\PID_CONTROLLER.integral_23__N_3509 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_12 (.CI(n27809), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n3223[10]), .CO(n27810));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n27763), 
            .O(duty_23__N_3609[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_9 (.CI(n27763), .I0(n106[7]), .I1(n155[7]), .CO(n27764));
    SB_LUT4 add_739_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n3223[9]), .I3(n27808), .O(\PID_CONTROLLER.integral_23__N_3509 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4636));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5211_13_lut (.I0(GND_net), .I1(n9529[10]), .I2(n904), 
            .I3(n28942), .O(n9513[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_11 (.CI(n27808), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n3223[9]), .CO(n27809));
    SB_CARRY sub_3_add_2_5 (.CI(n27880), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n27881));
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4635));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4634));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5211_13 (.CI(n28942), .I0(n9529[10]), .I1(n904), .CO(n28943));
    SB_LUT4 add_5211_12_lut (.I0(GND_net), .I1(n9529[9]), .I2(n831), .I3(n28941), 
            .O(n9513[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_12 (.CI(n28941), .I0(n9529[9]), .I1(n831), .CO(n28942));
    SB_LUT4 add_5211_11_lut (.I0(GND_net), .I1(n9529[8]), .I2(n758), .I3(n28940), 
            .O(n9513[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_11 (.CI(n28940), .I0(n9529[8]), .I1(n758), .CO(n28941));
    SB_LUT4 add_5211_10_lut (.I0(GND_net), .I1(n9529[7]), .I2(n685), .I3(n28939), 
            .O(n9513[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_10 (.CI(n28939), .I0(n9529[7]), .I1(n685), .CO(n28940));
    SB_LUT4 add_5211_9_lut (.I0(GND_net), .I1(n9529[6]), .I2(n612), .I3(n28938), 
            .O(n9513[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_9 (.CI(n28938), .I0(n9529[6]), .I1(n612), .CO(n28939));
    SB_LUT4 add_5211_8_lut (.I0(GND_net), .I1(n9529[5]), .I2(n539), .I3(n28937), 
            .O(n9513[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n27879), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_4 (.CI(n27879), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n27880));
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n27878), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n27878), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n27879));
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4633));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4632));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4631));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4629));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5211_8 (.CI(n28937), .I0(n9529[5]), .I1(n539), .CO(n28938));
    SB_LUT4 add_5211_7_lut (.I0(GND_net), .I1(n9529[4]), .I2(n466), .I3(n28936), 
            .O(n9513[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_7 (.CI(n28936), .I0(n9529[4]), .I1(n466), .CO(n28937));
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n27762), 
            .O(duty_23__N_3609[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5211_6_lut (.I0(GND_net), .I1(n9529[3]), .I2(n393), .I3(n28935), 
            .O(n9513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4665));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4628));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4666));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4626));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4625));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4668));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4623));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4669));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4622));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4620));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533_adj_4671));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606_adj_4672));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19377_2_lut (.I0(n28[1]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4674));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4675));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4619));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5211_6 (.CI(n28935), .I0(n9529[3]), .I1(n393), .CO(n28936));
    SB_LUT4 add_5211_5_lut (.I0(GND_net), .I1(n9529[2]), .I2(n320_adj_4676), 
            .I3(n28934), .O(n9513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n27878));
    SB_CARRY add_5211_5 (.CI(n28934), .I0(n9529[2]), .I1(n320_adj_4676), 
            .CO(n28935));
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5211_4_lut (.I0(GND_net), .I1(n9529[1]), .I2(n247_adj_4677), 
            .I3(n28933), .O(n9513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4617));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4616));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4614));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_8 (.CI(n27762), .I0(n106[6]), .I1(n155[6]), .CO(n27763));
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n27761), 
            .O(duty_23__N_3609[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n3223[8]), .I3(n27807), .O(\PID_CONTROLLER.integral_23__N_3509 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_4 (.CI(n28933), .I0(n9529[1]), .I1(n247_adj_4677), 
            .CO(n28934));
    SB_CARRY add_739_10 (.CI(n27807), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n3223[8]), .CO(n27808));
    SB_LUT4 add_5211_3_lut (.I0(GND_net), .I1(n9529[0]), .I2(n174_adj_4678), 
            .I3(n28932), .O(n9513[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n3223[7]), .I3(n27806), .O(\PID_CONTROLLER.integral_23__N_3509 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n27761), .I0(n106[5]), .I1(n155[5]), .CO(n27762));
    SB_CARRY add_739_9 (.CI(n27806), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n3223[7]), .CO(n27807));
    SB_LUT4 add_739_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n3223[6]), .I3(n27805), .O(\PID_CONTROLLER.integral_23__N_3509 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_3 (.CI(n28932), .I0(n9529[0]), .I1(n174_adj_4678), 
            .CO(n28933));
    SB_CARRY add_739_8 (.CI(n27805), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n3223[6]), .CO(n27806));
    SB_LUT4 add_5211_2_lut (.I0(GND_net), .I1(n32_adj_4679), .I2(n101_adj_4680), 
            .I3(GND_net), .O(n9513[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5211_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n3223[5]), .I3(n27804), .O(\PID_CONTROLLER.integral_23__N_3509 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n27760), 
            .O(duty_23__N_3609[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5211_2 (.CI(GND_net), .I0(n32_adj_4679), .I1(n101_adj_4680), 
            .CO(n28932));
    SB_LUT4 add_5210_16_lut (.I0(GND_net), .I1(n9513[13]), .I2(n1120_adj_4682), 
            .I3(n28931), .O(n9496[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5210_15_lut (.I0(GND_net), .I1(n9513[12]), .I2(n1047_adj_4683), 
            .I3(n28930), .O(n9496[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_7 (.CI(n27804), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n3223[5]), .CO(n27805));
    SB_CARRY add_5210_15 (.CI(n28930), .I0(n9513[12]), .I1(n1047_adj_4683), 
            .CO(n28931));
    SB_CARRY add_12_6 (.CI(n27760), .I0(n106[4]), .I1(n155[4]), .CO(n27761));
    SB_LUT4 add_739_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n3223[4]), .I3(n27803), .O(\PID_CONTROLLER.integral_23__N_3509 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n27759), 
            .O(duty_23__N_3609[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_5 (.CI(n27759), .I0(n106[3]), .I1(n155[3]), .CO(n27760));
    SB_LUT4 add_5210_14_lut (.I0(GND_net), .I1(n9513[11]), .I2(n974_adj_4684), 
            .I3(n28929), .O(n9496[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[23]), 
            .I3(n27951), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[22]), 
            .I3(n27950), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29667_3_lut_4_lut (.I0(duty_23__N_3609[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3609[2]), .O(n36063));   // verilog/motorControl.v(38[19:35])
    defparam i29667_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4611));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4610));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_739_6 (.CI(n27803), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n3223[4]), .CO(n27804));
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3609[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4499));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4608));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5210_14 (.CI(n28929), .I0(n9513[11]), .I1(n974_adj_4684), 
            .CO(n28930));
    SB_LUT4 i29703_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3609[3]), 
            .I2(duty_23__N_3609[2]), .I3(PWMLimit[2]), .O(n36099));   // verilog/motorControl.v(36[10:25])
    defparam i29703_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_739_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n3223[3]), .I3(n27802), .O(\PID_CONTROLLER.integral_23__N_3509 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3609[3]), 
            .I2(duty_23__N_3609[2]), .I3(GND_net), .O(n6_adj_4470));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4607));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_24 (.CI(n27950), .I0(GND_net), .I1(n1_adj_4708[22]), 
            .CO(n27951));
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4605));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4604));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[21]), 
            .I3(n27949), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n27949), .I0(GND_net), .I1(n1_adj_4708[21]), 
            .CO(n27950));
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4602));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_739_5 (.CI(n27802), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n3223[3]), .CO(n27803));
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4601));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4599));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n27758), 
            .O(duty_23__N_3609[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5210_13_lut (.I0(GND_net), .I1(n9513[10]), .I2(n901_adj_4688), 
            .I3(n28928), .O(n9496[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_13 (.CI(n28928), .I0(n9513[10]), .I1(n901_adj_4688), 
            .CO(n28929));
    SB_LUT4 add_739_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n3223[2]), .I3(n27801), .O(\PID_CONTROLLER.integral_23__N_3509 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5210_12_lut (.I0(GND_net), .I1(n9513[9]), .I2(n828_adj_4689), 
            .I3(n28927), .O(n9496[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n27758), .I0(n106[2]), .I1(n155[2]), .CO(n27759));
    SB_CARRY add_5210_12 (.CI(n28927), .I0(n9513[9]), .I1(n828_adj_4689), 
            .CO(n28928));
    SB_LUT4 add_5210_11_lut (.I0(GND_net), .I1(n9513[8]), .I2(n755_adj_4690), 
            .I3(n28926), .O(n9496[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_11 (.CI(n28926), .I0(n9513[8]), .I1(n755_adj_4690), 
            .CO(n28927));
    SB_LUT4 add_5210_10_lut (.I0(GND_net), .I1(n9513[7]), .I2(n682_adj_4691), 
            .I3(n28925), .O(n9496[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_10 (.CI(n28925), .I0(n9513[7]), .I1(n682_adj_4691), 
            .CO(n28926));
    SB_LUT4 add_5210_9_lut (.I0(GND_net), .I1(n9513[6]), .I2(n609_adj_4692), 
            .I3(n28924), .O(n9496[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_9 (.CI(n28924), .I0(n9513[6]), .I1(n609_adj_4692), 
            .CO(n28925));
    SB_LUT4 add_5210_8_lut (.I0(GND_net), .I1(n9513[5]), .I2(n536_adj_4693), 
            .I3(n28923), .O(n9496[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_8 (.CI(n28923), .I0(n9513[5]), .I1(n536_adj_4693), 
            .CO(n28924));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n27757), 
            .O(duty_23__N_3609[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4596));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5210_7_lut (.I0(GND_net), .I1(n9513[4]), .I2(n463_adj_4695), 
            .I3(n28922), .O(n9496[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_7 (.CI(n28922), .I0(n9513[4]), .I1(n463_adj_4695), 
            .CO(n28923));
    SB_LUT4 add_5210_6_lut (.I0(GND_net), .I1(n9513[3]), .I2(n390_adj_4696), 
            .I3(n28921), .O(n9496[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_6 (.CI(n28921), .I0(n9513[3]), .I1(n390_adj_4696), 
            .CO(n28922));
    SB_LUT4 add_5210_5_lut (.I0(GND_net), .I1(n9513[2]), .I2(n317_adj_4697), 
            .I3(n28920), .O(n9496[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4595));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5210_5 (.CI(n28920), .I0(n9513[2]), .I1(n317_adj_4697), 
            .CO(n28921));
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5210_4_lut (.I0(GND_net), .I1(n9513[1]), .I2(n244_adj_4698), 
            .I3(n28919), .O(n9496[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_4 (.CI(n27801), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n3223[2]), .CO(n27802));
    SB_CARRY add_5210_4 (.CI(n28919), .I0(n9513[1]), .I1(n244_adj_4698), 
            .CO(n28920));
    SB_LUT4 add_5210_3_lut (.I0(GND_net), .I1(n9513[0]), .I2(n171_adj_4699), 
            .I3(n28918), .O(n9496[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_3 (.CI(n28918), .I0(n9513[0]), .I1(n171_adj_4699), 
            .CO(n28919));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[20]), 
            .I3(n27948), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n27948), .I0(GND_net), .I1(n1_adj_4708[20]), 
            .CO(n27949));
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4593));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5210_2_lut (.I0(GND_net), .I1(n29_adj_4701), .I2(n98_adj_4702), 
            .I3(GND_net), .O(n9496[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5210_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5210_2 (.CI(GND_net), .I0(n29_adj_4701), .I1(n98_adj_4702), 
            .CO(n28918));
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4592));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5209_17_lut (.I0(GND_net), .I1(n9496[14]), .I2(GND_net), 
            .I3(n28917), .O(n9478[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5209_16_lut (.I0(GND_net), .I1(n9496[13]), .I2(n1117_adj_4703), 
            .I3(n28916), .O(n9478[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_16 (.CI(n28916), .I0(n9496[13]), .I1(n1117_adj_4703), 
            .CO(n28917));
    SB_LUT4 add_5209_15_lut (.I0(GND_net), .I1(n9496[12]), .I2(n1044_adj_4704), 
            .I3(n28915), .O(n9478[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_15 (.CI(n28915), .I0(n9496[12]), .I1(n1044_adj_4704), 
            .CO(n28916));
    SB_LUT4 add_5209_14_lut (.I0(GND_net), .I1(n9496[11]), .I2(n971_adj_4705), 
            .I3(n28914), .O(n9478[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_14 (.CI(n28914), .I0(n9496[11]), .I1(n971_adj_4705), 
            .CO(n28915));
    SB_LUT4 add_5209_13_lut (.I0(GND_net), .I1(n9496[10]), .I2(n898_adj_4706), 
            .I3(n28913), .O(n9478[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_13 (.CI(n28913), .I0(n9496[10]), .I1(n898_adj_4706), 
            .CO(n28914));
    SB_LUT4 add_5209_12_lut (.I0(GND_net), .I1(n9496[9]), .I2(n825_adj_4675), 
            .I3(n28912), .O(n9478[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_12 (.CI(n28912), .I0(n9496[9]), .I1(n825_adj_4675), 
            .CO(n28913));
    SB_LUT4 add_5209_11_lut (.I0(GND_net), .I1(n9496[8]), .I2(n752_adj_4674), 
            .I3(n28911), .O(n9478[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_11 (.CI(n28911), .I0(n9496[8]), .I1(n752_adj_4674), 
            .CO(n28912));
    SB_LUT4 add_5209_10_lut (.I0(GND_net), .I1(n9496[7]), .I2(n679_adj_4673), 
            .I3(n28910), .O(n9478[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_739_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3223[1]), .I3(n27800), .O(\PID_CONTROLLER.integral_23__N_3509 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_10 (.CI(n28910), .I0(n9496[7]), .I1(n679_adj_4673), 
            .CO(n28911));
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5209_9_lut (.I0(GND_net), .I1(n9496[6]), .I2(n606_adj_4672), 
            .I3(n28909), .O(n9478[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_9 (.CI(n28909), .I0(n9496[6]), .I1(n606_adj_4672), 
            .CO(n28910));
    SB_LUT4 add_5209_8_lut (.I0(GND_net), .I1(n9496[5]), .I2(n533_adj_4671), 
            .I3(n28908), .O(n9478[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_3 (.CI(n27800), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n3223[1]), .CO(n27801));
    SB_CARRY add_5209_8 (.CI(n28908), .I0(n9496[5]), .I1(n533_adj_4671), 
            .CO(n28909));
    SB_LUT4 add_5209_7_lut (.I0(GND_net), .I1(n9496[4]), .I2(n460_adj_4670), 
            .I3(n28907), .O(n9478[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4590));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5209_7 (.CI(n28907), .I0(n9496[4]), .I1(n460_adj_4670), 
            .CO(n28908));
    SB_LUT4 add_5209_6_lut (.I0(GND_net), .I1(n9496[3]), .I2(n387_adj_4669), 
            .I3(n28906), .O(n9478[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_6 (.CI(n28906), .I0(n9496[3]), .I1(n387_adj_4669), 
            .CO(n28907));
    SB_LUT4 add_5209_5_lut (.I0(GND_net), .I1(n9496[2]), .I2(n314_adj_4668), 
            .I3(n28905), .O(n9478[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_5 (.CI(n28905), .I0(n9496[2]), .I1(n314_adj_4668), 
            .CO(n28906));
    SB_LUT4 add_5209_4_lut (.I0(GND_net), .I1(n9496[1]), .I2(n241_adj_4667), 
            .I3(n28904), .O(n9478[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4589));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5209_4 (.CI(n28904), .I0(n9496[1]), .I1(n241_adj_4667), 
            .CO(n28905));
    SB_LUT4 add_5209_3_lut (.I0(GND_net), .I1(n9496[0]), .I2(n168_adj_4666), 
            .I3(n28903), .O(n9478[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5209_3 (.CI(n28903), .I0(n9496[0]), .I1(n168_adj_4666), 
            .CO(n28904));
    SB_LUT4 add_5209_2_lut (.I0(GND_net), .I1(n26_adj_4665), .I2(n95_adj_4664), 
            .I3(GND_net), .O(n9478[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5209_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5209_2 (.CI(GND_net), .I0(n26_adj_4665), .I1(n95_adj_4664), 
            .CO(n28903));
    SB_LUT4 add_5208_18_lut (.I0(GND_net), .I1(n9478[15]), .I2(GND_net), 
            .I3(n28902), .O(n9459[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5208_17_lut (.I0(GND_net), .I1(n9478[14]), .I2(GND_net), 
            .I3(n28901), .O(n9459[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4587));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5208_17 (.CI(n28901), .I0(n9478[14]), .I1(GND_net), .CO(n28902));
    SB_LUT4 add_5208_16_lut (.I0(GND_net), .I1(n9478[13]), .I2(n1114_adj_4662), 
            .I3(n28900), .O(n9459[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4586));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5208_16 (.CI(n28900), .I0(n9478[13]), .I1(n1114_adj_4662), 
            .CO(n28901));
    SB_LUT4 add_5208_15_lut (.I0(GND_net), .I1(n9478[12]), .I2(n1041_adj_4661), 
            .I3(n28899), .O(n9459[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_15 (.CI(n28899), .I0(n9478[12]), .I1(n1041_adj_4661), 
            .CO(n28900));
    SB_LUT4 add_5208_14_lut (.I0(GND_net), .I1(n9478[11]), .I2(n968_adj_4660), 
            .I3(n28898), .O(n9459[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_14 (.CI(n28898), .I0(n9478[11]), .I1(n968_adj_4660), 
            .CO(n28899));
    SB_LUT4 add_5208_13_lut (.I0(GND_net), .I1(n9478[10]), .I2(n895_adj_4659), 
            .I3(n28897), .O(n9459[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_13 (.CI(n28897), .I0(n9478[10]), .I1(n895_adj_4659), 
            .CO(n28898));
    SB_LUT4 add_5208_12_lut (.I0(GND_net), .I1(n9478[9]), .I2(n822_adj_4658), 
            .I3(n28896), .O(n9459[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_12 (.CI(n28896), .I0(n9478[9]), .I1(n822_adj_4658), 
            .CO(n28897));
    SB_LUT4 add_5208_11_lut (.I0(GND_net), .I1(n9478[8]), .I2(n749_adj_4657), 
            .I3(n28895), .O(n9459[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_11 (.CI(n28895), .I0(n9478[8]), .I1(n749_adj_4657), 
            .CO(n28896));
    SB_LUT4 add_5208_10_lut (.I0(GND_net), .I1(n9478[7]), .I2(n676_adj_4656), 
            .I3(n28894), .O(n9459[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_10 (.CI(n28894), .I0(n9478[7]), .I1(n676_adj_4656), 
            .CO(n28895));
    SB_LUT4 add_5208_9_lut (.I0(GND_net), .I1(n9478[6]), .I2(n603_adj_4655), 
            .I3(n28893), .O(n9459[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_9 (.CI(n28893), .I0(n9478[6]), .I1(n603_adj_4655), 
            .CO(n28894));
    SB_LUT4 add_5208_8_lut (.I0(GND_net), .I1(n9478[5]), .I2(n530_adj_4654), 
            .I3(n28892), .O(n9459[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_8 (.CI(n28892), .I0(n9478[5]), .I1(n530_adj_4654), 
            .CO(n28893));
    SB_LUT4 add_5208_7_lut (.I0(GND_net), .I1(n9478[4]), .I2(n457_adj_4653), 
            .I3(n28891), .O(n9459[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_7 (.CI(n28891), .I0(n9478[4]), .I1(n457_adj_4653), 
            .CO(n28892));
    SB_LUT4 add_5208_6_lut (.I0(GND_net), .I1(n9478[3]), .I2(n384_adj_4651), 
            .I3(n28890), .O(n9459[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_6 (.CI(n28890), .I0(n9478[3]), .I1(n384_adj_4651), 
            .CO(n28891));
    SB_LUT4 add_5208_5_lut (.I0(GND_net), .I1(n9478[2]), .I2(n311_adj_4650), 
            .I3(n28889), .O(n9459[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_5 (.CI(n28889), .I0(n9478[2]), .I1(n311_adj_4650), 
            .CO(n28890));
    SB_LUT4 add_5208_4_lut (.I0(GND_net), .I1(n9478[1]), .I2(n238_adj_4649), 
            .I3(n28888), .O(n9459[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[19]), 
            .I3(n27947), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_4 (.CI(n28888), .I0(n9478[1]), .I1(n238_adj_4649), 
            .CO(n28889));
    SB_LUT4 add_5208_3_lut (.I0(GND_net), .I1(n9478[0]), .I2(n165_adj_4643), 
            .I3(n28887), .O(n9459[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_3 (.CI(n28887), .I0(n9478[0]), .I1(n165_adj_4643), 
            .CO(n28888));
    SB_LUT4 add_5208_2_lut (.I0(GND_net), .I1(n23_adj_4642), .I2(n92_adj_4640), 
            .I3(GND_net), .O(n9459[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5208_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5208_2 (.CI(GND_net), .I0(n23_adj_4642), .I1(n92_adj_4640), 
            .CO(n28887));
    SB_LUT4 add_5207_19_lut (.I0(GND_net), .I1(n9459[16]), .I2(GND_net), 
            .I3(n28886), .O(n9439[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5207_18_lut (.I0(GND_net), .I1(n9459[15]), .I2(GND_net), 
            .I3(n28885), .O(n9439[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_18 (.CI(n28885), .I0(n9459[15]), .I1(GND_net), .CO(n28886));
    SB_LUT4 add_5207_17_lut (.I0(GND_net), .I1(n9459[14]), .I2(GND_net), 
            .I3(n28884), .O(n9439[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_17 (.CI(n28884), .I0(n9459[14]), .I1(GND_net), .CO(n28885));
    SB_LUT4 add_5207_16_lut (.I0(GND_net), .I1(n9459[13]), .I2(n1111_adj_4603), 
            .I3(n28883), .O(n9439[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_16 (.CI(n28883), .I0(n9459[13]), .I1(n1111_adj_4603), 
            .CO(n28884));
    SB_LUT4 add_5207_15_lut (.I0(GND_net), .I1(n9459[12]), .I2(n1038_adj_4600), 
            .I3(n28882), .O(n9439[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_15 (.CI(n28882), .I0(n9459[12]), .I1(n1038_adj_4600), 
            .CO(n28883));
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5207_14_lut (.I0(GND_net), .I1(n9459[11]), .I2(n965_adj_4597), 
            .I3(n28881), .O(n9439[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_14 (.CI(n28881), .I0(n9459[11]), .I1(n965_adj_4597), 
            .CO(n28882));
    SB_LUT4 add_5207_13_lut (.I0(GND_net), .I1(n9459[10]), .I2(n892_adj_4577), 
            .I3(n28880), .O(n9439[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_13 (.CI(n28880), .I0(n9459[10]), .I1(n892_adj_4577), 
            .CO(n28881));
    SB_LUT4 add_5207_12_lut (.I0(GND_net), .I1(n9459[9]), .I2(n819_adj_4573), 
            .I3(n28879), .O(n9439[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4584));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5207_12 (.CI(n28879), .I0(n9459[9]), .I1(n819_adj_4573), 
            .CO(n28880));
    SB_LUT4 add_5207_11_lut (.I0(GND_net), .I1(n9459[8]), .I2(n746_adj_4571), 
            .I3(n28878), .O(n9439[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_11 (.CI(n28878), .I0(n9459[8]), .I1(n746_adj_4571), 
            .CO(n28879));
    SB_LUT4 add_5207_10_lut (.I0(GND_net), .I1(n9459[7]), .I2(n673), .I3(n28877), 
            .O(n9439[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_10 (.CI(n28877), .I0(n9459[7]), .I1(n673), .CO(n28878));
    SB_LUT4 add_5207_9_lut (.I0(GND_net), .I1(n9459[6]), .I2(n600), .I3(n28876), 
            .O(n9439[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_9 (.CI(n28876), .I0(n9459[6]), .I1(n600), .CO(n28877));
    SB_LUT4 add_5207_8_lut (.I0(GND_net), .I1(n9459[5]), .I2(n527), .I3(n28875), 
            .O(n9439[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_8 (.CI(n28875), .I0(n9459[5]), .I1(n527), .CO(n28876));
    SB_LUT4 add_5207_7_lut (.I0(GND_net), .I1(n9459[4]), .I2(n454), .I3(n28874), 
            .O(n9439[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_7 (.CI(n28874), .I0(n9459[4]), .I1(n454), .CO(n28875));
    SB_LUT4 add_5207_6_lut (.I0(GND_net), .I1(n9459[3]), .I2(n381), .I3(n28873), 
            .O(n9439[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_6 (.CI(n28873), .I0(n9459[3]), .I1(n381), .CO(n28874));
    SB_LUT4 add_5207_5_lut (.I0(GND_net), .I1(n9459[2]), .I2(n308), .I3(n28872), 
            .O(n9439[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_5 (.CI(n28872), .I0(n9459[2]), .I1(n308), .CO(n28873));
    SB_LUT4 add_5207_4_lut (.I0(GND_net), .I1(n9459[1]), .I2(n235), .I3(n28871), 
            .O(n9439[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_4 (.CI(n28871), .I0(n9459[1]), .I1(n235), .CO(n28872));
    SB_LUT4 add_5207_3_lut (.I0(GND_net), .I1(n9459[0]), .I2(n162), .I3(n28870), 
            .O(n9439[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_3 (.CI(n28870), .I0(n9459[0]), .I1(n162), .CO(n28871));
    SB_LUT4 add_5207_2_lut (.I0(GND_net), .I1(n20_adj_4560), .I2(n89), 
            .I3(GND_net), .O(n9439[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5207_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5207_2 (.CI(GND_net), .I0(n20_adj_4560), .I1(n89), .CO(n28870));
    SB_LUT4 add_5206_20_lut (.I0(GND_net), .I1(n9439[17]), .I2(GND_net), 
            .I3(n28869), .O(n9418[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5206_19_lut (.I0(GND_net), .I1(n9439[16]), .I2(GND_net), 
            .I3(n28868), .O(n9418[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_19 (.CI(n28868), .I0(n9439[16]), .I1(GND_net), .CO(n28869));
    SB_LUT4 add_5206_18_lut (.I0(GND_net), .I1(n9439[15]), .I2(GND_net), 
            .I3(n28867), .O(n9418[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_18 (.CI(n28867), .I0(n9439[15]), .I1(GND_net), .CO(n28868));
    SB_LUT4 add_5206_17_lut (.I0(GND_net), .I1(n9439[14]), .I2(GND_net), 
            .I3(n28866), .O(n9418[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_17 (.CI(n28866), .I0(n9439[14]), .I1(GND_net), .CO(n28867));
    SB_LUT4 add_5206_16_lut (.I0(GND_net), .I1(n9439[13]), .I2(n1108), 
            .I3(n28865), .O(n9418[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_16 (.CI(n28865), .I0(n9439[13]), .I1(n1108), .CO(n28866));
    SB_LUT4 add_5206_15_lut (.I0(GND_net), .I1(n9439[12]), .I2(n1035), 
            .I3(n28864), .O(n9418[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_15 (.CI(n28864), .I0(n9439[12]), .I1(n1035), .CO(n28865));
    SB_LUT4 add_5206_14_lut (.I0(GND_net), .I1(n9439[11]), .I2(n962), 
            .I3(n28863), .O(n9418[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_14 (.CI(n28863), .I0(n9439[11]), .I1(n962), .CO(n28864));
    SB_LUT4 add_5206_13_lut (.I0(GND_net), .I1(n9439[10]), .I2(n889), 
            .I3(n28862), .O(n9418[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_13 (.CI(n28862), .I0(n9439[10]), .I1(n889), .CO(n28863));
    SB_LUT4 add_5206_12_lut (.I0(GND_net), .I1(n9439[9]), .I2(n816), .I3(n28861), 
            .O(n9418[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_12 (.CI(n28861), .I0(n9439[9]), .I1(n816), .CO(n28862));
    SB_LUT4 add_5206_11_lut (.I0(GND_net), .I1(n9439[8]), .I2(n743), .I3(n28860), 
            .O(n9418[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_11 (.CI(n28860), .I0(n9439[8]), .I1(n743), .CO(n28861));
    SB_LUT4 add_5206_10_lut (.I0(GND_net), .I1(n9439[7]), .I2(n670), .I3(n28859), 
            .O(n9418[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_10 (.CI(n28859), .I0(n9439[7]), .I1(n670), .CO(n28860));
    SB_LUT4 add_5206_9_lut (.I0(GND_net), .I1(n9439[6]), .I2(n597), .I3(n28858), 
            .O(n9418[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_9 (.CI(n28858), .I0(n9439[6]), .I1(n597), .CO(n28859));
    SB_LUT4 add_5206_8_lut (.I0(GND_net), .I1(n9439[5]), .I2(n524), .I3(n28857), 
            .O(n9418[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_8 (.CI(n28857), .I0(n9439[5]), .I1(n524), .CO(n28858));
    SB_LUT4 add_5206_7_lut (.I0(GND_net), .I1(n9439[4]), .I2(n451), .I3(n28856), 
            .O(n9418[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_7 (.CI(n28856), .I0(n9439[4]), .I1(n451), .CO(n28857));
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4583));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5206_6_lut (.I0(GND_net), .I1(n9439[3]), .I2(n378), .I3(n28855), 
            .O(n9418[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_6 (.CI(n28855), .I0(n9439[3]), .I1(n378), .CO(n28856));
    SB_LUT4 add_5206_5_lut (.I0(GND_net), .I1(n9439[2]), .I2(n305), .I3(n28854), 
            .O(n9418[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_5 (.CI(n28854), .I0(n9439[2]), .I1(n305), .CO(n28855));
    SB_LUT4 add_5206_4_lut (.I0(GND_net), .I1(n9439[1]), .I2(n232), .I3(n28853), 
            .O(n9418[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_4 (.CI(n28853), .I0(n9439[1]), .I1(n232), .CO(n28854));
    SB_LUT4 add_5206_3_lut (.I0(GND_net), .I1(n9439[0]), .I2(n159), .I3(n28852), 
            .O(n9418[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_3 (.CI(n28852), .I0(n9439[0]), .I1(n159), .CO(n28853));
    SB_LUT4 add_5206_2_lut (.I0(GND_net), .I1(n17_adj_4502), .I2(n86), 
            .I3(GND_net), .O(n9418[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5206_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5206_2 (.CI(GND_net), .I0(n17_adj_4502), .I1(n86), .CO(n28852));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n27947), .I0(GND_net), .I1(n1_adj_4708[19]), 
            .CO(n27948));
    SB_LUT4 add_5205_21_lut (.I0(GND_net), .I1(n9418[18]), .I2(GND_net), 
            .I3(n28851), .O(n9396[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5205_20_lut (.I0(GND_net), .I1(n9418[17]), .I2(GND_net), 
            .I3(n28850), .O(n9396[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_20 (.CI(n28850), .I0(n9418[17]), .I1(GND_net), .CO(n28851));
    SB_LUT4 add_739_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n3223[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3509 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_739_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4582));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5205_19_lut (.I0(GND_net), .I1(n9418[16]), .I2(GND_net), 
            .I3(n28849), .O(n9396[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_19 (.CI(n28849), .I0(n9418[16]), .I1(GND_net), .CO(n28850));
    SB_LUT4 add_5205_18_lut (.I0(GND_net), .I1(n9418[15]), .I2(GND_net), 
            .I3(n28848), .O(n9396[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_18 (.CI(n28848), .I0(n9418[15]), .I1(GND_net), .CO(n28849));
    SB_LUT4 add_5205_17_lut (.I0(GND_net), .I1(n9418[14]), .I2(GND_net), 
            .I3(n28847), .O(n9396[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_17 (.CI(n28847), .I0(n9418[14]), .I1(GND_net), .CO(n28848));
    SB_LUT4 add_5205_16_lut (.I0(GND_net), .I1(n9418[13]), .I2(n1105), 
            .I3(n28846), .O(n9396[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_16 (.CI(n28846), .I0(n9418[13]), .I1(n1105), .CO(n28847));
    SB_LUT4 add_5205_15_lut (.I0(GND_net), .I1(n9418[12]), .I2(n1032), 
            .I3(n28845), .O(n9396[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_15 (.CI(n28845), .I0(n9418[12]), .I1(n1032), .CO(n28846));
    SB_LUT4 add_5205_14_lut (.I0(GND_net), .I1(n9418[11]), .I2(n959), 
            .I3(n28844), .O(n9396[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_14 (.CI(n28844), .I0(n9418[11]), .I1(n959), .CO(n28845));
    SB_LUT4 add_5205_13_lut (.I0(GND_net), .I1(n9418[10]), .I2(n886), 
            .I3(n28843), .O(n9396[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_13 (.CI(n28843), .I0(n9418[10]), .I1(n886), .CO(n28844));
    SB_LUT4 add_5205_12_lut (.I0(GND_net), .I1(n9418[9]), .I2(n813), .I3(n28842), 
            .O(n9396[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_12 (.CI(n28842), .I0(n9418[9]), .I1(n813), .CO(n28843));
    SB_LUT4 add_5205_11_lut (.I0(GND_net), .I1(n9418[8]), .I2(n740), .I3(n28841), 
            .O(n9396[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4581));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5205_11 (.CI(n28841), .I0(n9418[8]), .I1(n740), .CO(n28842));
    SB_LUT4 add_5205_10_lut (.I0(GND_net), .I1(n9418[7]), .I2(n667), .I3(n28840), 
            .O(n9396[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_10 (.CI(n28840), .I0(n9418[7]), .I1(n667), .CO(n28841));
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4580));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5205_9_lut (.I0(GND_net), .I1(n9418[6]), .I2(n594), .I3(n28839), 
            .O(n9396[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_9 (.CI(n28839), .I0(n9418[6]), .I1(n594), .CO(n28840));
    SB_LUT4 add_5205_8_lut (.I0(GND_net), .I1(n9418[5]), .I2(n521), .I3(n28838), 
            .O(n9396[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_8 (.CI(n28838), .I0(n9418[5]), .I1(n521), .CO(n28839));
    SB_LUT4 add_5205_7_lut (.I0(GND_net), .I1(n9418[4]), .I2(n448), .I3(n28837), 
            .O(n9396[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_7 (.CI(n28837), .I0(n9418[4]), .I1(n448), .CO(n28838));
    SB_LUT4 add_5205_6_lut (.I0(GND_net), .I1(n9418[3]), .I2(n375), .I3(n28836), 
            .O(n9396[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_6 (.CI(n28836), .I0(n9418[3]), .I1(n375), .CO(n28837));
    SB_LUT4 add_5205_5_lut (.I0(GND_net), .I1(n9418[2]), .I2(n302), .I3(n28835), 
            .O(n9396[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_5 (.CI(n28835), .I0(n9418[2]), .I1(n302), .CO(n28836));
    SB_LUT4 add_5205_4_lut (.I0(GND_net), .I1(n9418[1]), .I2(n229), .I3(n28834), 
            .O(n9396[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_4 (.CI(n28834), .I0(n9418[1]), .I1(n229), .CO(n28835));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[18]), 
            .I3(n27946), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5205_3_lut (.I0(GND_net), .I1(n9418[0]), .I2(n156), .I3(n28833), 
            .O(n9396[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_3 (.CI(n28833), .I0(n9418[0]), .I1(n156), .CO(n28834));
    SB_LUT4 add_5205_2_lut (.I0(GND_net), .I1(n14_adj_4438), .I2(n83), 
            .I3(GND_net), .O(n9396[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5205_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5205_2 (.CI(GND_net), .I0(n14_adj_4438), .I1(n83), .CO(n28833));
    SB_LUT4 add_5204_22_lut (.I0(GND_net), .I1(n9396[19]), .I2(GND_net), 
            .I3(n28832), .O(n9373[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5204_21_lut (.I0(GND_net), .I1(n9396[18]), .I2(GND_net), 
            .I3(n28831), .O(n9373[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_21 (.CI(n28831), .I0(n9396[18]), .I1(GND_net), .CO(n28832));
    SB_LUT4 add_5204_20_lut (.I0(GND_net), .I1(n9396[17]), .I2(GND_net), 
            .I3(n28830), .O(n9373[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_20 (.CI(n28830), .I0(n9396[17]), .I1(GND_net), .CO(n28831));
    SB_LUT4 add_5204_19_lut (.I0(GND_net), .I1(n9396[16]), .I2(GND_net), 
            .I3(n28829), .O(n9373[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4579));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4578));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5204_19 (.CI(n28829), .I0(n9396[16]), .I1(GND_net), .CO(n28830));
    SB_LUT4 add_5204_18_lut (.I0(GND_net), .I1(n9396[15]), .I2(GND_net), 
            .I3(n28828), .O(n9373[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_18 (.CI(n28828), .I0(n9396[15]), .I1(GND_net), .CO(n28829));
    SB_LUT4 add_5204_17_lut (.I0(GND_net), .I1(n9396[14]), .I2(GND_net), 
            .I3(n28827), .O(n9373[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_17 (.CI(n28827), .I0(n9396[14]), .I1(GND_net), .CO(n28828));
    SB_LUT4 add_5204_16_lut (.I0(GND_net), .I1(n9396[13]), .I2(n1102), 
            .I3(n28826), .O(n9373[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_16 (.CI(n28826), .I0(n9396[13]), .I1(n1102), .CO(n28827));
    SB_LUT4 add_5204_15_lut (.I0(GND_net), .I1(n9396[12]), .I2(n1029), 
            .I3(n28825), .O(n9373[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_15 (.CI(n28825), .I0(n9396[12]), .I1(n1029), .CO(n28826));
    SB_LUT4 add_5204_14_lut (.I0(GND_net), .I1(n9396[11]), .I2(n956), 
            .I3(n28824), .O(n9373[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_14 (.CI(n28824), .I0(n9396[11]), .I1(n956), .CO(n28825));
    SB_LUT4 add_5204_13_lut (.I0(GND_net), .I1(n9396[10]), .I2(n883), 
            .I3(n28823), .O(n9373[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_13 (.CI(n28823), .I0(n9396[10]), .I1(n883), .CO(n28824));
    SB_LUT4 add_5204_12_lut (.I0(GND_net), .I1(n9396[9]), .I2(n810), .I3(n28822), 
            .O(n9373[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_12 (.CI(n28822), .I0(n9396[9]), .I1(n810), .CO(n28823));
    SB_LUT4 add_5204_11_lut (.I0(GND_net), .I1(n9396[8]), .I2(n737), .I3(n28821), 
            .O(n9373[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_11 (.CI(n28821), .I0(n9396[8]), .I1(n737), .CO(n28822));
    SB_LUT4 add_5204_10_lut (.I0(GND_net), .I1(n9396[7]), .I2(n664), .I3(n28820), 
            .O(n9373[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_10 (.CI(n28820), .I0(n9396[7]), .I1(n664), .CO(n28821));
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4576));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5204_9_lut (.I0(GND_net), .I1(n9396[6]), .I2(n591), .I3(n28819), 
            .O(n9373[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_9 (.CI(n28819), .I0(n9396[6]), .I1(n591), .CO(n28820));
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4706));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5204_8_lut (.I0(GND_net), .I1(n9396[5]), .I2(n518), .I3(n28818), 
            .O(n9373[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_8 (.CI(n28818), .I0(n9396[5]), .I1(n518), .CO(n28819));
    SB_LUT4 add_5204_7_lut (.I0(GND_net), .I1(n9396[4]), .I2(n445), .I3(n28817), 
            .O(n9373[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4575));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5204_7 (.CI(n28817), .I0(n9396[4]), .I1(n445), .CO(n28818));
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4574));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5204_6_lut (.I0(GND_net), .I1(n9396[3]), .I2(n372), .I3(n28816), 
            .O(n9373[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_6 (.CI(n28816), .I0(n9396[3]), .I1(n372), .CO(n28817));
    SB_LUT4 add_5204_5_lut (.I0(GND_net), .I1(n9396[2]), .I2(n299), .I3(n28815), 
            .O(n9373[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_5 (.CI(n28815), .I0(n9396[2]), .I1(n299), .CO(n28816));
    SB_LUT4 add_5204_4_lut (.I0(GND_net), .I1(n9396[1]), .I2(n226), .I3(n28814), 
            .O(n9373[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_739_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n3223[0]), .CO(n27800));
    SB_CARRY add_5204_4 (.CI(n28814), .I0(n9396[1]), .I1(n226), .CO(n28815));
    SB_LUT4 add_5204_3_lut (.I0(GND_net), .I1(n9396[0]), .I2(n153), .I3(n28813), 
            .O(n9373[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_3 (.CI(n28813), .I0(n9396[0]), .I1(n153), .CO(n28814));
    SB_LUT4 add_5204_2_lut (.I0(GND_net), .I1(n11_adj_4433), .I2(n80), 
            .I3(GND_net), .O(n9373[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5204_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5204_2 (.CI(GND_net), .I0(n11_adj_4433), .I1(n80), .CO(n28813));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n28[23]), .I1(n9349[21]), .I2(GND_net), 
            .I3(n28812), .O(n8060[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n9349[20]), .I2(GND_net), 
            .I3(n28811), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n28811), .I0(n9349[20]), .I1(GND_net), 
            .CO(n28812));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n9349[19]), .I2(GND_net), 
            .I3(n28810), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n28810), .I0(n9349[19]), .I1(GND_net), 
            .CO(n28811));
    SB_CARRY unary_minus_16_add_3_20 (.CI(n27946), .I0(GND_net), .I1(n1_adj_4708[18]), 
            .CO(n27947));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n9349[18]), .I2(GND_net), 
            .I3(n28809), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n28809), .I0(n9349[18]), .I1(GND_net), 
            .CO(n28810));
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4705));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n9349[17]), .I2(GND_net), 
            .I3(n28808), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_20 (.CI(n28808), .I0(n9349[17]), .I1(GND_net), 
            .CO(n28809));
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4572));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n9349[16]), .I2(GND_net), 
            .I3(n28807), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n28807), .I0(n9349[16]), .I1(GND_net), 
            .CO(n28808));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n9349[15]), .I2(GND_net), 
            .I3(n28806), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n28806), .I0(n9349[15]), .I1(GND_net), 
            .CO(n28807));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n9349[14]), .I2(GND_net), 
            .I3(n28805), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n28805), .I0(n9349[14]), .I1(GND_net), 
            .CO(n28806));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n9349[13]), .I2(n1096), 
            .I3(n28804), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n28804), .I0(n9349[13]), .I1(n1096), 
            .CO(n28805));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n9349[12]), .I2(n1023), 
            .I3(n28803), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n28803), .I0(n9349[12]), .I1(n1023), 
            .CO(n28804));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n9349[11]), .I2(n950), 
            .I3(n28802), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n28802), .I0(n9349[11]), .I1(n950), 
            .CO(n28803));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n9349[10]), .I2(n877), 
            .I3(n28801), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n28801), .I0(n9349[10]), .I1(n877), 
            .CO(n28802));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n9349[9]), .I2(n804), 
            .I3(n28800), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n28800), .I0(n9349[9]), .I1(n804), 
            .CO(n28801));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n9349[8]), .I2(n731), 
            .I3(n28799), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n28799), .I0(n9349[8]), .I1(n731), 
            .CO(n28800));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n9349[7]), .I2(n658), 
            .I3(n28798), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n28798), .I0(n9349[7]), .I1(n658), 
            .CO(n28799));
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4704));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n9349[6]), .I2(n585), 
            .I3(n28797), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n28797), .I0(n9349[6]), .I1(n585), 
            .CO(n28798));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n9349[5]), .I2(n512), 
            .I3(n28796), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_8 (.CI(n28796), .I0(n9349[5]), .I1(n512), 
            .CO(n28797));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n9349[4]), .I2(n439), 
            .I3(n28795), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n28795), .I0(n9349[4]), .I1(n439), 
            .CO(n28796));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[17]), 
            .I3(n27945), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n9349[3]), .I2(n366), 
            .I3(n28794), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n28794), .I0(n9349[3]), .I1(n366), 
            .CO(n28795));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n9349[2]), .I2(n293), 
            .I3(n28793), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n28793), .I0(n9349[2]), .I1(n293), 
            .CO(n28794));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n9349[1]), .I2(n220), 
            .I3(n28792), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n28792), .I0(n9349[1]), .I1(n220), 
            .CO(n28793));
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4703));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n9349[0]), .I2(n147), 
            .I3(n28791), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4702));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4701));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n27945), .I0(GND_net), .I1(n1_adj_4708[17]), 
            .CO(n27946));
    SB_CARRY mult_10_add_1225_3 (.CI(n28791), .I0(n9349[0]), .I1(n147), 
            .CO(n28792));
    SB_CARRY add_12_3 (.CI(n27757), .I0(n106[1]), .I1(n155[1]), .CO(n27758));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4413), .I2(n74), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4413), .I1(n74), 
            .CO(n28791));
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3609[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22716_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[20]), .I2(n27450), 
            .I3(n9639[0]), .O(n4_adj_4391));   // verilog/motorControl.v(34[16:22])
    defparam i22716_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4699));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4698));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1509 (.I0(\Kp[2] ), .I1(n28[20]), .I2(n9639[0]), 
            .I3(n27450), .O(n9634[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1509.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[16]), 
            .I3(n27944), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5203_23_lut (.I0(GND_net), .I1(n9373[20]), .I2(GND_net), 
            .I3(n28790), .O(n9349[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5203_22_lut (.I0(GND_net), .I1(n9373[19]), .I2(GND_net), 
            .I3(n28789), .O(n9349[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n27757));
    SB_CARRY add_5203_22 (.CI(n28789), .I0(n9373[19]), .I1(GND_net), .CO(n28790));
    SB_LUT4 i22703_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n9634[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22703_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_5203_21_lut (.I0(GND_net), .I1(n9373[18]), .I2(GND_net), 
            .I3(n28788), .O(n9349[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_21 (.CI(n28788), .I0(n9373[18]), .I1(GND_net), .CO(n28789));
    SB_LUT4 add_5203_20_lut (.I0(GND_net), .I1(n9373[17]), .I2(GND_net), 
            .I3(n28787), .O(n9349[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_20 (.CI(n28787), .I0(n9373[17]), .I1(GND_net), .CO(n28788));
    SB_LUT4 add_5203_19_lut (.I0(GND_net), .I1(n9373[16]), .I2(GND_net), 
            .I3(n28786), .O(n9349[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_19 (.CI(n28786), .I0(n9373[16]), .I1(GND_net), .CO(n28787));
    SB_LUT4 add_5203_18_lut (.I0(GND_net), .I1(n9373[15]), .I2(GND_net), 
            .I3(n28785), .O(n9349[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22705_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n27450));   // verilog/motorControl.v(34[16:22])
    defparam i22705_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n27944), .I0(GND_net), .I1(n1_adj_4708[16]), 
            .CO(n27945));
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4696));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463_adj_4695));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4693));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5203_18 (.CI(n28785), .I0(n9373[15]), .I1(GND_net), .CO(n28786));
    SB_LUT4 add_5203_17_lut (.I0(GND_net), .I1(n9373[14]), .I2(GND_net), 
            .I3(n28784), .O(n9349[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[15]), 
            .I3(n27943), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_17 (.CI(n28784), .I0(n9373[14]), .I1(GND_net), .CO(n28785));
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5203_16_lut (.I0(GND_net), .I1(n9373[13]), .I2(n1099), 
            .I3(n28783), .O(n9349[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_16 (.CI(n28783), .I0(n9373[13]), .I1(n1099), .CO(n28784));
    SB_LUT4 add_5203_15_lut (.I0(GND_net), .I1(n9373[12]), .I2(n1026), 
            .I3(n28782), .O(n9349[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_15 (.CI(n28782), .I0(n9373[12]), .I1(n1026), .CO(n28783));
    SB_LUT4 add_5203_14_lut (.I0(GND_net), .I1(n9373[11]), .I2(n953), 
            .I3(n28781), .O(n9349[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n27943), .I0(GND_net), .I1(n1_adj_4708[15]), 
            .CO(n27944));
    SB_CARRY add_5203_14 (.CI(n28781), .I0(n9373[11]), .I1(n953), .CO(n28782));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4708[14]), 
            .I3(n27942), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5203_13_lut (.I0(GND_net), .I1(n9373[10]), .I2(n880), 
            .I3(n28780), .O(n9349[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_13 (.CI(n28780), .I0(n9373[10]), .I1(n880), .CO(n28781));
    SB_LUT4 add_5203_12_lut (.I0(GND_net), .I1(n9373[9]), .I2(n807), .I3(n28779), 
            .O(n9349[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5203_12 (.CI(n28779), .I0(n9373[9]), .I1(n807), .CO(n28780));
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5203_11_lut (.I0(GND_net), .I1(n9373[8]), .I2(n734), .I3(n28778), 
            .O(n9349[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5203_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4565));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4692));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22685_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[19]), .I2(n27416), 
            .I3(n9634[0]), .O(n4_adj_4380));   // verilog/motorControl.v(34[16:22])
    defparam i22685_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4690));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4689));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19378_2_lut (.I0(n28[2]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19378_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19379_2_lut (.I0(n28[3]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19379_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1510 (.I0(\Kp[2] ), .I1(n28[19]), .I2(n9634[0]), 
            .I3(n27416), .O(n9628[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1510.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4708[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22672_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(n28[19]), 
            .I3(\Kp[1] ), .O(n9628[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22672_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i22674_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(n28[19]), 
            .I3(\Kp[1] ), .O(n27416));   // verilog/motorControl.v(34[16:22])
    defparam i22674_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4561));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4684));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19380_2_lut (.I0(n28[4]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19380_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22654_3_lut_4_lut (.I0(\Kp[3] ), .I1(n28[18]), .I2(n4_adj_4707), 
            .I3(n9628[1]), .O(n6_adj_4377));   // verilog/motorControl.v(34[16:22])
    defparam i22654_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1511 (.I0(\Kp[3] ), .I1(n28[18]), .I2(n9628[1]), 
            .I3(n4_adj_4707), .O(n9621[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1511.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1512 (.I0(\Kp[2] ), .I1(n28[18]), .I2(n9628[0]), 
            .I3(n27373), .O(n9621[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1512.LUT_INIT = 16'h8778;
    SB_LUT4 i22646_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[18]), .I2(n27373), 
            .I3(n9628[0]), .O(n4_adj_4707));   // verilog/motorControl.v(34[16:22])
    defparam i22646_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i22633_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n9621[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22633_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22635_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n27373));   // verilog/motorControl.v(34[16:22])
    defparam i22635_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4552));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4683));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19381_2_lut (.I0(n28[5]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19381_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4680));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19382_2_lut (.I0(n28[6]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19382_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19383_2_lut (.I0(n28[7]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19383_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4678));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19384_2_lut (.I0(n28[8]), .I1(\PID_CONTROLLER.integral_23__N_3557 ), 
            .I2(GND_net), .I3(GND_net), .O(n3223[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19384_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4550));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4549));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4677));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4547));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4546));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4544));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4543));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4538));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4537));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4535));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4534));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4531));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4528));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4525));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4522));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4520));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4519));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4517));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4516));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4514));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4513));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4512));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4511));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3509 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4510));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (CLK_c, GND_net, \state[3] , n6, n3567, \state[1] , 
            \state[0] , enable_slow_N_3964, n33160, n32413, read, 
            n23704, \state[2] , n7, n18643, rw, n32166, data_ready, 
            n32068, n32064, n10, n17058, n17053, n4867, \saved_addr[0] , 
            \state[0]_adj_13 , \state_7__N_3861[0] , n4, n35900, n4_adj_14, 
            scl_enable, sda_enable, \state_7__N_3877[3] , VCC_net, scl, 
            sda_out, n10_adj_15, n5300, n8, n18652, data, n18650, 
            n18649, n18648, n18647, n18646, n19174, n23726, n18633, 
            n18632) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    input GND_net;
    output \state[3] ;
    output n6;
    output [0:0]n3567;
    output \state[1] ;
    output \state[0] ;
    output enable_slow_N_3964;
    input n33160;
    output n32413;
    input read;
    output n23704;
    output \state[2] ;
    output n7;
    input n18643;
    output rw;
    input n32166;
    output data_ready;
    input n32068;
    input n32064;
    output n10;
    output n17058;
    output n17053;
    output n4867;
    output \saved_addr[0] ;
    output \state[0]_adj_13 ;
    output \state_7__N_3861[0] ;
    output n4;
    output n35900;
    output n4_adj_14;
    output scl_enable;
    output sda_enable;
    input \state_7__N_3877[3] ;
    input VCC_net;
    output scl;
    output sda_out;
    output n10_adj_15;
    input n5300;
    input n8;
    input n18652;
    output [7:0]data;
    input n18650;
    input n18649;
    input n18648;
    input n18647;
    input n18646;
    input n19174;
    output n23726;
    input n18633;
    input n18632;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3763;
    
    wire n18317;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n18558, n27798;
    wire [15:0]n3259;
    
    wire n27799, n27797, n16909, n27796, enable, n27795, n27794, 
        n27793, n27792, n27791, n27790, n27789, n27788, n27787, 
        n27786, n27785;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n28, n26, n27, n25;
    
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[15]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[12]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[11]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[10]), .S(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[9]), .S(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[8]), .S(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[7]), .S(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[6]), .S(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[5]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[4]), .S(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[3]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[2]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[1]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_CARRY add_743_16 (.CI(n27798), .I0(delay_counter[14]), .I1(n3259[14]), 
            .CO(n27799));
    SB_LUT4 add_743_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n3259[14]), 
            .I3(n27797), .O(delay_counter_15__N_3763[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_15 (.CI(n27797), .I0(delay_counter[13]), .I1(n3259[14]), 
            .CO(n27798));
    SB_LUT4 i2_2_lut (.I0(\state[3] ), .I1(n16909), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_743_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n3259[14]), 
            .I3(n27796), .O(delay_counter_15__N_3763[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_14 (.CI(n27796), .I0(delay_counter[12]), .I1(n3259[14]), 
            .CO(n27797));
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[14]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n3567[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_743_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n3259[14]), 
            .I3(n27795), .O(delay_counter_15__N_3763[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_13 (.CI(n27795), .I0(delay_counter[11]), .I1(n3259[14]), 
            .CO(n27796));
    SB_LUT4 add_743_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n3259[14]), 
            .I3(n27794), .O(delay_counter_15__N_3763[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_12 (.CI(n27794), .I0(delay_counter[10]), .I1(n3259[14]), 
            .CO(n27795));
    SB_LUT4 add_743_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n3259[14]), 
            .I3(n27793), .O(delay_counter_15__N_3763[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_11_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[13]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_CARRY add_743_11 (.CI(n27793), .I0(delay_counter[9]), .I1(n3259[14]), 
            .CO(n27794));
    SB_LUT4 add_743_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n3259[14]), 
            .I3(n27792), .O(delay_counter_15__N_3763[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_10 (.CI(n27792), .I0(delay_counter[8]), .I1(n3259[14]), 
            .CO(n27793));
    SB_LUT4 add_743_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n3259[14]), 
            .I3(n27791), .O(delay_counter_15__N_3763[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_9 (.CI(n27791), .I0(delay_counter[7]), .I1(n3259[14]), 
            .CO(n27792));
    SB_LUT4 add_743_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n3259[14]), 
            .I3(n27790), .O(delay_counter_15__N_3763[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_8 (.CI(n27790), .I0(delay_counter[6]), .I1(n3259[14]), 
            .CO(n27791));
    SB_LUT4 add_743_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n3259[14]), 
            .I3(n27789), .O(delay_counter_15__N_3763[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_7 (.CI(n27789), .I0(delay_counter[5]), .I1(n3259[14]), 
            .CO(n27790));
    SB_LUT4 add_743_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n3259[14]), 
            .I3(n27788), .O(delay_counter_15__N_3763[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_6 (.CI(n27788), .I0(delay_counter[4]), .I1(n3259[14]), 
            .CO(n27789));
    SB_LUT4 add_743_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n3259[14]), 
            .I3(n27787), .O(delay_counter_15__N_3763[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_5 (.CI(n27787), .I0(delay_counter[3]), .I1(n3259[14]), 
            .CO(n27788));
    SB_LUT4 add_743_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n3259[14]), 
            .I3(n27786), .O(delay_counter_15__N_3763[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_4 (.CI(n27786), .I0(delay_counter[2]), .I1(n3259[14]), 
            .CO(n27787));
    SB_LUT4 i13782_2_lut (.I0(n18317), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n18558));   // verilog/eeprom.v(26[8] 58[4])
    defparam i13782_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_3964), 
            .I3(n33160), .O(n32413));   // verilog/eeprom.v(51[5:9])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n18317));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i19099_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_3964), 
            .I3(GND_net), .O(n23704));   // verilog/eeprom.v(51[5:9])
    defparam i19099_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 add_743_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n3259[14]), 
            .I3(n27785), .O(delay_counter_15__N_3763[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_3 (.CI(n27785), .I0(delay_counter[1]), .I1(n3259[14]), 
            .CO(n27786));
    SB_LUT4 add_743_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n3259[14]), 
            .I3(GND_net), .O(delay_counter_15__N_3763[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_743_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n3259[14]), 
            .CO(n27785));
    SB_LUT4 mux_925_Mux_0_i1_4_lut (.I0(read), .I1(n16909), .I2(\state[0] ), 
            .I3(enable_slow_N_3964), .O(n3567[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_925_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i2_2_lut_adj_1496 (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut_adj_1496.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n16909));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30438_2_lut (.I0(n16909), .I1(enable_slow_N_3964), .I2(GND_net), 
            .I3(GND_net), .O(n3259[14]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i30438_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n18317), 
            .D(delay_counter_15__N_3763[0]), .R(n18558));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n18643));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n32166));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n32068));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n32064));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_743_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n3259[14]), 
            .I3(n27799), .O(delay_counter_15__N_3763[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_743_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n3259[14]), 
            .I3(n27798), .O(delay_counter_15__N_3763[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_743_16_lut.LUT_INIT = 16'hC33C;
    i2c_controller i2c (.CLK_c(CLK_c), .n10(n10), .n17058(n17058), .GND_net(GND_net), 
            .n17053(n17053), .n4867(n4867), .\saved_addr[0] (\saved_addr[0] ), 
            .\state[1] (state[1]), .\state[2] (\state[2] ), .\state[0] (\state[0]_adj_13 ), 
            .\state[3] (\state[3] ), .\state_7__N_3861[0] (\state_7__N_3861[0] ), 
            .enable_slow_N_3964(enable_slow_N_3964), .n4(n4), .n35900(n35900), 
            .n4_adj_11(n4_adj_14), .scl_enable(scl_enable), .sda_enable(sda_enable), 
            .\state_7__N_3877[3] (\state_7__N_3877[3] ), .VCC_net(VCC_net), 
            .scl(scl), .enable(enable), .sda_out(sda_out), .n10_adj_12(n10_adj_15), 
            .n5300(n5300), .n8(n8), .n18652(n18652), .data({data}), 
            .n18650(n18650), .n18649(n18649), .n18648(n18648), .n18647(n18647), 
            .n18646(n18646), .n19174(n19174), .n23726(n23726), .n18633(n18633), 
            .n18632(n18632)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (CLK_c, n10, n17058, GND_net, n17053, n4867, 
            \saved_addr[0] , \state[1] , \state[2] , \state[0] , \state[3] , 
            \state_7__N_3861[0] , enable_slow_N_3964, n4, n35900, n4_adj_11, 
            scl_enable, sda_enable, \state_7__N_3877[3] , VCC_net, scl, 
            enable, sda_out, n10_adj_12, n5300, n8, n18652, data, 
            n18650, n18649, n18648, n18647, n18646, n19174, n23726, 
            n18633, n18632) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    output n10;
    output n17058;
    input GND_net;
    output n17053;
    output n4867;
    output \saved_addr[0] ;
    output \state[1] ;
    output \state[2] ;
    output \state[0] ;
    output \state[3] ;
    output \state_7__N_3861[0] ;
    output enable_slow_N_3964;
    output n4;
    output n35900;
    output n4_adj_11;
    output scl_enable;
    output sda_enable;
    input \state_7__N_3877[3] ;
    input VCC_net;
    output scl;
    input enable;
    output sda_out;
    output n10_adj_12;
    input n5300;
    input n8;
    input n18652;
    output [7:0]data;
    input n18650;
    input n18649;
    input n18648;
    input n18647;
    input n18646;
    input n19174;
    output n23726;
    input n18633;
    input n18632;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n18552;
    wire [7:0]n119;
    
    wire n18362;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n18604, n9, n11, n24174, n35961, n35877, n11_adj_4270, 
        n35980, n7, n33, n37, n18487, n34, n39, enable_slow_N_3963, 
        i2c_clk_N_3950, n32132, n11_adj_4271, n15, n24476, scl_enable_N_3951, 
        n18254, n10190, n5184, sda_out_adj_4273, n11_adj_4274, n11_adj_4275, 
        n5, n23868, n28015, n28014, n28013, n28012, n28011, n28010, 
        n28009, state_7__N_3860, n4860, n24230, n10_adj_4276, n35965, 
        n32204, n10_adj_4277, n28422, n28421, n28420, n28419, n28418, 
        n33132, n12, n34179;
    
    SB_DFFSR counter2_1552_1553__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n18552));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n18362), .D(n119[7]), 
            .R(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n18362), .D(n119[6]), 
            .R(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n18362), .D(n119[5]), 
            .R(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n18362), .D(n119[4]), 
            .R(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n18362), .D(n119[3]), 
            .R(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n18362), .D(n119[2]), 
            .S(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n18362), .D(n119[1]), 
            .S(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n17058));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1491 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n17053));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_1491.LUT_INIT = 16'hfefe;
    SB_LUT4 i30585_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11), .I3(n4867), 
            .O(n24174));   // verilog/i2c_controller.v(151[5:14])
    defparam i30585_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 i29859_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n35961));   // verilog/i2c_controller.v(198[28:35])
    defparam i29859_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i29854_4_lut (.I0(n35961), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n35877));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i29854_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 i29774_4_lut (.I0(n35877), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(n11_adj_4270), .O(n35980));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i29774_4_lut.LUT_INIT = 16'h0322;
    SB_LUT4 i1_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n18487));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(n34), .I1(n37), .I2(GND_net), .I3(GND_net), 
            .O(n39));
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'heeee;
    SB_LUT4 i30436_2_lut (.I0(\state_7__N_3861[0] ), .I1(enable_slow_N_3964), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_3963));   // verilog/i2c_controller.v(62[6:32])
    defparam i30436_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_2_lut_adj_1493 (.I0(i2c_clk), .I1(n18552), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_3950));
    defparam i1_2_lut_adj_1493.LUT_INIT = 16'h6666;
    SB_LUT4 equal_150_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_150_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i30441_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n32132));
    defparam i30441_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i29862_3_lut_4_lut (.I0(n11_adj_4271), .I1(n11), .I2(enable_slow_N_3964), 
            .I3(\state_7__N_3861[0] ), .O(n35900));
    defparam i29862_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 equal_153_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_11));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_153_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i30583_3_lut_4_lut (.I0(n11_adj_4271), .I1(n11), .I2(n15), 
            .I3(n4867), .O(n24476));
    defparam i30583_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_3950));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_3951));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_DFFE enable_slow_120 (.Q(\state_7__N_3861[0] ), .C(CLK_c), .E(n18254), 
            .D(enable_slow_N_3963));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n5184), 
            .D(n10190), .S(n18487));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4273), .C(i2c_clk), .E(n32132), 
            .D(n35980));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_LUT4 i1_4_lut (.I0(n11_adj_4274), .I1(n11_adj_4275), .I2(\state_7__N_3877[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'h5755;
    SB_LUT4 i30521_2_lut (.I0(\state_7__N_3877[3] ), .I1(n11_adj_4275), 
            .I2(GND_net), .I3(GND_net), .O(n23868));
    defparam i30521_2_lut.LUT_INIT = 16'h1111;
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n18362), .D(n119[0]), 
            .S(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i30443_4_lut_4_lut (.I0(\state[2] ), .I1(n11_adj_4270), .I2(\state[1] ), 
            .I3(n39), .O(n5184));
    defparam i30443_4_lut_4_lut.LUT_INIT = 16'hef00;
    SB_LUT4 i30450_2_lut_3_lut (.I0(\state[2] ), .I1(n11_adj_4270), .I2(\state[0] ), 
            .I3(GND_net), .O(n10190));
    defparam i30450_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n28015), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n28014), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_8 (.CI(n28014), .I0(counter[6]), .I1(VCC_net), 
            .CO(n28015));
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n28013), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n28013), .I0(counter[5]), .I1(VCC_net), 
            .CO(n28014));
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n28012), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n28012), .I0(counter[4]), .I1(VCC_net), 
            .CO(n28013));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n28011), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n28011), .I0(counter[3]), .I1(VCC_net), 
            .CO(n28012));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n28010), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n28010), .I0(counter[2]), .I1(VCC_net), 
            .CO(n28011));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n28009), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i18938_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i18938_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i30409_4_lut (.I0(state_7__N_3860), .I1(n4860), .I2(n11_adj_4271), 
            .I3(n24230), .O(n4867));
    defparam i30409_4_lut.LUT_INIT = 16'h5111;
    SB_CARRY sub_39_add_2_3 (.CI(n28009), .I0(counter[1]), .I1(VCC_net), 
            .CO(n28010));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n28009));
    SB_LUT4 i29573_4_lut (.I0(n10_adj_4276), .I1(n10), .I2(\state_7__N_3877[3] ), 
            .I3(enable), .O(n35965));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i29573_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut_adj_1494 (.I0(\state[1] ), .I1(n7), .I2(n35965), 
            .I3(\state[0] ), .O(n32204));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_1494.LUT_INIT = 16'ha088;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_adj_4277));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_adj_4277), .I2(counter2[0]), 
            .I3(GND_net), .O(n18552));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 counter2_1552_1553_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n28422), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1552_1553_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1552_1553_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n28421), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1552_1553_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1552_1553_add_4_6 (.CI(n28421), .I0(GND_net), .I1(counter2[4]), 
            .CO(n28422));
    SB_LUT4 counter2_1552_1553_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n28420), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1552_1553_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1552_1553_add_4_5 (.CI(n28420), .I0(GND_net), .I1(counter2[3]), 
            .CO(n28421));
    SB_LUT4 counter2_1552_1553_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n28419), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1552_1553_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1552_1553_add_4_4 (.CI(n28419), .I0(GND_net), .I1(counter2[2]), 
            .CO(n28420));
    SB_LUT4 counter2_1552_1553_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n28418), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1552_1553_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1552_1553_add_4_3 (.CI(n28418), .I0(GND_net), .I1(counter2[1]), 
            .CO(n28419));
    SB_LUT4 counter2_1552_1553_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1552_1553_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1552_1553_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n28418));
    SB_LUT4 i1803_2_lut (.I0(sda_out_adj_4273), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i1803_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4275));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_LUT4 equal_95_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_95_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4274));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i28574_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_3964));   // verilog/i2c_controller.v(44[32:47])
    defparam i28574_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26806_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n33132), .O(n18604));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i26806_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_12));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_12), 
            .O(n4860));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i26749_2_lut (.I0(\state_7__N_3877[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n33132));
    defparam i26749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n4860), .I1(n33132), .I2(n5300), .I3(n37), 
            .O(n18362));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 equal_93_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4276));   // verilog/i2c_controller.v(44[32:47])
    defparam equal_93_i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i30588_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n4867), .O(n34179));
    defparam i30588_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4271));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i19453_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n24230));
    defparam i19453_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n4867), .D(n32204), 
            .S(n34179));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n4867), .D(n23868), 
            .S(n24174));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n4867), .D(n5), 
            .S(n24476));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n18652));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n18650));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n18649));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n18648));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n18647));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n18646));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1552_1553__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n18552));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i19599_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_3951));   // verilog/i2c_controller.v(44[32:47])
    defparam i19599_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i22_3_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n11_adj_4270));   // verilog/i2c_controller.v(44[32:47])
    defparam i22_3_lut_3_lut.LUT_INIT = 16'h1a1a;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut_adj_1495 (.I0(enable), .I1(\state_7__N_3861[0] ), 
            .I2(enable_slow_N_3964), .I3(GND_net), .O(n18254));
    defparam i1_2_lut_3_lut_adj_1495.LUT_INIT = 16'heaea;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n19174));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i18954_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n23726));
    defparam i18954_2_lut.LUT_INIT = 16'h8888;
    SB_DFFSR counter2_1552_1553__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n18552));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1552_1553__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n18552));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1552_1553__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n18552));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1552_1553__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n18552));   // verilog/i2c_controller.v(69[20:35])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n18633));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n18632));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i19645_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_3860));
    defparam i19645_3_lut_4_lut.LUT_INIT = 16'hf800;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, \data_in_frame[1] , \data_in_frame[2] , rx_data, 
            \data_out_frame[23] , \data_out_frame[25] , \data_out_frame[24] , 
            GND_net, \data_out_frame[20] , \data_out_frame[17] , \data_out_frame[19] , 
            \data_out_frame[15] , \data_out_frame[18] , n32658, \data_in_frame[19] , 
            \data_in_frame[3] , \data_out_frame[10] , \data_out_frame[13] , 
            \data_out_frame[11] , \data_out_frame[6] , \data_out_frame[4] , 
            \data_out_frame[8] , \data_out_frame[12] , \data_out_frame[5] , 
            \data_out_frame[7] , \data_out_frame[9] , \data_in_frame[6] , 
            \data_out_frame[16] , n30832, n32385, n32397, n30803, 
            n32722, n32920, \data_out_frame[14] , n32699, \FRAME_MATCHER.state[0] , 
            n32403, n32412, n66, \data_in_frame[13] , \data_in_frame[17] , 
            \data_in_frame[10] , \data_in_frame[11] , \data_in_frame[8] , 
            \data_in_frame[18] , \data_in_frame[12] , \data_in_frame[9] , 
            \data_in_frame[5] , n63, \FRAME_MATCHER.i_31__N_2461 , n3303, 
            n4452, n34405, rx_data_ready, \data_in_frame[21] , setpoint, 
            \data_in_frame[4] , n123, n1, n18735, n18734, n18733, 
            n18732, n18731, n18730, n18729, n18728, n18727, n18726, 
            n18725, n18724, n18723, n18722, n18721, n18720, n18719, 
            n18718, n18717, n18716, n18715, n18714, n18713, n18712, 
            n18703, n18702, n18701, n18700, n18699, n18698, n18697, 
            n18693, n18692, control_mode, n18691, n18690, n18689, 
            n18688, n18687, n18686, \data_in[0] , \data_in[1] , \data_in[2] , 
            \data_in[3] , n18685, PWMLimit, tx_active, \state[0] , 
            \state[2] , \state[3] , n5300, n32404, n34118, n34304, 
            DE_c, n18684, LED_c, n18683, n18682, n18681, n18680, 
            n18679, n18678, ID, n18677, n18676, n18675, n18674, 
            n18673, n18672, n18671, n18670, n18669, n18668, n18667, 
            n18666, n18665, n18664, n18663, n37934, n19173, IntegralLimit, 
            n19172, n19171, n19170, n19169, n19168, n19167, n19166, 
            n19165, n19164, n19163, n19162, n19161, n19160, n19159, 
            n19158, n19157, n19156, n19155, n19154, n19153, n19152, 
            n19151, n19118, n19117, n19116, n19115, n19114, n19113, 
            n19112, n19111, n19110, n19109, n19108, n19107, n19106, 
            n19105, n19104, n19103, n19102, n19101, n19100, n19099, 
            n19098, n19097, n19096, n19095, n19094, n19093, n19092, 
            n19091, n19090, n19089, n19088, n19087, \Kp[1] , n19086, 
            \Kp[2] , n19085, \Kp[3] , n19084, \Kp[4] , n19083, \Kp[5] , 
            n19082, \Kp[6] , n19081, \Kp[7] , n19080, \Kp[8] , n19079, 
            \Kp[9] , n19078, \Kp[10] , n19077, \Kp[11] , n19076, 
            \Kp[12] , n19075, \Kp[13] , n19074, \Kp[14] , n19073, 
            \Kp[15] , n19072, \Ki[1] , n19071, \Ki[2] , n19070, 
            \Ki[3] , n19069, \Ki[4] , n19068, \Ki[5] , n19067, \Ki[6] , 
            n19066, \Ki[7] , n19065, \Ki[8] , n19064, \Ki[9] , n19063, 
            \Ki[10] , n19062, \Ki[11] , n19061, \Ki[12] , n19060, 
            \Ki[13] , n19059, \Ki[14] , n19058, \Ki[15] , n19057, 
            n19056, n19055, n19054, n19053, n19052, n19051, n19050, 
            n19049, n19048, n19047, n19046, n19045, n19044, n19043, 
            n19042, n19041, n19040, n19039, n19038, n19037, n19036, 
            n19035, n19034, n19033, n19032, n19031, n19030, n19029, 
            n19028, n19027, n19026, n19025, n19024, n19023, n19022, 
            n19021, n19020, n19019, n19018, n19017, n19016, n19015, 
            n19014, n19013, n19012, n19011, n19010, n19009, n19008, 
            n19007, n19006, n19005, n19004, n19003, n19002, n19001, 
            n19000, n18999, n18998, n18997, n18996, n18994, n18993, 
            n18992, n18991, n18990, n18989, n18988, n18987, n18986, 
            n18985, n18984, n18983, n18982, n32395, n32400, n18981, 
            n32409, n18980, n18979, n18978, n18977, n18976, n18975, 
            n18974, n18973, n18972, n18971, n18970, n18969, n18968, 
            n18967, n18966, n18965, n18964, n18963, n18962, n18961, 
            n18960, n18959, n18958, n18957, n18956, n18955, n18954, 
            n18953, n18952, n18951, n18950, n18949, n18948, n18640, 
            n18639, n18637, neopxl_color, n18636, \Ki[0] , n18635, 
            \Kp[0] , n18634, n18947, n18946, n18945, n18944, n18943, 
            n18942, n18941, n18940, n18626, n18939, n18938, n18937, 
            n18936, n18935, n18934, n18933, n18932, n18931, n18930, 
            n18929, n18928, n18927, n18926, n18925, n18924, n18923, 
            n18922, n18921, n18920, n18919, n18918, n18917, n18916, 
            n18915, n18914, n18913, n18912, n18911, n18910, n18909, 
            n18908, n18907, n18906, n18905, n18904, n18903, n18902, 
            n18901, n18900, n18899, n18898, n18897, n18896, n18895, 
            n18894, n18893, n18892, n18891, n18890, n18889, n18888, 
            n18887, n18886, n18885, n18884, n18883, n18882, n18881, 
            n18880, n18879, n18878, n18877, n18876, n18875, n18874, 
            n18866, n18865, n18864, n18863, n18862, n18861, n18860, 
            n18859, n18850, n18849, n18848, n18847, n18846, n18845, 
            n18844, n18843, n18834, n18833, n18832, n18831, n18830, 
            n18829, n18828, n18827, n18802, n18801, n18800, n18799, 
            n18798, n18797, n18796, n18795, n18786, n18785, n18784, 
            n18783, n32831, n18782, n18781, n18780, n18779, n18770, 
            n18769, n18768, n18767, n18766, n18765, n18764, n18763, 
            n29929, n32394, n32410, n32402, n14410, r_SM_Main, n10125, 
            tx_o, \r_SM_Main_2__N_3450[1] , \r_Bit_Index[0] , n18336, 
            n18590, VCC_net, n4, n18644, n18660, n37939, tx_enable, 
            n23776, n4_adj_3, \r_Bit_Index[0]_adj_4 , n17079, n4_adj_5, 
            r_SM_Main_adj_10, \r_SM_Main_2__N_3379[2] , n17084, n4_adj_9, 
            n31970, r_Rx_Data, RX_N_10, n33211, n33251, n19204, 
            n19202, n19201, n19200, n19199, n19198, n19197, n18696, 
            n18995, n32359) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[2] ;
    output [7:0]rx_data;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[24] ;
    input GND_net;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[18] ;
    output n32658;
    output [7:0]\data_in_frame[19] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_out_frame[16] ;
    output n30832;
    output n32385;
    output n32397;
    output n30803;
    output n32722;
    output n32920;
    output [7:0]\data_out_frame[14] ;
    output n32699;
    output \FRAME_MATCHER.state[0] ;
    output n32403;
    output n32412;
    output n66;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[17] ;
    output [7:0]\data_in_frame[10] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[18] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]\data_in_frame[5] ;
    output n63;
    output \FRAME_MATCHER.i_31__N_2461 ;
    output n3303;
    output n4452;
    output n34405;
    output rx_data_ready;
    output [7:0]\data_in_frame[21] ;
    output [23:0]setpoint;
    output [7:0]\data_in_frame[4] ;
    output n123;
    output n1;
    input n18735;
    input n18734;
    input n18733;
    input n18732;
    input n18731;
    input n18730;
    input n18729;
    input n18728;
    input n18727;
    input n18726;
    input n18725;
    input n18724;
    input n18723;
    input n18722;
    input n18721;
    input n18720;
    input n18719;
    input n18718;
    input n18717;
    input n18716;
    input n18715;
    input n18714;
    input n18713;
    input n18712;
    input n18703;
    input n18702;
    input n18701;
    input n18700;
    input n18699;
    input n18698;
    input n18697;
    input n18693;
    input n18692;
    output [7:0]control_mode;
    input n18691;
    input n18690;
    input n18689;
    input n18688;
    input n18687;
    input n18686;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[3] ;
    input n18685;
    output [23:0]PWMLimit;
    output tx_active;
    input \state[0] ;
    input \state[2] ;
    input \state[3] ;
    output n5300;
    output n32404;
    output n34118;
    output n34304;
    output DE_c;
    input n18684;
    output LED_c;
    input n18683;
    input n18682;
    input n18681;
    input n18680;
    input n18679;
    input n18678;
    input [7:0]ID;
    input n18677;
    input n18676;
    input n18675;
    input n18674;
    input n18673;
    input n18672;
    input n18671;
    input n18670;
    input n18669;
    input n18668;
    input n18667;
    input n18666;
    input n18665;
    input n18664;
    input n18663;
    input n37934;
    input n19173;
    output [23:0]IntegralLimit;
    input n19172;
    input n19171;
    input n19170;
    input n19169;
    input n19168;
    input n19167;
    input n19166;
    input n19165;
    input n19164;
    input n19163;
    input n19162;
    input n19161;
    input n19160;
    input n19159;
    input n19158;
    input n19157;
    input n19156;
    input n19155;
    input n19154;
    input n19153;
    input n19152;
    input n19151;
    input n19118;
    input n19117;
    input n19116;
    input n19115;
    input n19114;
    input n19113;
    input n19112;
    input n19111;
    input n19110;
    input n19109;
    input n19108;
    input n19107;
    input n19106;
    input n19105;
    input n19104;
    input n19103;
    input n19102;
    input n19101;
    input n19100;
    input n19099;
    input n19098;
    input n19097;
    input n19096;
    input n19095;
    input n19094;
    input n19093;
    input n19092;
    input n19091;
    input n19090;
    input n19089;
    input n19088;
    input n19087;
    output \Kp[1] ;
    input n19086;
    output \Kp[2] ;
    input n19085;
    output \Kp[3] ;
    input n19084;
    output \Kp[4] ;
    input n19083;
    output \Kp[5] ;
    input n19082;
    output \Kp[6] ;
    input n19081;
    output \Kp[7] ;
    input n19080;
    output \Kp[8] ;
    input n19079;
    output \Kp[9] ;
    input n19078;
    output \Kp[10] ;
    input n19077;
    output \Kp[11] ;
    input n19076;
    output \Kp[12] ;
    input n19075;
    output \Kp[13] ;
    input n19074;
    output \Kp[14] ;
    input n19073;
    output \Kp[15] ;
    input n19072;
    output \Ki[1] ;
    input n19071;
    output \Ki[2] ;
    input n19070;
    output \Ki[3] ;
    input n19069;
    output \Ki[4] ;
    input n19068;
    output \Ki[5] ;
    input n19067;
    output \Ki[6] ;
    input n19066;
    output \Ki[7] ;
    input n19065;
    output \Ki[8] ;
    input n19064;
    output \Ki[9] ;
    input n19063;
    output \Ki[10] ;
    input n19062;
    output \Ki[11] ;
    input n19061;
    output \Ki[12] ;
    input n19060;
    output \Ki[13] ;
    input n19059;
    output \Ki[14] ;
    input n19058;
    output \Ki[15] ;
    input n19057;
    input n19056;
    input n19055;
    input n19054;
    input n19053;
    input n19052;
    input n19051;
    input n19050;
    input n19049;
    input n19048;
    input n19047;
    input n19046;
    input n19045;
    input n19044;
    input n19043;
    input n19042;
    input n19041;
    input n19040;
    input n19039;
    input n19038;
    input n19037;
    input n19036;
    input n19035;
    input n19034;
    input n19033;
    input n19032;
    input n19031;
    input n19030;
    input n19029;
    input n19028;
    input n19027;
    input n19026;
    input n19025;
    input n19024;
    input n19023;
    input n19022;
    input n19021;
    input n19020;
    input n19019;
    input n19018;
    input n19017;
    input n19016;
    input n19015;
    input n19014;
    input n19013;
    input n19012;
    input n19011;
    input n19010;
    input n19009;
    input n19008;
    input n19007;
    input n19006;
    input n19005;
    input n19004;
    input n19003;
    input n19002;
    input n19001;
    input n19000;
    input n18999;
    input n18998;
    input n18997;
    input n18996;
    input n18994;
    input n18993;
    input n18992;
    input n18991;
    input n18990;
    input n18989;
    input n18988;
    input n18987;
    input n18986;
    input n18985;
    input n18984;
    input n18983;
    input n18982;
    output n32395;
    output n32400;
    input n18981;
    output n32409;
    input n18980;
    input n18979;
    input n18978;
    input n18977;
    input n18976;
    input n18975;
    input n18974;
    input n18973;
    input n18972;
    input n18971;
    input n18970;
    input n18969;
    input n18968;
    input n18967;
    input n18966;
    input n18965;
    input n18964;
    input n18963;
    input n18962;
    input n18961;
    input n18960;
    input n18959;
    input n18958;
    input n18957;
    input n18956;
    input n18955;
    input n18954;
    input n18953;
    input n18952;
    input n18951;
    input n18950;
    input n18949;
    input n18948;
    input n18640;
    input n18639;
    input n18637;
    output [23:0]neopxl_color;
    input n18636;
    output \Ki[0] ;
    input n18635;
    output \Kp[0] ;
    input n18634;
    input n18947;
    input n18946;
    input n18945;
    input n18944;
    input n18943;
    input n18942;
    input n18941;
    input n18940;
    input n18626;
    input n18939;
    input n18938;
    input n18937;
    input n18936;
    input n18935;
    input n18934;
    input n18933;
    input n18932;
    input n18931;
    input n18930;
    input n18929;
    input n18928;
    input n18927;
    input n18926;
    input n18925;
    input n18924;
    input n18923;
    input n18922;
    input n18921;
    input n18920;
    input n18919;
    input n18918;
    input n18917;
    input n18916;
    input n18915;
    input n18914;
    input n18913;
    input n18912;
    input n18911;
    input n18910;
    input n18909;
    input n18908;
    input n18907;
    input n18906;
    input n18905;
    input n18904;
    input n18903;
    input n18902;
    input n18901;
    input n18900;
    input n18899;
    input n18898;
    input n18897;
    input n18896;
    input n18895;
    input n18894;
    input n18893;
    input n18892;
    input n18891;
    input n18890;
    input n18889;
    input n18888;
    input n18887;
    input n18886;
    input n18885;
    input n18884;
    input n18883;
    input n18882;
    input n18881;
    input n18880;
    input n18879;
    input n18878;
    input n18877;
    input n18876;
    input n18875;
    input n18874;
    input n18866;
    input n18865;
    input n18864;
    input n18863;
    input n18862;
    input n18861;
    input n18860;
    input n18859;
    input n18850;
    input n18849;
    input n18848;
    input n18847;
    input n18846;
    input n18845;
    input n18844;
    input n18843;
    input n18834;
    input n18833;
    input n18832;
    input n18831;
    input n18830;
    input n18829;
    input n18828;
    input n18827;
    input n18802;
    input n18801;
    input n18800;
    input n18799;
    input n18798;
    input n18797;
    input n18796;
    input n18795;
    input n18786;
    input n18785;
    input n18784;
    input n18783;
    output n32831;
    input n18782;
    input n18781;
    input n18780;
    input n18779;
    input n18770;
    input n18769;
    input n18768;
    input n18767;
    input n18766;
    input n18765;
    input n18764;
    input n18763;
    input n29929;
    output n32394;
    output n32410;
    output n32402;
    output n14410;
    output [2:0]r_SM_Main;
    output n10125;
    output tx_o;
    output \r_SM_Main_2__N_3450[1] ;
    output \r_Bit_Index[0] ;
    output n18336;
    output n18590;
    input VCC_net;
    output n4;
    input n18644;
    input n18660;
    input n37939;
    output tx_enable;
    output n23776;
    output n4_adj_3;
    output \r_Bit_Index[0]_adj_4 ;
    output n17079;
    output n4_adj_5;
    output [2:0]r_SM_Main_adj_10;
    output \r_SM_Main_2__N_3379[2] ;
    output n17084;
    output n4_adj_9;
    input n31970;
    output r_Rx_Data;
    input RX_N_10;
    output n33211;
    output n33251;
    input n19204;
    input n19202;
    input n19201;
    input n19200;
    input n19199;
    input n19198;
    input n19197;
    input n18696;
    input n18995;
    input n32359;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n18759;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n18758;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n17751, n10, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n18757, n18756, n8, n32398;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n18709, n18710, n32975, n32772, n34432, n34610, n15386, 
        n30801, n30046, n12, n2332, n30287, n33462, n32778, n7, 
        n30912, n32978, n34435, n32740, n32741, n30860, n32799, 
        n6, n34686, n32661, n32910, n30936, n32900, n30792, n30907, 
        n30836, n32507, n30788, n7_adj_3968, n33385, n32951, n34825, 
        n7_adj_3969, n30856, n16652, n18711, n29942, n33036, n32725, 
        n30090, n32788, n18755, n32529, n29901, n32728, n6_adj_3970, 
        n32914, n33038, n32664, n33044, n32923, n5063, n5064, 
        n17483, n32584, n32851, n17610, n14, n18108, n32564, n32860, 
        n15, n17101, n17678, n17104, n32550, n1193, n2394, n17250, 
        n32936, n16, n32687, n17, n30783, n32706, n32945, n54, 
        n32817, n32746, n32785, n42, n32990, n32690, n32814, n32511, 
        n40, n33078, n29940, n32891, n41, n32822, n39, n32854, 
        n48, n32872, n33030, n32999, n46, n32438, n18067, n47, 
        n33014, n45, n33027, n44, n32894, n43, n54_adj_3971, Kp_23__N_933, 
        n17376, Kp_23__N_1032, n49, n34766, n32546, n32443, n43_adj_3972, 
        n48_adj_3973, n30019, n32620, n17807, n28, n17534, n38, 
        n17693, n47_adj_3974, n32, n17664, n32674, n30, n18111, 
        n29979, n31, n32843, n17354, n29, n34718, n33521, n44_adj_3975, 
        n29870, n32671, n58, n29938, n62, n60, n32556, n61, 
        n32498, n59, n56, n30798, n34478, n64, n68, n32737, 
        n55, n6_adj_3976, n32837, n29984, n32608, n12_adj_3977, 
        n1130, n32840, n32981, n12_adj_3978, n16767, n33836, n30869, 
        n32539, n32596, n32617, n12_adj_3979, n33041, n10_adj_3980, 
        n32782, n30024, n32384, Kp_23__N_825, n16267, n17222;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n32590, n32391, n17297, n16793, n17886, n32993, n12_adj_3981, 
        n1169, n2063, n30867, n10_adj_3982, n32428, n6_adj_3983, 
        n32802, n10_adj_3984, n18754;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    
    wire n32939, n6_adj_3985, n15336, n32825, n29969, n18032, n17810, 
        n6_adj_3986, n34449, n33054, n29949, n10_adj_3987, n30811, 
        n33862, n32805, n33072, n6_adj_3988, n32463, n17098, n1191, 
        n1168, n32885, n10_adj_3989, n33569, n32996, n17207, n6_adj_3990, 
        n29953, n33011, n17883, n32984, n32460, n12_adj_3991, n32561, 
        n14_adj_3992, n10_adj_3993, n16700, n33517, n17711, n10_adj_3994, 
        n17108, n16_adj_3995, n17_adj_3996, n14_adj_3997, n10_adj_3998, 
        n33075, n15_adj_3999, n14_adj_4000, n16_adj_4001, n17_adj_4002, 
        n6_adj_4003, n32425, n8_adj_4004;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n8_adj_4005, n24776, n32378, n18277, n33621, n32491, n6_adj_4006, 
        Kp_23__N_806, n32478, n26, n17177, n24, n29_adj_4007, n21, 
        n4_c, n14565, n32_adj_4008, n32505, n27, n34988;
    wire [31:0]\FRAME_MATCHER.state_31__N_2561 ;
    
    wire n4_adj_4009, n2_adj_4010, n1_c, n5, n17092, n31898, n32406, 
        n5_adj_4011, n31890, n31888, n31832, n31834, n31886, n31884, 
        n31882, n31880, n31878, n31876, n31874, n31836, n31838, 
        n31820, n31872, n31870, n31868, n18753, n31866, n8_adj_4012, 
        n8_adj_4013, n31864, n31862, n31860, n31892, n31858, n8_adj_4014, 
        n8_adj_4015, \FRAME_MATCHER.i_31__N_2463 , n8_adj_4016, n18752, 
        n18751, n18750, n18749, n32452, n6_adj_4017, n32766, n10_adj_4018;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n30504, n17198, n30884, n33063, n46_adj_4019, n32655, n32794, 
        n32455, n42_adj_4020;
    wire [7:0]n8825;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n27756, n32757, n17187, n28_adj_4021, n33084, n32494, n32927, 
        n26_adj_4022, n17427, n33081, n17447, n32933, n27_adj_4023, 
        n34667, n33050, n25, n34390, Kp_23__N_1335, n34, n32888, 
        n30314, n33005, n43_adj_4024, n32501, n36, n32650, n50, 
        n33069, n33066, n48_adj_4025, n32828, n32763, n49_adj_4026, 
        n17758, n47_adj_4027, n17579, n6_adj_4028, Kp_23__N_698, n32791, 
        n32905, n5_adj_4029, n32611, n32693, n12_adj_4030, n32942, 
        n34750, n6_adj_4031, n33060, n30809, n32743, n32957, n10_adj_4032, 
        n5_adj_4033, n32714, n34722, n32987, Kp_23__N_1170, n6_adj_4034, 
        n32963, n33047, n29843, n6_adj_4035, n32966, n15471, n12_adj_4036, 
        n30921, n10_adj_4037, n15478, n32972, n18035, n5087, n5086, 
        n5085, n32834, n10_adj_4038, n17842, Kp_23__N_1373, n32760, 
        n30777, n29856, n12_adj_4039, n33033, n5084, n5083, n5082, 
        n30005, n6_adj_4040, n32731, n10_adj_4041, n17434, n30823, 
        n17705, n5081, n5080, n5079, n32614, n5078, n5077, n5076, 
        n32577, n5075, n17814, n17128, n12_adj_4042, n5074, n30259, 
        n33438, n13, n32623, n5073, n5072, n17364, n32647, n32845, 
        n18, n17396, n20, n33008, n16_adj_4043, n32677, n32775, 
        n27755, n17342, n32645, n12_adj_4044, n5071, n28_adj_4045, 
        n5070, n33017, n26_adj_4046, n33024, n32863, n27_adj_4047, 
        n30001, n25_adj_4048, n5069, n34613, n32683, n5068, n5067, 
        n5066, n32930, n17358, n6_adj_4049, n17246, n6_adj_4050, 
        n17316, n17867, n16_adj_4051, n30028, n32880, n17745, n17_adj_4052, 
        n29907, n29854, n32571, n4_adj_4053, n10_adj_4054, n17212, 
        n17370, n33002, n10_adj_4055, n32602, n32475, n10_adj_4056, 
        n18748, n63_c, n63_adj_4057;
    wire [31:0]n92;
    
    wire n38282, n30543, n10_adj_4059, n5_adj_4060, n10_adj_4061, 
        Kp_23__N_1167, n1_adj_4062, n33978, n8_adj_4063, n5_adj_4064, 
        n37935, n17589, n17926, n6_adj_4065, n17418, n29850, n32667, 
        n12_adj_4066, n32917, n6_adj_4067, n8_adj_4068;
    wire [0:0]n3519;
    wire [2:0]r_SM_Main_2__N_3453;
    
    wire n3482, n32960, n14_adj_4069, n10_adj_4070, n17699, \FRAME_MATCHER.rx_data_ready_prev , 
        n31814, n33985, n18744, n18216, n20456, n30854, n38031, 
        n12_adj_4071, n8_adj_4072, n10_adj_4073, n18743, n10_adj_4074, 
        n6_adj_4075, n32709, n10_adj_4076, n12_adj_4077, n11, n6_adj_4078, 
        n34561, n34494, n19, n16_adj_4079, n17_adj_4080, n35893, 
        n35892, n10_adj_4081, n12_adj_4082, n16_adj_4083, n34814, 
        n8_adj_4084, n33574, Kp_23__N_901, n38040, n14_adj_4085, n13_adj_4086, 
        n18241, n34784, n23, n18742, n13_adj_4087, n16_adj_4088, 
        n11_adj_4089, n10_adj_4090, n2_adj_4091, n27717, n2236, n34764, 
        n18741, n6_adj_4092, n10_adj_4093, n33866, n34823, n5065, 
        n34774, n26_adj_4094, n32808, n17_adj_4095, n27718, n22, 
        n28_adj_4096, n21_adj_4097, n17768, n29_adj_4098, n31_adj_4099, 
        n27754, n6_adj_4100, n32487, n6_adj_4101, n30895, n32638, 
        n32866, n17590, n32848, n17742, n6_adj_4102, n32877, n32567, 
        n12_adj_4103, n32574, n32642, n29905, n17466, Kp_23__N_930, 
        n8_adj_4104, n18736, n18737, n17324, n18738, n2_adj_4105, 
        n27716, n18739, n17731, n17237, n18740, n27753, n2_adj_4106, 
        n27715, n2_adj_4107, n27714, n27752, n2_adj_4108, n27713, 
        n7_adj_4109, n7_adj_4110, n7_adj_4111, n31964, n31962, n31960, 
        n31958, n31956, n7_adj_4112, n7_adj_4113, n31954, n31952, 
        n31950, n31948, n31946, n31944, n31942, n31940, n31938, 
        n31936, n31934, n31932, n31930, n31928, n31926, n31924, 
        n31922, n31920, n31816, n771, n32373, \FRAME_MATCHER.i_31__N_2457 , 
        n27751;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n18102, n32587, n32826, n34574, n33844, n33843;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n32721, n33395, n2_adj_4115, n3_adj_4116, n2_adj_4117, n27712, 
        n17785, n10_adj_4118, n15437, n32521, n17761, n32525, n32518, 
        n32534, n2_adj_4119, n3_adj_4120, n2_adj_4121, n3_adj_4122, 
        n2_adj_4123, n3_adj_4124, n2_adj_4125, n3_adj_4126, n2_adj_4127, 
        n3_adj_4128, n2_adj_4129, n3_adj_4130, n2_adj_4131, n3_adj_4132, 
        n2_adj_4133, n3_adj_4134, n35078, n35079, n2_adj_4135, n3_adj_4136, 
        n3_adj_4137, n3_adj_4138, n3_adj_4139, n3_adj_4140, n3_adj_4141, 
        n3_adj_4142, n2_adj_4143, n3_adj_4144, n2_adj_4145, n3_adj_4146, 
        n2_adj_4147, n3_adj_4148, n2_adj_4149, n3_adj_4150, n35077, 
        n2_adj_4151, n3_adj_4152, n2_adj_4153, n3_adj_4154, n2_adj_4155, 
        n3_adj_4156, n2_adj_4157, n3_adj_4158, n27750, n2_adj_4159, 
        n3_adj_4160, n2_adj_4161, n3_adj_4162, n2_adj_4163, n3_adj_4164, 
        n2_adj_4165, n3_adj_4166, n2_adj_4167, n3_adj_4168, n2_adj_4169, 
        n3_adj_4170, n2_adj_4171, n3_adj_4172, n37469, n37613, n14_adj_4173, 
        n37589, n35901, n16_adj_4174, n17_adj_4175, n35875, n35874, 
        n16_adj_4176, n17_adj_4177, n35903, n35902, n27711, n16_adj_4178, 
        tx_transmit_N_3350, n17_adj_4179, n27710, n35869, n35868, 
        n27709, n32553, n16_adj_4180, n17_adj_4181, n10_adj_4182, 
        n14_adj_4183, n24578, n24390, n20_adj_4184, n19_adj_4185, 
        n38_adj_4186, n21_adj_4187, n24690, n17001, n1_adj_4188, n10_adj_4189, 
        n17017, n34324, n161, n17068, n17089, n24219, n10_adj_4190, 
        n27708, n27707, n18708, n18707, n5202, n5_adj_4191, n6_adj_4192, 
        n32337, n18706, n18705, n18704, n32605, n32869, n30_adj_4193, 
        n34_adj_4194, n27706, n32_adj_4195, n35909, n35908, n27705, 
        n77, n33, n31_adj_4196, n27704, n24682, n10932, n34998, 
        \FRAME_MATCHER.i_31__N_2460 , n17014, n16911, n5_adj_4197, n34138, 
        n17065, n12_adj_4198, n16914, n10_adj_4199, n16_adj_4200, 
        n17_adj_4201, n27703, n7_adj_4202, n17011, n10_adj_4203, n14_adj_4204, 
        n17008, n18_adj_4205, n20_adj_4206, n15_adj_4207, n16_adj_4208, 
        n17_adj_4209, n14_adj_4210, n34684, n15_adj_4211, n44_adj_4212, 
        n42_adj_4213, n43_adj_4214, n41_adj_4215, n40_adj_4216, n39_adj_4217, 
        n50_adj_4218, n35112, n35110, n7_adj_4219, n45_adj_4220, n8_adj_4221, 
        n14278;
    wire [31:0]\FRAME_MATCHER.state_31__N_2497 ;
    
    wire n33875, n4_adj_4222, n35103, n35101, n7_adj_4223, n35097, 
        n35095, n7_adj_4224, n23655, n24235, n74, n47_adj_4225, 
        n34921, n62_adj_4226, n35073, n35071, n7_adj_4227, n8_adj_4228, 
        n7_adj_4229, n10_adj_4230, n35085, n35083, n7_adj_4231, n27702, 
        n27701, n6_adj_4232, n27700, n35091, n35089, n7_adj_4233, 
        n27699, n35070, n35068, n7_adj_4234, n18867, n27698, n18868, 
        n27697, n18869, n37610, n37349, n35870, n37604, n14_adj_4235;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n37598, n37601, n37361, n35864, n37592, n14_adj_4236, n37586, 
        n37580, n18870, n18460, n18871, n37583, n1_adj_4237, n37574, 
        n37577, n37568, n37571, n37562, n37565, n37556, n37559, 
        n37550, n37553, n18872, n18873, n31_adj_4238, n18638, n37532, 
        n37535, n37526, n37529, n37520, n37523, n37514, n37517, 
        n37508, n37511, n37502, n37505, n17391, n37496, n37499, 
        n37490, n10_adj_4239, n18851, n18852, n18853, n18854, n18855, 
        n18856, n37493, n18857, n37367, n35907, n37484, n14_adj_4240, 
        n37466, n37454, n37457, n37448, n37451, n17820, n37439, 
        n35904, n37442, n14_adj_4241, n18858, n35905, n35906, n37436, 
        n17_adj_4242, n16_adj_4243, n37430, n37433, n37373, n35861, 
        n37412, n14_adj_4244, n37406, n37409, n12_adj_4245, n34602, 
        n18835, n18836, n18837, n18838, n18839, n37379, n35912, 
        n37400, n14_adj_4246, n37385, n35891, n37394, n14_adj_4247, 
        n18840, n37388, n18841, n18470, n34936, n18_adj_4248, n18842, 
        n26_adj_4249, n37391, n27727, n35002, n23_adj_4250, n27_adj_4251, 
        n29_adj_4252, n27726, n27725, n37382, n8_adj_4253, n18819, 
        n12_adj_4254, n18820, n18821, n18822, n18823, n18824, n27724, 
        n18825, n18826, n33579, n18811, n18812, n10_adj_4255, n18813, 
        n11_adj_4256, n9, n32415, n18814, n18815, n18816, n18817, 
        n18818, n18803, n18804, n18805, n18806, n14047, n18807, 
        n18808, n18809, n18810, n27723, n27722, n32580, n16_adj_4257, 
        n17_adj_4258, n35927, n35928, n37376, n18787, n18788, n18789, 
        n18790, n18791, n18792, n18793, n27721, n18794, n27720, 
        n27719, n17_adj_4259, n16_adj_4260, n18760, n18761, n35096, 
        n18762, n35862, n35863, n37370, n18771, n18772, n18773, 
        n18774, n18775, n18776, n18777, n18778, n37364, n35069, 
        n37331, n37358, n37352, n36443, n37346, n35090, n35084, 
        n37328, n37322;
    
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n18759));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n18758));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(n17751), .O(n10));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n18757));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n18756));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13920_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n18709));
    defparam i13920_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13921_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n18710));
    defparam i13921_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut (.I0(\data_out_frame[23] [6]), .I1(n32975), .I2(n32772), 
            .I3(\data_out_frame[25] [7]), .O(n34432));
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n34610), .I1(n15386), .I2(n30801), .I3(n30046), 
            .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut (.I0(n2332), .I1(n12), .I2(n30287), .I3(\data_out_frame[25] [7]), 
            .O(n33462));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut (.I0(\data_out_frame[24] [1]), .I1(n32778), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_843 (.I0(n7), .I1(\data_out_frame[24] [0]), .I2(n30912), 
            .I3(n32978), .O(n34435));
    defparam i4_4_lut_adj_843.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut (.I0(n30287), .I1(n32740), .I2(GND_net), .I3(GND_net), 
            .O(n32741));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_844 (.I0(n30860), .I1(\data_out_frame[24] [2]), 
            .I2(n32799), .I3(n6), .O(n34686));
    defparam i4_4_lut_adj_844.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut (.I0(n32661), .I1(n32910), .I2(n30936), .I3(GND_net), 
            .O(n34610));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_845 (.I0(n32900), .I1(\data_out_frame[20] [2]), 
            .I2(n32778), .I3(GND_net), .O(n32661));
    defparam i2_3_lut_adj_845.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_846 (.I0(n30792), .I1(\data_out_frame[20] [1]), 
            .I2(n30907), .I3(GND_net), .O(n15386));
    defparam i2_3_lut_adj_846.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_847 (.I0(n30836), .I1(n32507), .I2(n30801), .I3(n30788), 
            .O(n30046));
    defparam i3_4_lut_adj_847.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_848 (.I0(n7_adj_3968), .I1(n30046), .I2(n33385), 
            .I3(n32951), .O(n34825));
    defparam i4_4_lut_adj_848.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_849 (.I0(\data_out_frame[24] [0]), .I1(\data_out_frame[23] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_3969));
    defparam i2_2_lut_adj_849.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_850 (.I0(n7_adj_3969), .I1(n30856), .I2(n16652), 
            .I3(n30912), .O(n32507));
    defparam i4_4_lut_adj_850.LUT_INIT = 16'h6996;
    SB_LUT4 i13922_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n18711));
    defparam i13922_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_851 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[19] [6]), 
            .I2(n29942), .I3(GND_net), .O(n32778));
    defparam i2_3_lut_adj_851.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_852 (.I0(\data_out_frame[23] [7]), .I1(n33036), 
            .I2(GND_net), .I3(GND_net), .O(n32725));
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_853 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n32740));
    defparam i1_2_lut_adj_853.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut (.I0(\data_out_frame[19] [4]), .I1(n30090), .I2(n32788), 
            .I3(\data_out_frame[17] [3]), .O(n30860));
    defparam i1_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n18755));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_854 (.I0(n30912), .I1(n30860), .I2(GND_net), 
            .I3(GND_net), .O(n32772));
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_855 (.I0(\data_out_frame[15] [2]), .I1(n32529), 
            .I2(\data_out_frame[15] [1]), .I3(n29901), .O(n30090));
    defparam i3_4_lut_adj_855.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_856 (.I0(\data_out_frame[19] [5]), .I1(n30090), 
            .I2(n29942), .I3(GND_net), .O(n32728));
    defparam i2_3_lut_adj_856.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_857 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[15] [5]), 
            .I2(n6_adj_3970), .I3(\data_out_frame[17] [6]), .O(n32900));
    defparam i1_4_lut_adj_857.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_out_frame[18] [0]), .I1(\data_out_frame[19] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n32914));
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_859 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [4]), 
            .I2(n32658), .I3(\data_out_frame[20] [3]), .O(n32910));
    defparam i1_4_lut_adj_859.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_860 (.I0(\data_out_frame[20] [2]), .I1(n32910), 
            .I2(GND_net), .I3(GND_net), .O(n33038));
    defparam i1_2_lut_adj_860.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_861 (.I0(n32664), .I1(n33044), .I2(n32923), .I3(n32914), 
            .O(n30792));
    defparam i3_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1351_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n5063), .I3(GND_net), .O(n5064));
    defparam mux_1351_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_862 (.I0(n33036), .I1(n30792), .I2(n33038), .I3(\data_out_frame[20] [1]), 
            .O(n30936));
    defparam i1_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_863 (.I0(\data_out_frame[24] [3]), .I1(n30936), 
            .I2(GND_net), .I3(GND_net), .O(n32799));
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_864 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17483));
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_865 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n32584));
    defparam i1_2_lut_adj_865.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_866 (.I0(\data_out_frame[15] [3]), .I1(n32529), 
            .I2(GND_net), .I3(GND_net), .O(n32851));
    defparam i1_2_lut_adj_866.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[13] [1]), 
            .I2(n17610), .I3(GND_net), .O(n14));   // verilog/coms.v(76[16:43])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_867 (.I0(\data_out_frame[11] [0]), .I1(n18108), 
            .I2(n32564), .I3(n32860), .O(n15));   // verilog/coms.v(76[16:43])
    defparam i6_4_lut_adj_867.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(n17101), .I2(n14), .I3(n17678), 
            .O(n32529));   // verilog/coms.v(76[16:43])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_868 (.I0(\data_out_frame[6] [1]), .I1(n17104), 
            .I2(GND_net), .I3(GND_net), .O(n17101));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_869 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32550));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_870 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(n1193), .O(n32564));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_871 (.I0(n2394), .I1(\data_out_frame[25] [2]), 
            .I2(n17250), .I3(n32936), .O(n16));
    defparam i6_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n30788), .I1(n32687), .I2(\data_out_frame[25] [1]), 
            .I3(\data_out_frame[25] [7]), .O(n17));
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(n30856), .I2(n16), .I3(n30783), 
            .O(n32951));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 equal_127_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_127_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i19_4_lut (.I0(\data_out_frame[24] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(n32706), .I3(n32945), .O(n54));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n32817), .I1(n32746), .I2(n32785), .I3(n32564), 
            .O(n42));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n32990), .I1(n32690), .I2(n32814), .I3(n32511), 
            .O(n40));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(\data_out_frame[12] [0]), .I1(n33078), .I2(n29940), 
            .I3(n32891), .O(n41));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(\data_out_frame[11] [2]), .I1(n32550), .I2(n32822), 
            .I3(\data_out_frame[8] [4]), .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[4] [6]), .I3(n32854), .O(n48));   // verilog/coms.v(75[16:43])
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(n32872), .I1(n33030), .I2(\data_out_frame[7] [7]), 
            .I3(n32999), .O(n46));   // verilog/coms.v(75[16:43])
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_872 (.I0(n32438), .I1(\data_out_frame[7] [1]), 
            .I2(n18067), .I3(n32550), .O(n47));   // verilog/coms.v(75[16:43])
    defparam i19_4_lut_adj_872.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_873 (.I0(\data_out_frame[9] [4]), .I1(n33014), 
            .I2(\data_out_frame[9] [2]), .I3(\data_out_frame[7] [4]), .O(n45));   // verilog/coms.v(75[16:43])
    defparam i17_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_874 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[8] [5]), 
            .I2(n33027), .I3(\data_out_frame[9] [6]), .O(n44));   // verilog/coms.v(75[16:43])
    defparam i16_4_lut_adj_874.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_875 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[9] [3]), 
            .I2(n32894), .I3(\data_out_frame[9] [0]), .O(n43));   // verilog/coms.v(75[16:43])
    defparam i15_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54_adj_3971));   // verilog/coms.v(75[16:43])
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_876 (.I0(Kp_23__N_933), .I1(\data_in_frame[6] [4]), 
            .I2(n17376), .I3(GND_net), .O(Kp_23__N_1032));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_LUT4 i21_4_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [7]), 
            .I2(\data_out_frame[6] [3]), .I3(n17101), .O(n49));   // verilog/coms.v(75[16:43])
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54_adj_3971), .I2(n43), .I3(n44), 
            .O(n34766));   // verilog/coms.v(75[16:43])
    defparam i27_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_877 (.I0(n32546), .I1(n34766), .I2(n32443), 
            .I3(\data_out_frame[11] [3]), .O(n43_adj_3972));
    defparam i18_4_lut_adj_877.LUT_INIT = 16'h9669;
    SB_LUT4 i23_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n48_adj_3973));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n30019), .I1(n32620), .I2(n32923), .I3(n17807), 
            .O(n28));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n43_adj_3972), .I1(n17534), .I2(n38), .I3(n17693), 
            .O(n47_adj_3974));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_878 (.I0(n47_adj_3974), .I1(n28), .I2(n32584), 
            .I3(n48_adj_3973), .O(n32));
    defparam i14_4_lut_adj_878.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut (.I0(n17664), .I1(\data_out_frame[16] [1]), .I2(n32674), 
            .I3(\data_out_frame[17] [2]), .O(n30));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut (.I0(n18111), .I1(n29979), .I2(n32511), .I3(\data_out_frame[17] [1]), 
            .O(n31));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut (.I0(\data_out_frame[17] [5]), .I1(n32843), .I2(n17354), 
            .I3(\data_out_frame[17] [6]), .O(n29));
    defparam i11_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i17_4_lut_adj_879 (.I0(n29), .I1(n31), .I2(n30), .I3(n32), 
            .O(n34718));
    defparam i17_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 i9_2_lut (.I0(n33521), .I1(n16652), .I2(GND_net), .I3(GND_net), 
            .O(n44_adj_3975));
    defparam i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i23_4_lut_adj_880 (.I0(\data_out_frame[24] [4]), .I1(n29870), 
            .I2(n32671), .I3(n32778), .O(n58));
    defparam i23_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i27_4_lut_adj_881 (.I0(\data_out_frame[18] [6]), .I1(n54), .I2(n29938), 
            .I3(n32799), .O(n62));
    defparam i27_4_lut_adj_881.LUT_INIT = 16'h9669;
    SB_LUT4 i25_4_lut (.I0(\data_out_frame[19] [1]), .I1(n32851), .I2(n34718), 
            .I3(n32772), .O(n60));
    defparam i25_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut_adj_882 (.I0(n32674), .I1(\data_out_frame[18] [1]), 
            .I2(n32556), .I3(\data_out_frame[18] [7]), .O(n61));
    defparam i26_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(\data_out_frame[18] [3]), .I1(n32728), .I2(n32914), 
            .I3(n32498), .O(n59));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_883 (.I0(n32978), .I1(n32740), .I2(n32900), 
            .I3(n32725), .O(n56));
    defparam i21_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n30798), .I1(n58), .I2(n44_adj_3975), .I3(n34478), 
            .O(n64));
    defparam i29_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i33_4_lut (.I0(n59), .I1(n61), .I2(n60), .I3(n62), .O(n68));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_884 (.I0(n32737), .I1(n30832), .I2(\data_out_frame[18] [2]), 
            .I3(\data_out_frame[24] [5]), .O(n55));
    defparam i20_4_lut_adj_884.LUT_INIT = 16'h9669;
    SB_LUT4 i34_4_lut (.I0(n55), .I1(n68), .I2(n64), .I3(n56), .O(n30801));
    defparam i34_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_885 (.I0(n30801), .I1(n32951), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3976));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_886 (.I0(n30836), .I1(n30788), .I2(n32507), .I3(n6_adj_3976), 
            .O(n32837));
    defparam i4_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_887 (.I0(n29984), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33044));
    defparam i1_2_lut_adj_887.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_888 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[11] [0]), .I3(GND_net), .O(n32891));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_888.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_889 (.I0(n32608), .I1(n32891), .I2(\data_out_frame[13] [2]), 
            .I3(\data_out_frame[6] [6]), .O(n12_adj_3977));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_890 (.I0(\data_out_frame[9] [0]), .I1(n12_adj_3977), 
            .I2(n33030), .I3(n1130), .O(n17534));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_891 (.I0(\data_out_frame[15] [4]), .I1(n17534), 
            .I2(n32511), .I3(GND_net), .O(n32840));
    defparam i2_3_lut_adj_891.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_892 (.I0(n32840), .I1(n32981), .I2(\data_out_frame[18] [0]), 
            .I3(n17693), .O(n12_adj_3978));
    defparam i5_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_893 (.I0(\data_out_frame[17] [7]), .I1(n12_adj_3978), 
            .I2(n33044), .I3(\data_out_frame[17] [6]), .O(n16652));
    defparam i6_4_lut_adj_893.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_894 (.I0(n16652), .I1(n30836), .I2(GND_net), 
            .I3(GND_net), .O(n16767));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_895 (.I0(n29938), .I1(\data_out_frame[23] [0]), 
            .I2(n33836), .I3(\data_out_frame[24] [6]), .O(n32706));
    defparam i3_4_lut_adj_895.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_896 (.I0(\data_out_frame[25] [0]), .I1(n32706), 
            .I2(n16767), .I3(n30907), .O(n33385));
    defparam i3_4_lut_adj_896.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_897 (.I0(\data_out_frame[25] [1]), .I1(n33385), 
            .I2(GND_net), .I3(GND_net), .O(n30869));
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_898 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32923));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_899 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n32539));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_900 (.I0(n32596), .I1(n32617), .I2(\data_out_frame[13] [3]), 
            .I3(n32539), .O(n12_adj_3979));
    defparam i5_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_901 (.I0(\data_out_frame[10] [7]), .I1(n12_adj_3979), 
            .I2(n32894), .I3(\data_out_frame[11] [1]), .O(n17693));
    defparam i6_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_902 (.I0(n32511), .I1(n29984), .I2(GND_net), 
            .I3(GND_net), .O(n32843));
    defparam i1_2_lut_adj_902.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_903 (.I0(\data_out_frame[18] [1]), .I1(n33041), 
            .I2(n32843), .I3(n17693), .O(n10_adj_3980));
    defparam i4_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_904 (.I0(n32782), .I1(n32981), .I2(n30024), .I3(GND_net), 
            .O(n34478));
    defparam i2_3_lut_adj_904.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_905 (.I0(\data_out_frame[20] [3]), .I1(n34478), 
            .I2(GND_net), .I3(GND_net), .O(n30907));
    defparam i1_2_lut_adj_905.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_906 (.I0(\data_out_frame[20] [6]), .I1(\data_out_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n32658));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n32384), .O(n32385));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i2_3_lut_adj_907 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_825), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n16267));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_907.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_908 (.I0(n17222), .I1(\data_in_frame[7] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n32590));
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32391), .I3(\FRAME_MATCHER.i [0]), .O(n32397));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_adj_909 (.I0(\data_out_frame[11] [2]), .I1(n18108), 
            .I2(n18067), .I3(GND_net), .O(n32617));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_909.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_910 (.I0(\data_out_frame[13] [6]), .I1(n17297), 
            .I2(n16793), .I3(\data_out_frame[11] [5]), .O(n33041));
    defparam i1_4_lut_adj_910.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_911 (.I0(n17886), .I1(n32993), .I2(\data_out_frame[9] [0]), 
            .I3(n32617), .O(n12_adj_3981));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_912 (.I0(n1169), .I1(n12_adj_3981), .I2(\data_out_frame[13] [4]), 
            .I3(n32854), .O(n32511));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_912.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_913 (.I0(n17664), .I1(\data_out_frame[18] [2]), 
            .I2(n32511), .I3(n33041), .O(n32782));
    defparam i3_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_914 (.I0(\data_out_frame[18] [3]), .I1(n32782), 
            .I2(n30803), .I3(\data_out_frame[16] [2]), .O(n33521));
    defparam i3_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_915 (.I0(n33836), .I1(n2063), .I2(GND_net), .I3(GND_net), 
            .O(n32722));
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_916 (.I0(\data_out_frame[20] [5]), .I1(n30867), 
            .I2(\data_out_frame[23] [0]), .I3(n32722), .O(n10_adj_3982));
    defparam i4_4_lut_adj_916.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_917 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [5]), .I3(GND_net), .O(n17610));
    defparam i2_3_lut_adj_917.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_918 (.I0(n17610), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[11] [3]), .I3(\data_out_frame[7] [1]), .O(n32993));
    defparam i3_4_lut_adj_918.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_919 (.I0(n32993), .I1(n32428), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3983));
    defparam i2_2_lut_adj_919.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_920 (.I0(\data_out_frame[13] [5]), .I1(\data_out_frame[9] [1]), 
            .I2(n6_adj_3983), .I3(n32802), .O(n29984));
    defparam i1_4_lut_adj_920.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_921 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(n29984), .I3(n32690), .O(n10_adj_3984));
    defparam i4_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n18754));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_922 (.I0(\data_out_frame[16] [1]), .I1(n32939), 
            .I2(n10_adj_3984), .I3(n16793), .O(n30024));
    defparam i1_4_lut_adj_922.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_923 (.I0(\data_out_frame[18] [4]), .I1(n30024), 
            .I2(\data_out_frame[16] [3]), .I3(n6_adj_3985), .O(n2063));
    defparam i4_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_924 (.I0(n2063), .I1(\data_out_frame[23] [2]), 
            .I2(\data_out_frame[23] [1]), .I3(GND_net), .O(n32671));
    defparam i2_3_lut_adj_924.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_925 (.I0(n15336), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [6]), .I3(n30867), .O(n32920));
    defparam i1_4_lut_adj_925.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_926 (.I0(n32920), .I1(\data_out_frame[25] [3]), 
            .I2(n32671), .I3(GND_net), .O(n32825));
    defparam i2_3_lut_adj_926.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_927 (.I0(\data_out_frame[16] [5]), .I1(n29969), 
            .I2(GND_net), .I3(GND_net), .O(n32556));
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_928 (.I0(\data_out_frame[16] [7]), .I1(n18032), 
            .I2(n29979), .I3(n17810), .O(n30798));
    defparam i3_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_929 (.I0(\data_out_frame[19] [1]), .I1(n30798), 
            .I2(GND_net), .I3(GND_net), .O(n30856));
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_930 (.I0(\data_out_frame[25] [4]), .I1(n32825), 
            .I2(n29938), .I3(GND_net), .O(n32687));
    defparam i2_3_lut_adj_930.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_931 (.I0(\data_out_frame[23] [3]), .I1(n30783), 
            .I2(n30856), .I3(n6_adj_3986), .O(n34449));
    defparam i4_4_lut_adj_931.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_932 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n18111));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_932.LUT_INIT = 16'h6666;
    SB_LUT4 i342_2_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1130));   // verilog/coms.v(76[16:27])
    defparam i342_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_out_frame[9] [3]), .I1(n17886), 
            .I2(GND_net), .I3(GND_net), .O(n32990));
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_934 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[14] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33054));
    defparam i1_2_lut_adj_934.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_935 (.I0(n32802), .I1(n32990), .I2(GND_net), 
            .I3(GND_net), .O(n17297));
    defparam i1_2_lut_adj_935.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_936 (.I0(n32939), .I1(n29949), .I2(n17297), .I3(n33054), 
            .O(n10_adj_3987));
    defparam i4_4_lut_adj_936.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32498));
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_938 (.I0(n15336), .I1(n29938), .I2(\data_out_frame[20] [6]), 
            .I3(GND_net), .O(n33836));
    defparam i2_3_lut_adj_938.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_939 (.I0(\data_out_frame[23] [2]), .I1(n33836), 
            .I2(GND_net), .I3(GND_net), .O(n30783));
    defparam i1_2_lut_adj_939.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_940 (.I0(\data_out_frame[25] [4]), .I1(\data_out_frame[25] [5]), 
            .I2(n30783), .I3(n30811), .O(n33862));
    defparam i3_4_lut_adj_940.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_941 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17354));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_942 (.I0(n30912), .I1(n29938), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n30811));
    defparam i2_3_lut_adj_942.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_943 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n32805));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_943.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_944 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[8] [0]), 
            .I2(n33072), .I3(n6_adj_3988), .O(n32443));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_944.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_945 (.I0(\data_out_frame[5] [3]), .I1(n32463), 
            .I2(n17098), .I3(n1191), .O(n1168));   // verilog/coms.v(71[16:62])
    defparam i3_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i381_2_lut (.I0(n1168), .I1(\data_out_frame[4] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n1169));   // verilog/coms.v(71[16:69])
    defparam i381_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_946 (.I0(\data_out_frame[9] [4]), .I1(n32596), 
            .I2(n32428), .I3(\data_out_frame[7] [1]), .O(n32885));
    defparam i3_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_947 (.I0(n32885), .I1(\data_out_frame[11] [7]), 
            .I2(\data_out_frame[13] [7]), .I3(n33027), .O(n10_adj_3989));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_948 (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n32746));
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_949 (.I0(\data_out_frame[16] [5]), .I1(\data_out_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17807));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_949.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_950 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[6] [0]), .I3(GND_net), .O(n33569));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_950.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_951 (.I0(n32443), .I1(n33569), .I2(n32996), .I3(n32805), 
            .O(n17207));   // verilog/coms.v(74[16:27])
    defparam i3_4_lut_adj_951.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_952 (.I0(n17207), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3990));
    defparam i1_2_lut_adj_952.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_953 (.I0(n17807), .I1(n29969), .I2(n29953), .I3(n6_adj_3990), 
            .O(n32699));
    defparam i4_4_lut_adj_953.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_954 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n32872));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_954.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33011));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17098));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_out_frame[4] [7]), .I1(n32438), 
            .I2(GND_net), .I3(GND_net), .O(n17883));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33072));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_959 (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[12] [1]), 
            .I2(\data_out_frame[11] [7]), .I3(GND_net), .O(n32814));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_959.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_960 (.I0(n32814), .I1(n32984), .I2(\data_out_frame[9] [5]), 
            .I3(n32460), .O(n12_adj_3991));   // verilog/coms.v(75[16:27])
    defparam i5_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_961 (.I0(\data_out_frame[9] [6]), .I1(n12_adj_3991), 
            .I2(n33072), .I3(n17883), .O(n29969));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_962 (.I0(n33011), .I1(\data_out_frame[9] [5]), 
            .I2(n32561), .I3(\data_out_frame[7] [6]), .O(n14_adj_3992));
    defparam i6_4_lut_adj_962.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_963 (.I0(\data_out_frame[12] [1]), .I1(n14_adj_3992), 
            .I2(n10_adj_3993), .I3(n32463), .O(n16700));
    defparam i7_4_lut_adj_963.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_964 (.I0(n16700), .I1(\data_out_frame[14] [2]), 
            .I2(n29969), .I3(GND_net), .O(n33517));
    defparam i2_3_lut_adj_964.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_965 (.I0(\data_out_frame[18] [7]), .I1(n17711), 
            .I2(n17207), .I3(GND_net), .O(n18032));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_965.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_966 (.I0(\data_out_frame[19] [0]), .I1(n18032), 
            .I2(n33517), .I3(\data_out_frame[16] [4]), .O(n10_adj_3994));
    defparam i4_4_lut_adj_966.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_967 (.I0(\data_out_frame[18] [6]), .I1(n10_adj_3994), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n29938));
    defparam i5_3_lut_adj_967.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\data_out_frame[18] [5]), .I1(n32699), 
            .I2(GND_net), .I3(GND_net), .O(n32945));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\data_out_frame[23] [4]), .I1(\data_out_frame[23] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17250));
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32546));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_971 (.I0(n17108), .I1(\data_out_frame[10] [6]), 
            .I2(\data_out_frame[13] [0]), .I3(n32860), .O(n16_adj_3995));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_972 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[10] [4]), 
            .I2(n33014), .I3(\data_out_frame[6] [0]), .O(n17_adj_3996));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_973 (.I0(n17_adj_3996), .I1(\data_out_frame[8] [5]), 
            .I2(n16_adj_3995), .I3(\data_out_frame[12] [6]), .O(n29940));   // verilog/coms.v(85[17:28])
    defparam i9_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_974 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32620));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_974.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_975 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32463));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_976 (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n32822));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_976.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_977 (.I0(n32822), .I1(\data_out_frame[8] [2]), 
            .I2(n17104), .I3(\data_out_frame[12] [4]), .O(n14_adj_3997));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_978 (.I0(n32999), .I1(n14_adj_3997), .I2(n10_adj_3998), 
            .I3(\data_out_frame[10] [4]), .O(n17810));   // verilog/coms.v(85[17:63])
    defparam i7_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33075));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_980 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n32817));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_980.LUT_INIT = 16'h6666;
    SB_LUT4 i375_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1191));   // verilog/coms.v(71[16:27])
    defparam i375_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_981 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n32460));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_981.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_982 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32996));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_982.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_983 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[4] [0]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n17104));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_983.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_out_frame[8] [4]), .I1(n17104), 
            .I2(GND_net), .I3(GND_net), .O(n32608));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1193));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_986 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n32984));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_986.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_987 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[12] [5]), 
            .I2(\data_out_frame[6] [2]), .I3(\data_out_frame[14] [7]), .O(n32785));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_988 (.I0(n32785), .I1(n32984), .I2(\data_out_frame[10] [5]), 
            .I3(n1193), .O(n15_adj_3999));   // verilog/coms.v(73[16:42])
    defparam i6_4_lut_adj_988.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_989 (.I0(n15_adj_3999), .I1(\data_out_frame[12] [6]), 
            .I2(n14_adj_4000), .I3(n17678), .O(n29901));   // verilog/coms.v(73[16:42])
    defparam i8_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_990 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[14] [5]), 
            .I2(n32996), .I3(n32460), .O(n16_adj_4001));   // verilog/coms.v(75[16:27])
    defparam i6_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_991 (.I0(\data_out_frame[8] [2]), .I1(n32817), 
            .I2(n33075), .I3(\data_out_frame[4] [0]), .O(n17_adj_4002));   // verilog/coms.v(75[16:27])
    defparam i7_4_lut_adj_991.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_992 (.I0(n17_adj_4002), .I1(\data_out_frame[10] [3]), 
            .I2(n16_adj_4001), .I3(\data_out_frame[12] [4]), .O(n17711));   // verilog/coms.v(75[16:27])
    defparam i9_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_993 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4003));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_994 (.I0(\data_out_frame[15] [0]), .I1(n17711), 
            .I2(n29901), .I3(n6_adj_4003), .O(n32425));
    defparam i4_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_995 (.I0(\data_out_frame[17] [2]), .I1(n17810), 
            .I2(n32620), .I3(n29940), .O(n32788));   // verilog/coms.v(71[16:62])
    defparam i3_4_lut_adj_995.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_996 (.I0(n32788), .I1(\data_out_frame[19] [3]), 
            .I2(n32425), .I3(GND_net), .O(n29870));
    defparam i2_3_lut_adj_996.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut (.I0(n17810), .I1(\data_out_frame[17] [0]), .I2(n32425), 
            .I3(GND_net), .O(n8_adj_4004));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_997 (.I0(\data_out_frame[19] [2]), .I1(n17354), 
            .I2(n8_adj_4004), .I3(n17207), .O(n30912));
    defparam i1_4_lut_adj_997.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_998 (.I0(n30912), .I1(n29870), .I2(GND_net), 
            .I3(GND_net), .O(n30788));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_999 (.I0(\data_out_frame[25] [5]), .I1(n32975), 
            .I2(GND_net), .I3(GND_net), .O(n32936));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h6666;
    SB_LUT4 i22_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4005));   // verilog/coms.v(127[12] 300[6])
    defparam i22_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1000 (.I0(n24776), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n8_adj_4005), .I3(\FRAME_MATCHER.state [2]), .O(n32378));
    defparam i3_4_lut_adj_1000.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\FRAME_MATCHER.state [1]), .I1(n32378), 
            .I2(GND_net), .I3(GND_net), .O(n18277));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h4444;
    SB_LUT4 i3_4_lut_adj_1002 (.I0(n30867), .I1(n32936), .I2(n32737), 
            .I3(n30788), .O(n33621));
    defparam i3_4_lut_adj_1002.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1003 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32398), .I3(\FRAME_MATCHER.i [0]), .O(n32403));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1003.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_1004 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(n32491), .I3(n6_adj_4006), .O(Kp_23__N_806));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1004.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1005 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_806), 
            .I2(GND_net), .I3(GND_net), .O(n32478));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_1005.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1006 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[1] [5]), 
            .I2(n32478), .I3(\data_in_frame[1] [4]), .O(n26));
    defparam i9_4_lut_adj_1006.LUT_INIT = 16'h8400;
    SB_LUT4 i12_4_lut_adj_1007 (.I0(n17177), .I1(n24), .I2(Kp_23__N_806), 
            .I3(\data_in_frame[2] [1]), .O(n29_adj_4007));
    defparam i12_4_lut_adj_1007.LUT_INIT = 16'h0440;
    SB_LUT4 i4_4_lut_adj_1008 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [1]), .I3(n32478), .O(n21));
    defparam i4_4_lut_adj_1008.LUT_INIT = 16'h2184;
    SB_LUT4 i15_4_lut_adj_1009 (.I0(n29_adj_4007), .I1(n4_c), .I2(n26), 
            .I3(n14565), .O(n32_adj_4008));
    defparam i15_4_lut_adj_1009.LUT_INIT = 16'h0020;
    SB_LUT4 i10_4_lut_adj_1010 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [6]), .I3(n32505), .O(n27));
    defparam i10_4_lut_adj_1010.LUT_INIT = 16'h0080;
    SB_LUT4 i16_4_lut_adj_1011 (.I0(n27), .I1(n32_adj_4008), .I2(n21), 
            .I3(n34988), .O(\FRAME_MATCHER.state_31__N_2561 [3]));
    defparam i16_4_lut_adj_1011.LUT_INIT = 16'h0080;
    SB_LUT4 i1_4_lut_adj_1012 (.I0(\FRAME_MATCHER.state [3]), .I1(n4_adj_4009), 
            .I2(n2_adj_4010), .I3(n1_c), .O(n5));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1012.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_4_lut_adj_1013 (.I0(n17092), .I1(n5), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state_31__N_2561 [3]), .O(n31898));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'hcdcc;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1014 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32406), .I3(\FRAME_MATCHER.i [0]), .O(n32412));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1014.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\FRAME_MATCHER.state [4]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31890));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1016 (.I0(\FRAME_MATCHER.state [5]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31888));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(\FRAME_MATCHER.state [6]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31832));
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\FRAME_MATCHER.state [7]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31834));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(\FRAME_MATCHER.state [8]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31886));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1020 (.I0(\FRAME_MATCHER.state [9]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31884));
    defparam i1_2_lut_adj_1020.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(\FRAME_MATCHER.state [10]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31882));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(\FRAME_MATCHER.state [11]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31880));
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\FRAME_MATCHER.state [12]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31878));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1024 (.I0(\FRAME_MATCHER.state [13]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31876));
    defparam i1_2_lut_adj_1024.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1025 (.I0(\FRAME_MATCHER.state [14]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31874));
    defparam i1_2_lut_adj_1025.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\FRAME_MATCHER.state [15]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31836));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\FRAME_MATCHER.state [16]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31838));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\FRAME_MATCHER.state [17]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31820));
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\FRAME_MATCHER.state [18]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31872));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\FRAME_MATCHER.state [19]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31870));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\FRAME_MATCHER.state [20]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31868));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n18753));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\FRAME_MATCHER.state [21]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31866));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1033 (.I0(\FRAME_MATCHER.state [22]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4012));
    defparam i1_2_lut_adj_1033.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1034 (.I0(\FRAME_MATCHER.state [23]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4013));
    defparam i1_2_lut_adj_1034.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\FRAME_MATCHER.state [24]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31864));
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(\FRAME_MATCHER.state [25]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31862));
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1037 (.I0(\FRAME_MATCHER.state [26]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31860));
    defparam i1_2_lut_adj_1037.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1038 (.I0(\FRAME_MATCHER.state [27]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31892));
    defparam i1_2_lut_adj_1038.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(\FRAME_MATCHER.state [28]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n31858));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(\FRAME_MATCHER.state [29]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4014));
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(\FRAME_MATCHER.state [30]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4015));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(\FRAME_MATCHER.state[0] ), .I1(n66), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2463 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\FRAME_MATCHER.state [31]), .I1(n5_adj_4011), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4016));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n18752));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(n17483), .I1(n32728), .I2(n32725), .I3(n29870), 
            .O(n30287));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n18751));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n18750));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n18749));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1044 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [7]), 
            .I2(n32452), .I3(n6_adj_4017), .O(Kp_23__N_825));   // verilog/coms.v(73[16:34])
    defparam i4_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1045 (.I0(n32766), .I1(n10_adj_4018), .I2(\data_in_frame[16] [6]), 
            .I3(GND_net), .O(n30504));
    defparam i5_3_lut_adj_1045.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(n17198), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[13] [5]), .I3(n30884), .O(n33063));
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'h9669;
    SB_LUT4 i19_4_lut_adj_1047 (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[17] [4]), 
            .I2(\data_in_frame[13] [2]), .I3(\data_in_frame[14] [3]), .O(n46_adj_4019));
    defparam i19_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1048 (.I0(n32655), .I1(n32794), .I2(\data_in_frame[13] [7]), 
            .I3(n32455), .O(n42_adj_4020));
    defparam i15_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n27756), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i12_4_lut_adj_1049 (.I0(n32757), .I1(n17187), .I2(\data_in_frame[10] [2]), 
            .I3(\data_in_frame[11] [2]), .O(n28_adj_4021));
    defparam i12_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1050 (.I0(\data_in_frame[11] [0]), .I1(n33084), 
            .I2(n32494), .I3(n32927), .O(n26_adj_4022));
    defparam i10_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1051 (.I0(n17427), .I1(n33081), .I2(n17447), 
            .I3(n32933), .O(n27_adj_4023));
    defparam i11_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1052 (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(n34667), .I3(n33050), .O(n25));
    defparam i9_4_lut_adj_1052.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1053 (.I0(n25), .I1(n27_adj_4023), .I2(n26_adj_4022), 
            .I3(n28_adj_4021), .O(n34390));
    defparam i15_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1054 (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[18] [1]), 
            .I2(\data_in_frame[16] [1]), .I3(Kp_23__N_1335), .O(n34));
    defparam i7_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1055 (.I0(n34390), .I1(n32888), .I2(n30314), 
            .I3(n33005), .O(n43_adj_4024));
    defparam i16_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1056 (.I0(n32501), .I1(n46_adj_4019), .I2(n36), 
            .I3(n32650), .O(n50));
    defparam i23_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1057 (.I0(n33069), .I1(n42_adj_4020), .I2(n33066), 
            .I3(\data_in_frame[10] [5]), .O(n48_adj_4025));
    defparam i21_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1058 (.I0(n43_adj_4024), .I1(n32828), .I2(n34), 
            .I3(n32763), .O(n49_adj_4026));
    defparam i22_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1059 (.I0(\data_in_frame[15] [5]), .I1(n17758), 
            .I2(\data_in_frame[18] [3]), .I3(\data_in_frame[18] [7]), .O(n47_adj_4027));
    defparam i20_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i26_4_lut_adj_1060 (.I0(n47_adj_4027), .I1(n49_adj_4026), .I2(n48_adj_4025), 
            .I3(n50), .O(n17579));
    defparam i26_4_lut_adj_1060.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[19] [6]), .I3(\data_in_frame[19] [2]), .O(n6_adj_4028));   // verilog/coms.v(85[17:28])
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1061 (.I0(\data_in_frame[19] [1]), .I1(n6_adj_4028), 
            .I2(\data_in_frame[19] [4]), .I3(\data_in_frame[19] [5]), .O(Kp_23__N_698));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1062 (.I0(n30314), .I1(Kp_23__N_698), .I2(n32791), 
            .I3(n17579), .O(n32905));
    defparam i2_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1063 (.I0(\data_in_frame[11] [1]), .I1(n5_adj_4029), 
            .I2(n32611), .I3(n32693), .O(n12_adj_4030));
    defparam i5_4_lut_adj_1063.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1064 (.I0(\data_in_frame[10] [6]), .I1(n12_adj_4030), 
            .I2(\data_in_frame[15] [4]), .I3(n32942), .O(n34750));
    defparam i6_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4031));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1066 (.I0(n33060), .I1(n30809), .I2(\data_in_frame[15] [6]), 
            .I3(n6_adj_4031), .O(n32791));
    defparam i4_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1067 (.I0(n32743), .I1(n32957), .I2(\data_in_frame[17] [5]), 
            .I3(\data_in_frame[13] [1]), .O(n10_adj_4032));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1067.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1068 (.I0(n34750), .I1(n10_adj_4032), .I2(\data_in_frame[10] [6]), 
            .I3(GND_net), .O(n30314));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1068.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4033));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1070 (.I0(\data_in_frame[18] [5]), .I1(n5_adj_4033), 
            .I2(n32714), .I3(n34722), .O(n32987));
    defparam i1_4_lut_adj_1070.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1071 (.I0(\data_in_frame[14] [0]), .I1(n30884), 
            .I2(Kp_23__N_1170), .I3(n6_adj_4034), .O(n32963));
    defparam i4_4_lut_adj_1071.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1072 (.I0(n32987), .I1(n33047), .I2(\data_in_frame[16] [2]), 
            .I3(GND_net), .O(n32455));
    defparam i2_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_in_frame[10] [1]), .I1(n29843), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4035));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1074 (.I0(\data_in_frame[12] [1]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[11] [7]), .I3(n6_adj_4035), .O(n32757));
    defparam i4_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1075 (.I0(\data_in_frame[12] [2]), .I1(n32966), 
            .I2(n15471), .I3(\data_in_frame[9] [6]), .O(n12_adj_4036));
    defparam i5_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1076 (.I0(\data_in_frame[9] [5]), .I1(n12_adj_4036), 
            .I2(\data_in_frame[14] [3]), .I3(n32757), .O(n34722));
    defparam i6_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1077 (.I0(n30921), .I1(\data_in_frame[14] [5]), 
            .I2(n34722), .I3(\data_in_frame[10] [3]), .O(n10_adj_4037));
    defparam i4_4_lut_adj_1077.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1078 (.I0(\data_in_frame[14] [4]), .I1(n15478), 
            .I2(n10_adj_4037), .I3(\data_in_frame[12] [4]), .O(n32766));
    defparam i1_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1079 (.I0(\data_in_frame[16] [7]), .I1(n32972), 
            .I2(n32766), .I3(\data_in_frame[16] [5]), .O(n32763));
    defparam i3_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(\data_in_frame[10] [3]), .I1(n18035), 
            .I2(GND_net), .I3(GND_net), .O(n17187));
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1351_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n5063), .I3(GND_net), .O(n5087));
    defparam mux_1351_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1081 (.I0(n17187), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[17] [3]), .I3(\data_in_frame[14] [7]), .O(n33005));
    defparam i3_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1351_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n5063), .I3(GND_net), .O(n5086));
    defparam mux_1351_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n5063), .I3(GND_net), .O(n5085));
    defparam mux_1351_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1082 (.I0(n32834), .I1(\data_in_frame[13] [1]), 
            .I2(\data_in_frame[12] [6]), .I3(n33005), .O(n10_adj_4038));
    defparam i4_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1083 (.I0(n32611), .I1(n10_adj_4038), .I2(n15478), 
            .I3(GND_net), .O(n17842));
    defparam i5_3_lut_adj_1083.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1373));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1084 (.I0(n32760), .I1(\data_in_frame[9] [1]), 
            .I2(n30777), .I3(n29856), .O(n12_adj_4039));
    defparam i5_4_lut_adj_1084.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1085 (.I0(\data_in_frame[11] [1]), .I1(n12_adj_4039), 
            .I2(n33033), .I3(n29843), .O(n34667));
    defparam i6_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(n34667), .I1(\data_in_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32693));
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h9999;
    SB_LUT4 mux_1351_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n5063), .I3(GND_net), .O(n5084));
    defparam mux_1351_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n5063), .I3(GND_net), .O(n5083));
    defparam mux_1351_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n5063), .I3(GND_net), .O(n5082));
    defparam mux_1351_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1087 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[9] [2]), 
            .I2(n30005), .I3(n6_adj_4040), .O(n30809));
    defparam i4_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1088 (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[15] [5]), 
            .I2(n32731), .I3(\data_in_frame[17] [7]), .O(n10_adj_4041));
    defparam i4_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1089 (.I0(n30809), .I1(n10_adj_4041), .I2(n17434), 
            .I3(n32693), .O(n30823));
    defparam i5_4_lut_adj_1089.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1090 (.I0(Kp_23__N_1032), .I1(n32650), .I2(GND_net), 
            .I3(GND_net), .O(n17705));
    defparam i1_2_lut_adj_1090.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1351_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n5063), .I3(GND_net), .O(n5081));
    defparam mux_1351_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n5063), .I3(GND_net), .O(n5080));
    defparam mux_1351_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n5063), .I3(GND_net), .O(n5079));
    defparam mux_1351_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1091 (.I0(\data_in_frame[13] [4]), .I1(n33033), 
            .I2(\data_in_frame[11] [3]), .I3(GND_net), .O(n32614));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1091.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1351_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n5063), .I3(GND_net), .O(n5078));
    defparam mux_1351_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1092 (.I0(\data_in_frame[13] [5]), .I1(n32933), 
            .I2(GND_net), .I3(GND_net), .O(n32655));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1351_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n5063), .I3(GND_net), .O(n5077));
    defparam mux_1351_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n5063), .I3(GND_net), .O(n5076));
    defparam mux_1351_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1093 (.I0(n17434), .I1(\data_in_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n33060));
    defparam i1_2_lut_adj_1093.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1094 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[5] [3]), .I3(GND_net), .O(n32577));
    defparam i2_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1351_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n5063), .I3(GND_net), .O(n5075));
    defparam mux_1351_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(n29843), .I1(n17814), .I2(GND_net), 
            .I3(GND_net), .O(n29856));
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1096 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17128));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h6666;
    SB_LUT4 i4_3_lut (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n12_adj_4042));   // verilog/coms.v(85[17:28])
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1351_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n5063), .I3(GND_net), .O(n5074));
    defparam mux_1351_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1097 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[9] [6]), 
            .I2(n30259), .I3(n33438), .O(n13));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_1097.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1098 (.I0(n13), .I1(n17128), .I2(n12_adj_4042), 
            .I3(n32623), .O(n33084));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1351_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n5063), .I3(GND_net), .O(n5073));
    defparam mux_1351_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n5063), .I3(GND_net), .O(n5072));
    defparam mux_1351_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1099 (.I0(\data_in_frame[9] [1]), .I1(n17364), 
            .I2(GND_net), .I3(GND_net), .O(n32647));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1099.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1100 (.I0(n32845), .I1(n32647), .I2(\data_in_frame[9] [0]), 
            .I3(\data_in_frame[8] [2]), .O(n18));   // verilog/coms.v(70[16:69])
    defparam i7_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1101 (.I0(n17396), .I1(n18), .I2(\data_in_frame[6] [3]), 
            .I3(n33084), .O(n20));   // verilog/coms.v(70[16:69])
    defparam i9_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1102 (.I0(n33008), .I1(n20), .I2(n16_adj_4043), 
            .I3(n32677), .O(n32775));   // verilog/coms.v(70[16:69])
    defparam i10_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n27755), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1103 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17342));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1104 (.I0(n17342), .I1(n32775), .I2(\data_in_frame[11] [7]), 
            .I3(n32645), .O(n12_adj_4044));
    defparam i5_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1105 (.I0(\data_in_frame[9] [2]), .I1(n12_adj_4044), 
            .I2(\data_in_frame[14] [1]), .I3(n29856), .O(n32714));
    defparam i6_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1351_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n5063), .I3(GND_net), .O(n5071));
    defparam mux_1351_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1106 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[5] [0]), 
            .I2(n17177), .I3(\data_in_frame[9] [6]), .O(n28_adj_4045));
    defparam i12_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1351_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n5063), .I3(GND_net), .O(n5070));
    defparam mux_1351_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1107 (.I0(n33017), .I1(n30259), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[3] [0]), .O(n26_adj_4046));
    defparam i10_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1108 (.I0(n33024), .I1(n32577), .I2(n32863), 
            .I3(\data_in_frame[12] [1]), .O(n27_adj_4047));
    defparam i11_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1109 (.I0(n30001), .I1(n32775), .I2(\data_in_frame[11] [6]), 
            .I3(n17128), .O(n25_adj_4048));
    defparam i9_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1351_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n5063), .I3(GND_net), .O(n5069));
    defparam mux_1351_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15_4_lut_adj_1110 (.I0(n25_adj_4048), .I1(n27_adj_4047), .I2(n26_adj_4046), 
            .I3(n28_adj_4045), .O(n34613));
    defparam i15_4_lut_adj_1110.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1111 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32683));
    defparam i1_2_lut_adj_1111.LUT_INIT = 16'h6666;
    SB_LUT4 mux_1351_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n5063), .I3(GND_net), .O(n5068));
    defparam mux_1351_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n5063), .I3(GND_net), .O(n5067));
    defparam mux_1351_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1351_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n5063), .I3(GND_net), .O(n5066));
    defparam mux_1351_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1112 (.I0(\data_in_frame[18] [4]), .I1(n34613), 
            .I2(n32714), .I3(\data_in_frame[14] [2]), .O(n33047));
    defparam i1_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1113 (.I0(\data_in_frame[18] [3]), .I1(n30005), 
            .I2(\data_in_frame[15] [7]), .I3(n17342), .O(n32930));
    defparam i3_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[8] [0]), .I1(n17358), 
            .I2(GND_net), .I3(GND_net), .O(n32966));
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1115 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[12] [3]), 
            .I2(\data_in_frame[9] [7]), .I3(n6_adj_4049), .O(n32794));
    defparam i4_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(n15471), .I1(n32794), .I2(GND_net), 
            .I3(GND_net), .O(n30921));
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[16] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n32888));
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n33081));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1119 (.I0(n17246), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[14] [6]), .I3(n6_adj_4050), .O(n32501));
    defparam i4_4_lut_adj_1119.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n32623));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1121 (.I0(n17316), .I1(\data_in_frame[10] [2]), 
            .I2(n32590), .I3(n17867), .O(n16_adj_4051));
    defparam i6_4_lut_adj_1121.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1122 (.I0(n30028), .I1(\data_in_frame[1] [2]), 
            .I2(n32880), .I3(n17745), .O(n17_adj_4052));
    defparam i7_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1123 (.I0(n17_adj_4052), .I1(n29907), .I2(n16_adj_4051), 
            .I3(\data_in_frame[3] [4]), .O(n29854));
    defparam i9_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1124 (.I0(\data_in_frame[12] [2]), .I1(n30001), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n33050));
    defparam i2_3_lut_adj_1124.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1125 (.I0(\data_in_frame[17] [0]), .I1(n32571), 
            .I2(n4_adj_4053), .I3(\data_in_frame[14] [6]), .O(n10_adj_4054));
    defparam i4_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[8] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17396));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1127 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n32834));
    defparam i2_3_lut_adj_1127.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1128 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17447));
    defparam i1_2_lut_adj_1128.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1129 (.I0(n17212), .I1(\data_in_frame[14] [5]), 
            .I2(n17370), .I3(n33002), .O(n10_adj_4055));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1130 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[16] [7]), 
            .I2(n32602), .I3(n17447), .O(n32475));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1131 (.I0(n32834), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[17] [2]), .I3(n33002), .O(n10_adj_4056));
    defparam i4_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n18748));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19048_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_c), .I2(n63_adj_4057), 
            .I3(GND_net), .O(n92[2]));   // verilog/coms.v(139[4] 141[7])
    defparam i19048_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i19038_rep_320_2_lut (.I0(n92[2]), .I1(n63), .I2(GND_net), 
            .I3(GND_net), .O(n38282));   // verilog/coms.v(142[4] 144[7])
    defparam i19038_rep_320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_3_lut_adj_1132 (.I0(n32501), .I1(n10_adj_4056), .I2(n29854), 
            .I3(GND_net), .O(n30543));
    defparam i5_3_lut_adj_1132.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1133 (.I0(n32972), .I1(n32602), .I2(\data_in_frame[14] [4]), 
            .I3(n33050), .O(n10_adj_4059));
    defparam i4_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 select_441_Select_2_i5_4_lut (.I0(n92[2]), .I1(\FRAME_MATCHER.i_31__N_2461 ), 
            .I2(n3303), .I3(n63), .O(n5_adj_4060));
    defparam select_441_Select_2_i5_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i1_2_lut_adj_1134 (.I0(n17364), .I1(n10_adj_4061), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1167));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1135 (.I0(n10_adj_4061), .I1(n17814), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1170));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1136 (.I0(\data_in_frame[9] [0]), .I1(n30777), 
            .I2(n18035), .I3(GND_net), .O(n33438));
    defparam i2_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1137 (.I0(n17745), .I1(\data_in_frame[7] [7]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n32677));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1137.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1138 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17316));
    defparam i1_2_lut_adj_1138.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1139 (.I0(\FRAME_MATCHER.i_31__N_2463 ), .I1(n92[2]), 
            .I2(n4452), .I3(n63), .O(n1_adj_4062));   // verilog/coms.v(201[5:24])
    defparam i1_4_lut_adj_1139.LUT_INIT = 16'ha8a0;
    SB_LUT4 i3_4_lut_adj_1140 (.I0(n1_adj_4062), .I1(n5_adj_4060), .I2(n38282), 
            .I3(n33978), .O(n8_adj_4063));   // verilog/coms.v(201[5:24])
    defparam i3_4_lut_adj_1140.LUT_INIT = 16'heefe;
    SB_LUT4 i4_4_lut_adj_1141 (.I0(n92[2]), .I1(n8_adj_4063), .I2(n34405), 
            .I3(n5_adj_4064), .O(n37935));   // verilog/coms.v(201[5:24])
    defparam i4_4_lut_adj_1141.LUT_INIT = 16'hefcf;
    SB_LUT4 i4_4_lut_adj_1142 (.I0(n17589), .I1(n17926), .I2(n32577), 
            .I3(n6_adj_4065), .O(n17418));
    defparam i4_4_lut_adj_1142.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(n29843), .I1(n17418), .I2(GND_net), 
            .I3(GND_net), .O(n29850));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1144 (.I0(n32667), .I1(n33008), .I2(n17427), 
            .I3(n17246), .O(n12_adj_4066));
    defparam i5_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1145 (.I0(n29850), .I1(n12_adj_4066), .I2(n5_adj_4029), 
            .I3(n29907), .O(n32917));
    defparam i6_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1146 (.I0(n33438), .I1(Kp_23__N_1170), .I2(\data_in_frame[10] [7]), 
            .I3(GND_net), .O(n32760));
    defparam i2_3_lut_adj_1146.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17758));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n33066));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1149 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n32957));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1149.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1150 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17212));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1151 (.I0(\data_in_frame[13] [2]), .I1(n17364), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4067));
    defparam i1_2_lut_adj_1151.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1152 (.I0(n32760), .I1(n8_adj_4068), .I2(n32917), 
            .I3(n6_adj_4067), .O(n32942));
    defparam i4_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1153 (.I0(n17246), .I1(n32942), .I2(\data_in_frame[15] [3]), 
            .I3(GND_net), .O(n32743));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1153.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_17__7__I_0_3899_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1335));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_17__7__I_0_3899_2_lut.LUT_INIT = 16'h6666;
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3453[0]), .C(clk32MHz), 
            .D(n3519[0]), .R(n3482));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1154 (.I0(n32960), .I1(n17212), .I2(n32494), 
            .I3(\data_in_frame[15] [2]), .O(n14_adj_4069));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1155 (.I0(\data_in_frame[17] [4]), .I1(n14_adj_4069), 
            .I2(n10_adj_4070), .I3(\data_in_frame[13] [0]), .O(n17699));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_1155.LUT_INIT = 16'h6996;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
            .D(n31814), .S(n33985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n18744));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1156 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17867));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1156.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n18216), .D(n8825[7]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_rep_69_3_lut (.I0(n30854), .I1(n30543), .I2(n32475), .I3(GND_net), 
            .O(n38031));
    defparam i1_rep_69_3_lut.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n18216), .D(n8825[6]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1157 (.I0(n32930), .I1(n33047), .I2(\data_in_frame[20] [5]), 
            .I3(n32683), .O(n12_adj_4071));
    defparam i5_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1158 (.I0(\data_in_frame[15] [6]), .I1(n8_adj_4072), 
            .I2(\data_in_frame[20] [2]), .I3(n30823), .O(n10_adj_4073));
    defparam i4_4_lut_adj_1158.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n18743));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1159 (.I0(\data_in_frame[16] [3]), .I1(n32455), 
            .I2(n32963), .I3(\data_in_frame[20] [6]), .O(n10_adj_4074));
    defparam i4_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1160 (.I0(\data_in_frame[20] [1]), .I1(n30314), 
            .I2(n32791), .I3(GND_net), .O(n6_adj_4075));
    defparam i2_3_lut_adj_1160.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1161 (.I0(n32709), .I1(n17699), .I2(n30543), 
            .I3(GND_net), .O(n10_adj_4076));
    defparam i3_3_lut_adj_1161.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1162 (.I0(n30543), .I1(n10_adj_4076), .I2(n30854), 
            .I3(n32475), .O(n12_adj_4077));
    defparam i5_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1163 (.I0(\data_in_frame[21] [1]), .I1(n32905), 
            .I2(n30314), .I3(n17699), .O(n11));
    defparam i4_4_lut_adj_1163.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1164 (.I0(\data_in_frame[21] [5]), .I1(\data_in_frame[19] [4]), 
            .I2(\data_in_frame[19] [3]), .I3(n6_adj_4078), .O(n34561));
    defparam i4_4_lut_adj_1164.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1165 (.I0(n30823), .I1(n34494), .I2(n6_adj_4075), 
            .I3(\data_in_frame[19] [7]), .O(n19));
    defparam i3_4_lut_adj_1165.LUT_INIT = 16'hb77b;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4079));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4080));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29850_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35893));
    defparam i29850_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29852_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35892));
    defparam i29852_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[18] [2]), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n10_adj_4081));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_adj_1166 (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[15] [6]), 
            .I2(n30823), .I3(GND_net), .O(n12_adj_4082));
    defparam i3_3_lut_adj_1166.LUT_INIT = 16'h6969;
    SB_LUT4 i7_4_lut_adj_1167 (.I0(Kp_23__N_1373), .I1(\data_in_frame[18] [1]), 
            .I2(n17705), .I3(n10_adj_4081), .O(n16_adj_4083));
    defparam i7_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1168 (.I0(n33063), .I1(n16_adj_4083), .I2(n12_adj_4082), 
            .I3(\data_in_frame[16] [0]), .O(n34814));
    defparam i8_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1169 (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[19] [2]), 
            .I2(n32709), .I3(GND_net), .O(n8_adj_4084));
    defparam i3_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_1170 (.I0(\data_in_frame[19] [3]), .I1(n38031), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[21] [4]), .O(n33574));
    defparam i2_4_lut_adj_1170.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_1__4__I_0_2_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_901));   // verilog/coms.v(75[16:27])
    defparam data_in_frame_1__4__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_rep_78_2_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n38040));
    defparam i1_rep_78_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1171 (.I0(n32963), .I1(\data_in_frame[16] [0]), 
            .I2(n32614), .I3(\data_in_frame[18] [2]), .O(n14_adj_4085));
    defparam i6_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1172 (.I0(\data_in_frame[20] [4]), .I1(n32930), 
            .I2(\data_in_frame[16] [2]), .I3(\data_in_frame[15] [6]), .O(n13_adj_4086));
    defparam i5_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n18241), .D(n5064));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_4_lut_adj_1173 (.I0(n17699), .I1(n38040), .I2(n30543), 
            .I3(\data_in_frame[21] [6]), .O(n34784));
    defparam i2_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1174 (.I0(\data_in_frame[21] [3]), .I1(n33574), 
            .I2(n8_adj_4084), .I3(n30854), .O(n23));
    defparam i7_4_lut_adj_1174.LUT_INIT = 16'hedde;
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n18742));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1175 (.I0(n13_adj_4087), .I1(n30823), .I2(n34750), 
            .I3(\data_in_frame[16] [0]), .O(n16_adj_4088));
    defparam i7_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1176 (.I0(\data_in_frame[19] [7]), .I1(n30809), 
            .I2(\data_in_frame[19] [6]), .I3(GND_net), .O(n11_adj_4089));
    defparam i2_3_lut_adj_1176.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1177 (.I0(n32791), .I1(\data_in_frame[19] [0]), 
            .I2(Kp_23__N_698), .I3(n32987), .O(n10_adj_4090));
    defparam i4_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_23_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n27717), .O(n2_adj_4091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i8_4_lut_adj_1178 (.I0(n11_adj_4089), .I1(n16_adj_4088), .I2(\data_in_frame[20] [0]), 
            .I3(n32731), .O(n34764));
    defparam i8_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n18741));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1179 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4092));
    defparam i1_2_lut_adj_1179.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1180 (.I0(n38031), .I1(n30314), .I2(\data_in_frame[21] [0]), 
            .I3(n32905), .O(n10_adj_4093));
    defparam i4_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1181 (.I0(\data_in_frame[21] [7]), .I1(n30314), 
            .I2(n17842), .I3(n6_adj_4092), .O(n33866));
    defparam i4_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1182 (.I0(\data_in_frame[16] [3]), .I1(n12_adj_4071), 
            .I2(n33063), .I3(\data_in_frame[16] [1]), .O(n34823));
    defparam i6_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1351_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n5063), .I3(GND_net), .O(n5065));
    defparam mux_1351_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1183 (.I0(\data_in_frame[18] [1]), .I1(n10_adj_4073), 
            .I2(n34750), .I3(Kp_23__N_1335), .O(n34774));
    defparam i5_4_lut_adj_1183.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1184 (.I0(n19), .I1(n34561), .I2(n11), .I3(n12_adj_4077), 
            .O(n26_adj_4094));
    defparam i10_4_lut_adj_1184.LUT_INIT = 16'hbffb;
    SB_LUT4 i3_4_lut_adj_1185 (.I0(n17867), .I1(n32808), .I2(n32452), 
            .I3(\data_in_frame[5] [7]), .O(n17358));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1186 (.I0(n30543), .I1(n33866), .I2(n10_adj_4093), 
            .I3(n30504), .O(n17_adj_4095));
    defparam i1_4_lut_adj_1186.LUT_INIT = 16'hb77b;
    SB_CARRY add_43_23 (.CI(n27717), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n27718));
    SB_LUT4 i6_4_lut_adj_1187 (.I0(n34814), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[21] [2]), .I3(n30504), .O(n22));
    defparam i6_4_lut_adj_1187.LUT_INIT = 16'hebbe;
    SB_LUT4 i12_4_lut_adj_1188 (.I0(n23), .I1(n34784), .I2(n13_adj_4086), 
            .I3(n14_adj_4085), .O(n28_adj_4096));
    defparam i12_4_lut_adj_1188.LUT_INIT = 16'hfbbf;
    SB_LUT4 i5_4_lut_adj_1189 (.I0(n34764), .I1(n17579), .I2(n10_adj_4090), 
            .I3(\data_in_frame[20] [7]), .O(n21_adj_4097));
    defparam i5_4_lut_adj_1189.LUT_INIT = 16'hebbe;
    SB_LUT4 i3_4_lut_adj_1190 (.I0(\data_in_frame[1] [3]), .I1(n32677), 
            .I2(n17867), .I3(n17768), .O(n15471));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_1190.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1191 (.I0(n17_adj_4095), .I1(n26_adj_4094), .I2(n34774), 
            .I3(n34823), .O(n29_adj_4098));
    defparam i13_4_lut_adj_1191.LUT_INIT = 16'hffef;
    SB_CARRY add_3971_8 (.CI(n27755), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n27756));
    SB_LUT4 i15_4_lut_adj_1192 (.I0(n29_adj_4098), .I1(n21_adj_4097), .I2(n28_adj_4096), 
            .I3(n22), .O(n31_adj_4099));
    defparam i15_4_lut_adj_1192.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(n17358), .I1(\data_in_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4053));   // verilog/coms.v(236[9:81])
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'h6666;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n27754), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1194 (.I0(\data_in_frame[6] [1]), .I1(n17768), 
            .I2(Kp_23__N_901), .I3(n6_adj_4100), .O(n17370));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1195 (.I0(\data_in_frame[8] [3]), .I1(n32487), 
            .I2(GND_net), .I3(GND_net), .O(n32828));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1195.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4101));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1197 (.I0(n17483), .I1(n32728), .I2(n32900), 
            .I3(n30895), .O(n33036));
    defparam i2_3_lut_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1198 (.I0(n32638), .I1(n17376), .I2(n32866), 
            .I3(n6_adj_4101), .O(n8_adj_4068));   // verilog/coms.v(77[16:43])
    defparam i4_4_lut_adj_1198.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1199 (.I0(n17589), .I1(\data_in_frame[0] [7]), 
            .I2(Kp_23__N_825), .I3(GND_net), .O(n17590));   // verilog/coms.v(71[16:69])
    defparam i2_3_lut_adj_1199.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1200 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[4] [1]), 
            .I2(n32848), .I3(\data_in_frame[1] [7]), .O(n32487));   // verilog/coms.v(78[16:27])
    defparam i3_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_7 (.CI(n27754), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n27755));
    SB_LUT4 i3_4_lut_adj_1201 (.I0(\data_in_frame[5] [2]), .I1(n32863), 
            .I2(n17590), .I3(\data_in_frame[4] [7]), .O(n29843));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_1201.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1202 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[5] [4]), 
            .I2(n17742), .I3(n6_adj_4102), .O(n30259));
    defparam i4_4_lut_adj_1202.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_in_frame[5] [1]), .I1(n32877), 
            .I2(GND_net), .I3(GND_net), .O(n32567));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1204 (.I0(\data_in_frame[2] [7]), .I1(n32567), 
            .I2(\data_in_frame[7] [2]), .I3(n16267), .O(n12_adj_4103));
    defparam i5_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1205 (.I0(\data_in_frame[5] [0]), .I1(n12_adj_4103), 
            .I2(n32574), .I3(n17926), .O(n17814));
    defparam i6_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1206 (.I0(n32642), .I1(n29905), .I2(\data_in_frame[6] [0]), 
            .I3(GND_net), .O(n33017));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1206.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1207 (.I0(n17466), .I1(n17742), .I2(\data_in_frame[5] [5]), 
            .I3(GND_net), .O(n17745));
    defparam i2_3_lut_adj_1207.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1208 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n33024));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1208.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(n32845), .I3(GND_net), .O(Kp_23__N_930));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13947_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n18736));
    defparam i13947_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13948_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n18737));
    defparam i13948_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n17324));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_LUT4 i13949_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n18738));
    defparam i13949_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_22_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n27716), .O(n2_adj_4105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13950_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n18739));
    defparam i13950_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1210 (.I0(\data_in_frame[4] [3]), .I1(n17731), 
            .I2(\data_in_frame[2] [0]), .I3(n17237), .O(Kp_23__N_933));   // verilog/coms.v(73[16:42])
    defparam i3_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_CARRY add_43_22 (.CI(n27716), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n27717));
    SB_LUT4 i13951_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n18740));
    defparam i13951_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13952_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n18741));
    defparam i13952_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n18740));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13953_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n18742));
    defparam i13953_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13954_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32398), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n18743));
    defparam i13954_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1211 (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_930), 
            .I2(n17396), .I3(\data_in_frame[15] [0]), .O(n33002));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n27753), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_adj_1212 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n17731));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1212.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_21_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n27715), .O(n2_adj_4106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 equal_1541_i5_3_lut_4_lut (.I0(\data_in_frame[6] [3]), .I1(Kp_23__N_930), 
            .I2(n32487), .I3(\data_in_frame[8] [4]), .O(n5_adj_4029));   // verilog/coms.v(74[16:43])
    defparam equal_1541_i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1213 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n17177));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1213.LUT_INIT = 16'h9696;
    SB_CARRY add_43_21 (.CI(n27715), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n27716));
    SB_LUT4 add_43_20_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n27714), .O(n2_adj_4107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n27714), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n27715));
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_in_frame[4] [4]), .I1(n17731), 
            .I2(GND_net), .I3(GND_net), .O(n32866));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_CARRY add_3971_6 (.CI(n27753), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n27754));
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n27752), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_43_19_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n27713), .O(n2_adj_4108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_4109), .S(n8_adj_4016));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n7_adj_4110), .S(n8_adj_4015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n7_adj_4111), .S(n8_adj_4014));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n31964), .S(n31858));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n31962), .S(n31892));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n31960), .S(n31860));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n31958), .S(n31862));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n31956), .S(n31864));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n7_adj_4112), .S(n8_adj_4013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n7_adj_4113), .S(n8_adj_4012));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n31954), .S(n31866));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n31952), .S(n31868));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n31950), .S(n31870));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n31948), .S(n31872));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n31946), .S(n31820));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n31944), .S(n31838));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n31942), .S(n31836));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n31940), .S(n31874));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n31938), .S(n31876));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n31936), .S(n31878));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n31934), .S(n31880));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n31932), .S(n31882));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n31930), .S(n31884));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n31928), .S(n31886));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n31926), .S(n31834));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n31924), .S(n31832));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n31922), .S(n31888));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n31920), .S(n31890));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n31816), .S(n31898));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_5 (.CI(n27752), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n27753));
    SB_LUT4 i1_4_lut_4_lut (.I0(n63), .I1(n771), .I2(n32373), .I3(\FRAME_MATCHER.i_31__N_2457 ), 
            .O(n5_adj_4064));   // verilog/coms.v(157[6] 159[9])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'ha2a0;
    SB_CARRY add_43_19 (.CI(n27713), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n27714));
    SB_LUT4 select_441_Select_1_i1_3_lut_4_lut (.I0(n63), .I1(n771), .I2(\FRAME_MATCHER.i_31__N_2457 ), 
            .I3(n123), .O(n1));   // verilog/coms.v(157[6] 159[9])
    defparam select_441_Select_1_i1_3_lut_4_lut.LUT_INIT = 16'hf0d0;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n27751), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n18277), .D(n33621));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_3971_4 (.CI(n27751), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n27752));
    SB_LUT4 i3_4_lut_adj_1215 (.I0(\data_in_frame[8] [5]), .I1(Kp_23__N_930), 
            .I2(Kp_23__N_933), .I3(n17324), .O(n18035));
    defparam i3_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1216 (.I0(n18102), .I1(n33024), .I2(n32877), 
            .I3(n32587), .O(n10_adj_4061));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1217 (.I0(\data_in_frame[8] [6]), .I1(n8_adj_4068), 
            .I2(Kp_23__N_1032), .I3(n17316), .O(n33008));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1217.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1218 (.I0(\data_in_frame[8] [6]), .I1(n8_adj_4068), 
            .I2(\data_in_frame[9] [0]), .I3(\data_in_frame[11] [2]), .O(n32650));   // verilog/coms.v(77[16:43])
    defparam i2_3_lut_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_4_lut (.I0(n17418), .I1(n32623), .I2(n17427), .I3(\data_in_frame[3] [7]), 
            .O(n16_adj_4043));   // verilog/coms.v(85[17:28])
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n18277), .D(n33862));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n18277), .D(n34449));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n18277), .D(n32826));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n18277), .D(n34574));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n18277), .D(n30869));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n18277), .D(n33844));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n18277), .D(n33843));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n18277), .D(n34825));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n18277), .D(n32721));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n18277), .D(n33395));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n18277), .D(n34686));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n18277), .D(n32741));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n18277), .D(n34435));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n18277), .D(n33462));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n18277), .D(n34432));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4115), .S(n3_adj_4116));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1219 (.I0(n17418), .I1(n32623), .I2(n17427), 
            .I3(\data_in_frame[10] [0]), .O(n30001));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_18_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n27712), .O(n2_adj_4117)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1220 (.I0(n32574), .I1(n17785), .I2(n17751), 
            .I3(n32866), .O(n10_adj_4118));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1221 (.I0(n17177), .I1(n10_adj_4118), .I2(\data_in_frame[7] [0]), 
            .I3(GND_net), .O(n17364));   // verilog/coms.v(75[16:43])
    defparam i5_3_lut_adj_1221.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32491));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1223 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n17751));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1223.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(n17751), .I1(n32638), .I2(GND_net), 
            .I3(GND_net), .O(n18102));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n17785));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1226 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n17768));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1226.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1227 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[5] [4]), 
            .I2(n15437), .I3(\data_in_frame[3] [2]), .O(n17222));
    defparam i3_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1228 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(GND_net), .O(n32521));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1229 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17761));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1229.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1230 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n32452));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1230.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1231 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32525));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1231.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1232 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32518));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1232.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1233 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n32587));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1233.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1234 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n32534));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1234.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1235 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[2] [0]), 
            .I2(n32525), .I3(n32452), .O(n32848));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[11] [4]), .I1(Kp_23__N_1167), 
            .I2(n10_adj_4074), .I3(Kp_23__N_1373), .O(n34494));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_3_lut (.I0(n32763), .I1(n33069), .I2(\data_in_frame[19] [0]), 
            .I3(GND_net), .O(n10_adj_4018));
    defparam i4_4_lut_3_lut.LUT_INIT = 16'h6969;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4119), .S(n3_adj_4120));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4121), .S(n3_adj_4122));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4123), .S(n3_adj_4124));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4125), .S(n3_adj_4126));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4127), .S(n3_adj_4128));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4129), .S(n3_adj_4130));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4131), .S(n3_adj_4132));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4133), .S(n3_adj_4134));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28682_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35078));
    defparam i28682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28683_4_lut (.I0(n35078), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n35079));
    defparam i28683_4_lut.LUT_INIT = 16'ha0a3;
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4135), .S(n3_adj_4136));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4091), .S(n3_adj_4137));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4105), .S(n3_adj_4138));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4106), .S(n3_adj_4139));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4107), .S(n3_adj_4140));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4108), .S(n3_adj_4141));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4117), .S(n3_adj_4142));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4143), .S(n3_adj_4144));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4145), .S(n3_adj_4146));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4147), .S(n3_adj_4148));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4149), .S(n3_adj_4150));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28681_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35077));
    defparam i28681_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4151), .S(n3_adj_4152));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4153), .S(n3_adj_4154));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4155), .S(n3_adj_4156));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4157), .S(n3_adj_4158));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n27750), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_43_18 (.CI(n27712), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n27713));
    SB_CARRY add_3971_3 (.CI(n27750), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n27751));
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4159), .S(n3_adj_4160));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4161), .S(n3_adj_4162));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_4163), .S(n3_adj_4164));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_4165), .S(n3_adj_4166));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_4167), .S(n3_adj_4168));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_4169), .S(n3_adj_4170));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_4171), .S(n3_adj_4172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n18739));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2009866_i1_3_lut (.I0(n37469), .I1(n37613), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4173));
    defparam i2009866_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29571_2_lut (.I0(n37589), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35901));
    defparam i29571_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4174));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4175));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29838_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35875));
    defparam i29838_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29856_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35874));
    defparam i29856_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut_4_lut (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[14] [2]), 
            .I2(n34613), .I3(\data_in_frame[18] [6]), .O(n33069));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4176));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_2_lut_3_lut (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[14] [2]), 
            .I2(n30543), .I3(GND_net), .O(n36));
    defparam i9_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4177));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29834_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35903));
    defparam i29834_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29836_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35902));
    defparam i29836_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_43_17_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n27711), .O(n2_adj_4143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4178));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3350), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3350), 
            .CO(n27750));
    SB_CARRY add_43_17 (.CI(n27711), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n27712));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4179));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_16_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n27710), .O(n2_adj_4145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i29841_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35869));
    defparam i29841_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29819_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35868));
    defparam i29819_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_16 (.CI(n27710), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n27711));
    SB_LUT4 add_43_15_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n27709), .O(n2_adj_4147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_4_lut_adj_1236 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(n32553), .I3(n32645), .O(n29907));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1236.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1237 (.I0(\data_out_frame[24] [5]), .I1(n15386), 
            .I2(n2332), .I3(\data_out_frame[24] [4]), .O(n32721));
    defparam i1_2_lut_3_lut_4_lut_adj_1237.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4180));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4181));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_adj_1238 (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4182));
    defparam i2_2_lut_adj_1238.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1239 (.I0(\FRAME_MATCHER.state [13]), .I1(\FRAME_MATCHER.state [9]), 
            .I2(\FRAME_MATCHER.state [11]), .I3(\FRAME_MATCHER.state [12]), 
            .O(n14_adj_4183));
    defparam i6_4_lut_adj_1239.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1240 (.I0(\FRAME_MATCHER.state [10]), .I1(n14_adj_4183), 
            .I2(n10_adj_4182), .I3(\FRAME_MATCHER.state [8]), .O(n24578));
    defparam i7_4_lut_adj_1240.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1241 (.I0(\FRAME_MATCHER.state [6]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n24390));
    defparam i3_4_lut_adj_1241.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1242 (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [22]), 
            .I2(\FRAME_MATCHER.state [21]), .I3(\FRAME_MATCHER.state [25]), 
            .O(n20_adj_4184));
    defparam i8_4_lut_adj_1242.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1243 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [23]), 
            .I2(\FRAME_MATCHER.state [31]), .I3(\FRAME_MATCHER.state [30]), 
            .O(n19_adj_4185));
    defparam i7_4_lut_adj_1243.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1244 (.I0(\FRAME_MATCHER.state [18]), .I1(\FRAME_MATCHER.state [20]), 
            .I2(\FRAME_MATCHER.state [17]), .I3(\FRAME_MATCHER.state [24]), 
            .O(n38_adj_4186));
    defparam i3_4_lut_adj_1244.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1245 (.I0(\FRAME_MATCHER.state [19]), .I1(\FRAME_MATCHER.state [28]), 
            .I2(\FRAME_MATCHER.state [27]), .I3(\FRAME_MATCHER.state [26]), 
            .O(n21_adj_4187));
    defparam i9_4_lut_adj_1245.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1246 (.I0(n21_adj_4187), .I1(n38_adj_4186), .I2(n19_adj_4185), 
            .I3(n20_adj_4184), .O(n24690));
    defparam i1_4_lut_adj_1246.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_15 (.CI(n27709), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n27710));
    SB_LUT4 i1_3_lut_adj_1247 (.I0(n24690), .I1(n24390), .I2(n24578), 
            .I3(GND_net), .O(n24776));
    defparam i1_3_lut_adj_1247.LUT_INIT = 16'hfefe;
    SB_LUT4 i30428_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17001));   // verilog/coms.v(145[4] 299[11])
    defparam i30428_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_3_lut_adj_1248 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [4]), .I3(GND_net), .O(n31920));
    defparam i1_2_lut_3_lut_adj_1248.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1249 (.I0(n24578), .I1(n24390), .I2(n17001), 
            .I3(n24690), .O(n10_adj_4189));
    defparam i4_4_lut_adj_1249.LUT_INIT = 16'hffef;
    SB_LUT4 i30889_3_lut (.I0(n17017), .I1(n10_adj_4189), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(GND_net), .O(n34324));
    defparam i30889_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i19609_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n66), .I2(n17068), 
            .I3(n17089), .O(n2236));
    defparam i19609_4_lut.LUT_INIT = 16'h2aaa;
    SB_LUT4 i1_2_lut_3_lut_adj_1250 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [5]), .I3(GND_net), .O(n31922));
    defparam i1_2_lut_3_lut_adj_1250.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(n24219), .I1(n10_adj_4190), .I2(GND_net), 
            .I3(GND_net), .O(n32406));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_adj_1252 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [6]), .I3(GND_net), .O(n31924));
    defparam i1_2_lut_3_lut_adj_1252.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1253 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [7]), .I3(GND_net), .O(n31926));
    defparam i1_2_lut_3_lut_adj_1253.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n18738));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_14_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n27708), .O(n2_adj_4149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_14 (.CI(n27708), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n27709));
    SB_LUT4 add_43_13_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n27707), .O(n2_adj_4151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n18737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n18736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n18735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n18734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n18733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n18732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n18731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n18730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n18729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n18728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n18727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n18726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n18725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n18724));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n18723));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n18722));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n18721));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n18720));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n18719));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n18718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n18717));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n18716));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n18715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n18714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n18713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n18712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n18711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n18710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n18709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n18708));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n18707));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30886_4_lut (.I0(n17017), .I1(n5202), .I2(n5_adj_4191), .I3(n6_adj_4192), 
            .O(n32337));
    defparam i30886_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_in_frame[5] [6]), .I1(n17466), 
            .I2(GND_net), .I3(GND_net), .O(n32808));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1255 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [8]), .I3(GND_net), .O(n31928));
    defparam i1_2_lut_3_lut_adj_1255.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n18706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n18705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n18704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n18703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n18702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n18701));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n18700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n18699));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n18698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n18697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n18693));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[24] [5]), .I1(n15386), .I2(\data_out_frame[24] [6]), 
            .I3(GND_net), .O(n7_adj_3968));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY add_43_13 (.CI(n27707), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n27708));
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[3] [1]), .I1(\data_in_frame[5] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n32605));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [9]), .I3(GND_net), .O(n31930));
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'he0e0;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n18692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n18691));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n18690));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n18689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n18688));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n18687));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i11_4_lut_adj_1258 (.I0(n32869), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[2] [2]), .I3(n32605), .O(n30_adj_4193));   // verilog/coms.v(78[16:27])
    defparam i11_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1259 (.I0(\data_in_frame[3] [7]), .I1(n30_adj_4193), 
            .I2(\data_in_frame[5] [1]), .I3(n32553), .O(n34_adj_4194));   // verilog/coms.v(78[16:27])
    defparam i15_4_lut_adj_1259.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1260 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [10]), .I3(GND_net), .O(n31932));
    defparam i1_2_lut_3_lut_adj_1260.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_12_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n27706), .O(n2_adj_4153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13_4_lut_adj_1261 (.I0(n32848), .I1(n32534), .I2(n32587), 
            .I3(n32518), .O(n32_adj_4195));   // verilog/coms.v(78[16:27])
    defparam i13_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1262 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [11]), .I3(GND_net), .O(n31934));
    defparam i1_2_lut_3_lut_adj_1262.LUT_INIT = 16'he0e0;
    SB_LUT4 i29793_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35909));
    defparam i29793_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29791_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35908));
    defparam i29791_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_12 (.CI(n27706), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n27707));
    SB_LUT4 add_43_11_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n27705), .O(n2_adj_4155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1263 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [12]), .I3(GND_net), .O(n31936));
    defparam i1_2_lut_3_lut_adj_1263.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_adj_1264 (.I0(\FRAME_MATCHER.state [2]), .I1(n18216), 
            .I2(n77), .I3(GND_net), .O(n20456));   // verilog/coms.v(112[11:16])
    defparam i1_3_lut_adj_1264.LUT_INIT = 16'hc4c4;
    SB_LUT4 i14_4_lut_adj_1265 (.I0(\data_in_frame[0] [2]), .I1(n17761), 
            .I2(\data_in_frame[5] [7]), .I3(\data_in_frame[3] [0]), .O(n33));   // verilog/coms.v(78[16:27])
    defparam i14_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1266 (.I0(n17745), .I1(n17751), .I2(n32638), 
            .I3(n33017), .O(n30028));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_CARRY add_43_11 (.CI(n27705), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n27706));
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1267 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(n32529), .I3(\data_out_frame[17] [5]), .O(n32664));
    defparam i1_2_lut_3_lut_4_lut_adj_1267.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1268 (.I0(n32521), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[2] [7]), .I3(n17222), .O(n31_adj_4196));   // verilog/coms.v(78[16:27])
    defparam i12_4_lut_adj_1268.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1269 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[4] [5]), .O(n32638));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1270 (.I0(n31_adj_4196), .I1(n33), .I2(n32_adj_4195), 
            .I3(n34_adj_4194), .O(n29905));   // verilog/coms.v(78[16:27])
    defparam i18_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i28594_2_lut_3_lut_4_lut (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(n17751), .O(n34988));   // verilog/coms.v(166[9:87])
    defparam i28594_2_lut_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1271 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[4] [6]), .O(n32574));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1272 (.I0(\data_out_frame[20] [4]), .I1(n33521), 
            .I2(\data_out_frame[20] [3]), .I3(n34478), .O(n30832));
    defparam i1_2_lut_3_lut_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_10_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n27704), .O(n2_adj_4157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_10 (.CI(n27704), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n27705));
    SB_LUT4 i30883_2_lut (.I0(n24682), .I1(n10932), .I2(GND_net), .I3(GND_net), 
            .O(tx_transmit_N_3350));
    defparam i30883_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1273 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n24776), .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n17089));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1273.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1274 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[5] [4]), .I3(\data_out_frame[7] [5]), .O(n33027));
    defparam i1_2_lut_3_lut_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1275 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[5] [7]), .I3(\data_out_frame[5] [6]), .O(n33014));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i28603_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17001), .I3(n24776), .O(n34998));
    defparam i28603_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i2_3_lut_adj_1276 (.I0(n34998), .I1(\FRAME_MATCHER.i_31__N_2460 ), 
            .I2(n2236), .I3(GND_net), .O(n33978));
    defparam i2_3_lut_adj_1276.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\FRAME_MATCHER.i [4]), .I1(n17014), .I2(GND_net), 
            .I3(GND_net), .O(n16911));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'heeee;
    SB_LUT4 i19017_4_lut (.I0(n5_adj_4197), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(\FRAME_MATCHER.i [3]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i19017_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i19022_4_lut (.I0(n8_adj_4104), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n16911), .I3(\FRAME_MATCHER.i [3]), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i19022_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i1_2_lut_adj_1278 (.I0(\FRAME_MATCHER.state[0] ), .I1(n17089), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2457 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1278.LUT_INIT = 16'h2222;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n18686));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1279 (.I0(\FRAME_MATCHER.state[0] ), .I1(n17068), 
            .I2(GND_net), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2461 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1279.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1280 (.I0(\data_in[0] [3]), .I1(\data_in[1] [0]), 
            .I2(\data_in[2] [2]), .I3(GND_net), .O(n34138));
    defparam i2_3_lut_adj_1280.LUT_INIT = 16'h8080;
    SB_LUT4 i5_4_lut_adj_1281 (.I0(\data_in[0] [6]), .I1(n17065), .I2(\data_in[2] [4]), 
            .I3(n34138), .O(n12_adj_4198));
    defparam i5_4_lut_adj_1281.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1282 (.I0(\data_in[3] [0]), .I1(n12_adj_4198), 
            .I2(\data_in[1] [4]), .I3(\data_in[1] [5]), .O(n16914));
    defparam i6_4_lut_adj_1282.LUT_INIT = 16'hfdff;
    SB_LUT4 i4_4_lut_adj_1283 (.I0(\data_in[0] [4]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [7]), .I3(\data_in[3] [4]), .O(n10_adj_4199));
    defparam i4_4_lut_adj_1283.LUT_INIT = 16'hdfff;
    SB_LUT4 i5_3_lut_adj_1284 (.I0(\data_in[1] [1]), .I1(n10_adj_4199), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n17065));
    defparam i5_3_lut_adj_1284.LUT_INIT = 16'hefef;
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n18685));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_1285 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4200));
    defparam i6_4_lut_adj_1285.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1286 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4201));
    defparam i7_4_lut_adj_1286.LUT_INIT = 16'hfffd;
    SB_LUT4 add_43_9_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n27703), .O(n2_adj_4159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n18216), .D(n8825[0]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35079), .I3(n35077), .O(n7_adj_4202));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i9_4_lut_adj_1287 (.I0(n17_adj_4201), .I1(\data_in[1] [6]), 
            .I2(n16_adj_4200), .I3(\data_in[3] [7]), .O(n17011));
    defparam i9_4_lut_adj_1287.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_2_lut_adj_1288 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4203));
    defparam i2_2_lut_adj_1288.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1289 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4204));
    defparam i6_4_lut_adj_1289.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1290 (.I0(\data_in[3] [6]), .I1(n14_adj_4204), 
            .I2(n10_adj_4203), .I3(\data_in[2] [1]), .O(n17008));
    defparam i7_4_lut_adj_1290.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1291 (.I0(\data_in[2] [4]), .I1(\data_in[2] [2]), 
            .I2(n17008), .I3(\data_in[1] [0]), .O(n18_adj_4205));
    defparam i7_4_lut_adj_1291.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1292 (.I0(\data_in[1] [4]), .I1(n18_adj_4205), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n20_adj_4206));
    defparam i9_4_lut_adj_1292.LUT_INIT = 16'hfffd;
    SB_LUT4 i10_4_lut_adj_1293 (.I0(n15_adj_4207), .I1(n20_adj_4206), .I2(n17011), 
            .I3(\data_in[0] [6]), .O(n63_c));
    defparam i10_4_lut_adj_1293.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1294 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n16914), .O(n16_adj_4208));
    defparam i6_4_lut_adj_1294.LUT_INIT = 16'hffef;
    SB_LUT4 i7_4_lut_adj_1295 (.I0(n17011), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [1]), .O(n17_adj_4209));
    defparam i7_4_lut_adj_1295.LUT_INIT = 16'hbfff;
    SB_LUT4 i9_4_lut_adj_1296 (.I0(n17_adj_4209), .I1(\data_in[3] [5]), 
            .I2(n16_adj_4208), .I3(\data_in[3] [3]), .O(n63_adj_4057));
    defparam i9_4_lut_adj_1296.LUT_INIT = 16'hfbff;
    SB_LUT4 i5_3_lut_adj_1297 (.I0(\data_in[0] [5]), .I1(\data_in[2] [6]), 
            .I2(\data_in[3] [7]), .I3(GND_net), .O(n14_adj_4210));
    defparam i5_3_lut_adj_1297.LUT_INIT = 16'hfdfd;
    SB_LUT4 i3_4_lut_adj_1298 (.I0(\data_in[1] [3]), .I1(\data_in[3] [2]), 
            .I2(\data_in[1] [2]), .I3(\data_in[2] [5]), .O(n34684));
    defparam i3_4_lut_adj_1298.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_1299 (.I0(\data_in[1] [6]), .I1(n17008), .I2(\data_in[0] [1]), 
            .I3(n16914), .O(n15_adj_4211));
    defparam i6_4_lut_adj_1299.LUT_INIT = 16'hffef;
    SB_LUT4 i8_4_lut_adj_1300 (.I0(n15_adj_4211), .I1(n34684), .I2(n14_adj_4210), 
            .I3(\data_in[2] [0]), .O(n63));
    defparam i8_4_lut_adj_1300.LUT_INIT = 16'hfbff;
    SB_LUT4 i18_4_lut_adj_1301 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_4212));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut_adj_1301.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1302 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [13]), .I3(GND_net), .O(n31938));
    defparam i1_2_lut_3_lut_adj_1302.LUT_INIT = 16'he0e0;
    SB_LUT4 i16_4_lut_adj_1303 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_4213));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut_adj_1303.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1304 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_4214));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut_adj_1304.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1305 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_4215));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut_adj_1305.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1306 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_4216));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut_adj_1306.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4217));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut_adj_1307 (.I0(n41_adj_4215), .I1(n43_adj_4214), .I2(n42_adj_4213), 
            .I3(n44_adj_4212), .O(n50_adj_4218));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut_adj_1307.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35112), .I3(n35110), .O(n7_adj_4219));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i19_4_lut_adj_1308 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45_adj_4220));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut_adj_1308.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1309 (.I0(n45_adj_4220), .I1(n50_adj_4218), .I2(n39_adj_4217), 
            .I3(n40_adj_4216), .O(n17014));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut_adj_1309.LUT_INIT = 16'hfffe;
    SB_LUT4 i19023_4_lut (.I0(n8_adj_4221), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n17014), .I3(\FRAME_MATCHER.i [4]), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i19023_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i19025_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n14278), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2497 [0]));
    defparam i19025_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_1310 (.I0(\FRAME_MATCHER.state [2]), .I1(n77), 
            .I2(\FRAME_MATCHER.state_31__N_2497 [0]), .I3(n4452), .O(n33875));   // verilog/coms.v(112[11:16])
    defparam i3_4_lut_adj_1310.LUT_INIT = 16'hffef;
    SB_LUT4 i1_4_lut_adj_1311 (.I0(\FRAME_MATCHER.i_31__N_2461 ), .I1(\FRAME_MATCHER.i_31__N_2457 ), 
            .I2(n3303), .I3(n771), .O(n4_adj_4222));
    defparam i1_4_lut_adj_1311.LUT_INIT = 16'h0ace;
    SB_LUT4 i2_4_lut_adj_1312 (.I0(\FRAME_MATCHER.state_31__N_2497 [0]), .I1(n34405), 
            .I2(n4_adj_4222), .I3(n33875), .O(n33985));
    defparam i2_4_lut_adj_1312.LUT_INIT = 16'hb3ff;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35103), .I3(n35101), .O(n7_adj_4223));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35097), .I3(n35095), .O(n7_adj_4224));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i18883_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3453[0]), .I2(GND_net), 
            .I3(GND_net), .O(n23655));
    defparam i18883_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19458_2_lut (.I0(byte_transmit_counter[0]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n24235));
    defparam i19458_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1313 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n24235), .I3(byte_transmit_counter[2]), .O(n24682));
    defparam i2_4_lut_adj_1313.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut_adj_1314 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n74));
    defparam i1_2_lut_adj_1314.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1315 (.I0(byte_transmit_counter[5]), .I1(byte_transmit_counter[7]), 
            .I2(byte_transmit_counter[6]), .I3(GND_net), .O(n10932));   // verilog/coms.v(214[11:56])
    defparam i2_3_lut_adj_1315.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4225));
    defparam i15_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_3_lut_adj_1316 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [14]), .I3(GND_net), .O(n31940));
    defparam i1_2_lut_3_lut_adj_1316.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_4_lut_adj_1317 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [3]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n34921));
    defparam i2_4_lut_adj_1317.LUT_INIT = 16'h0504;
    SB_LUT4 i30432_4_lut (.I0(n62_adj_4226), .I1(n24776), .I2(n47_adj_4225), 
            .I3(n34921), .O(n3482));
    defparam i30432_4_lut.LUT_INIT = 16'hccce;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35073), .I3(n35071), .O(n7_adj_4227));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i3_3_lut_adj_1318 (.I0(n10932), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n74), .I3(GND_net), .O(n8_adj_4228));
    defparam i3_3_lut_adj_1318.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_2_lut_adj_1319 (.I0(n24682), .I1(n23655), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4229));
    defparam i2_2_lut_adj_1319.LUT_INIT = 16'heeee;
    SB_LUT4 mux_899_i1_4_lut (.I0(n7_adj_4229), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n5202), .I3(n8_adj_4228), .O(n3519[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_899_i1_4_lut.LUT_INIT = 16'h0c5c;
    SB_LUT4 i30412_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n10_adj_4230), .I3(n24578), .O(n18241));
    defparam i30412_3_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1320 (.I0(\data_in_frame[10] [7]), .I1(Kp_23__N_1032), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[8] [6]), .O(n32611));
    defparam i1_2_lut_3_lut_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35085), .I3(n35083), .O(n7_adj_4231));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_CARRY add_43_9 (.CI(n27703), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n27704));
    SB_LUT4 add_43_8_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n27702), .O(n2_adj_4161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_8 (.CI(n27702), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n27703));
    SB_LUT4 add_43_7_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n27701), .O(n2_adj_4163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1321 (.I0(n17370), .I1(n17358), .I2(\data_in_frame[8] [2]), 
            .I3(n15471), .O(n32667));
    defparam i1_2_lut_3_lut_4_lut_adj_1321.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1322 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[6] [1]), .I3(GND_net), .O(n6_adj_4232));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1322.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1323 (.I0(n17370), .I1(\data_in_frame[8] [3]), 
            .I2(n32487), .I3(n18035), .O(n17246));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1323.LUT_INIT = 16'h6996;
    SB_CARRY add_43_7 (.CI(n27701), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n27702));
    SB_LUT4 add_43_6_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n27700), .O(n2_adj_4165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_6 (.CI(n27700), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n27701));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35091), .I3(n35089), .O(n7_adj_4233));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_43_5_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n27699), .O(n2_adj_4167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n5300));
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'h0202;
    SB_LUT4 i19995_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n24776), .O(n5202));
    defparam i19995_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1325 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n62_adj_4226));
    defparam i1_2_lut_3_lut_adj_1325.LUT_INIT = 16'hfefe;
    SB_CARRY add_43_5 (.CI(n27699), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n27700));
    SB_LUT4 i1_2_lut_3_lut_adj_1326 (.I0(\FRAME_MATCHER.state[0] ), .I1(n14278), 
            .I2(n32404), .I3(GND_net), .O(n31814));
    defparam i1_2_lut_3_lut_adj_1326.LUT_INIT = 16'hb0b0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n35070), .I3(n35068), .O(n7_adj_4234));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i14078_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n18867));
    defparam i14078_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_in[1] [1]), .I1(n10_adj_4199), .I2(\data_in[2] [7]), 
            .I3(\data_in[3] [0]), .O(n15_adj_4207));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_1327 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n32880));
    defparam i1_2_lut_3_lut_adj_1327.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1328 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [15]), .I3(GND_net), .O(n31942));
    defparam i1_2_lut_3_lut_adj_1328.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_4_lut_adj_1329 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n17014), .I3(\FRAME_MATCHER.i [1]), .O(n5_adj_4197));
    defparam i1_3_lut_4_lut_adj_1329.LUT_INIT = 16'hfefc;
    SB_LUT4 add_43_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n27698), .O(n2_adj_4169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_4 (.CI(n27698), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n27699));
    SB_LUT4 i1_2_lut_3_lut_adj_1330 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [16]), .I3(GND_net), .O(n31944));
    defparam i1_2_lut_3_lut_adj_1330.LUT_INIT = 16'he0e0;
    SB_LUT4 i14079_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n18868));
    defparam i14079_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_3_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n27697), .O(n2_adj_4171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_4_lut_adj_1331 (.I0(n33978), .I1(tx_transmit_N_3350), 
            .I2(n23655), .I3(\FRAME_MATCHER.i_31__N_2460 ), .O(n32404));
    defparam i1_2_lut_4_lut_adj_1331.LUT_INIT = 16'hfd55;
    SB_LUT4 i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n17001), 
            .I2(n24776), .I3(\FRAME_MATCHER.state [3]), .O(n34405));   // verilog/coms.v(201[5:24])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_3_lut_adj_1332 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [17]), .I3(GND_net), .O(n31946));
    defparam i1_2_lut_3_lut_adj_1332.LUT_INIT = 16'he0e0;
    SB_CARRY add_43_3 (.CI(n27697), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n27698));
    SB_LUT4 i14080_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n18869));
    defparam i14080_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n37610));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37610_bdd_4_lut (.I0(n37610), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n37613));
    defparam n37610_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n37349), .I2(n35870), .I3(byte_transmit_counter[4]), .O(n37604));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37604_bdd_4_lut (.I0(n37604), .I1(n14_adj_4235), .I2(n7_adj_4231), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n37604_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31164 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n37598));
    defparam byte_transmit_counter_0__bdd_4_lut_31164.LUT_INIT = 16'he4aa;
    SB_LUT4 n37598_bdd_4_lut (.I0(n37598), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n37601));
    defparam n37598_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31159 (.I0(byte_transmit_counter[3]), 
            .I1(n37361), .I2(n35864), .I3(byte_transmit_counter[4]), .O(n37592));
    defparam byte_transmit_counter_3__bdd_4_lut_31159.LUT_INIT = 16'he4aa;
    SB_LUT4 n37592_bdd_4_lut (.I0(n37592), .I1(n14_adj_4236), .I2(n7_adj_4233), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n37592_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31154 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n37586));
    defparam byte_transmit_counter_0__bdd_4_lut_31154.LUT_INIT = 16'he4aa;
    SB_LUT4 n37586_bdd_4_lut (.I0(n37586), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n37589));
    defparam n37586_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_adj_1333 (.I0(n34405), .I1(\FRAME_MATCHER.i_31__N_2460 ), 
            .I2(tx_active), .I3(r_SM_Main_2__N_3453[0]), .O(n18216));   // verilog/coms.v(201[5:24])
    defparam i1_3_lut_4_lut_adj_1333.LUT_INIT = 16'h555d;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31144 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n37580));
    defparam byte_transmit_counter_0__bdd_4_lut_31144.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1334 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [18]), .I3(GND_net), .O(n31948));
    defparam i1_2_lut_3_lut_adj_1334.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1335 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[2] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [4]), .O(n32869));
    defparam i1_2_lut_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i14081_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n18870));
    defparam i14081_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1336 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [6]), 
            .I2(n17466), .I3(GND_net), .O(n32553));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1336.LUT_INIT = 16'h9696;
    SB_LUT4 i30896_2_lut_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n18460));
    defparam i30896_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i14082_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n18871));
    defparam i14082_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n37580_bdd_4_lut (.I0(n37580), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n37583));
    defparam n37580_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n1_adj_4237), .I3(GND_net), .O(n5_adj_4191));
    defparam i1_4_lut_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31139 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n37574));
    defparam byte_transmit_counter_0__bdd_4_lut_31139.LUT_INIT = 16'he4aa;
    SB_LUT4 n37574_bdd_4_lut (.I0(n37574), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n37577));
    defparam n37574_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31134 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n37568));
    defparam byte_transmit_counter_0__bdd_4_lut_31134.LUT_INIT = 16'he4aa;
    SB_LUT4 n37568_bdd_4_lut (.I0(n37568), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n37571));
    defparam n37568_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1337 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [19]), .I3(GND_net), .O(n31950));
    defparam i1_2_lut_3_lut_adj_1337.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31129 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n37562));
    defparam byte_transmit_counter_0__bdd_4_lut_31129.LUT_INIT = 16'he4aa;
    SB_LUT4 n37562_bdd_4_lut (.I0(n37562), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n37565));
    defparam n37562_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [20]), .I3(GND_net), .O(n31952));
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31124 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n37556));
    defparam byte_transmit_counter_0__bdd_4_lut_31124.LUT_INIT = 16'he4aa;
    SB_LUT4 n37556_bdd_4_lut (.I0(n37556), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n37559));
    defparam n37556_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31119 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n37550));
    defparam byte_transmit_counter_0__bdd_4_lut_31119.LUT_INIT = 16'he4aa;
    SB_LUT4 n37550_bdd_4_lut (.I0(n37550), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n37553));
    defparam n37550_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i19444_2_lut_3_lut (.I0(n2236), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n24219));
    defparam i19444_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i14083_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n18872));
    defparam i14083_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14084_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n18873));
    defparam i14084_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19340_2_lut_4_lut (.I0(n14565), .I1(n31_adj_4099), .I2(n31_adj_4238), 
            .I3(\FRAME_MATCHER.state [1]), .O(n1_adj_4237));
    defparam i19340_2_lut_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i13849_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32391), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n18638));
    defparam i13849_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [21]), .I3(GND_net), .O(n31954));
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_2_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_3_lut_4_lut_adj_1340 (.I0(n3482), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n62_adj_4226), .I3(n24776), .O(n17017));
    defparam i1_3_lut_4_lut_adj_1340.LUT_INIT = 16'haaae;
    SB_LUT4 i2_3_lut_4_lut_adj_1341 (.I0(n31_adj_4238), .I1(n14565), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n17092), .O(n34118));
    defparam i2_3_lut_4_lut_adj_1341.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [22]), .I3(GND_net), .O(n7_adj_4113));
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31114 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n37532));
    defparam byte_transmit_counter_0__bdd_4_lut_31114.LUT_INIT = 16'he4aa;
    SB_LUT4 n37532_bdd_4_lut (.I0(n37532), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n37535));
    defparam n37532_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31099 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n37526));
    defparam byte_transmit_counter_0__bdd_4_lut_31099.LUT_INIT = 16'he4aa;
    SB_LUT4 n37526_bdd_4_lut (.I0(n37526), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n37529));
    defparam n37526_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31094 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n37520));
    defparam byte_transmit_counter_0__bdd_4_lut_31094.LUT_INIT = 16'he4aa;
    SB_LUT4 n37520_bdd_4_lut (.I0(n37520), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n37523));
    defparam n37520_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [23]), .I3(GND_net), .O(n7_adj_4112));
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'he0e0;
    SB_LUT4 i1351_2_lut_3_lut (.I0(n31_adj_4238), .I1(n14565), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n5063));
    defparam i1351_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut_3_lut_adj_1344 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [24]), .I3(GND_net), .O(n31956));
    defparam i1_2_lut_3_lut_adj_1344.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1345 (.I0(n32763), .I1(n29854), .I2(n33050), 
            .I3(\data_in_frame[18] [7]), .O(n32709));
    defparam i1_2_lut_3_lut_4_lut_adj_1345.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31089 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n37514));
    defparam byte_transmit_counter_0__bdd_4_lut_31089.LUT_INIT = 16'he4aa;
    SB_LUT4 n37514_bdd_4_lut (.I0(n37514), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n37517));
    defparam n37514_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1346 (.I0(\data_in_frame[11] [4]), .I1(n17364), 
            .I2(n10_adj_4061), .I3(\data_in_frame[11] [5]), .O(n6_adj_4040));
    defparam i1_2_lut_3_lut_4_lut_adj_1346.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31084 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n37508));
    defparam byte_transmit_counter_0__bdd_4_lut_31084.LUT_INIT = 16'he4aa;
    SB_LUT4 n37508_bdd_4_lut (.I0(n37508), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n37511));
    defparam n37508_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31079 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n37502));
    defparam byte_transmit_counter_0__bdd_4_lut_31079.LUT_INIT = 16'he4aa;
    SB_LUT4 n37502_bdd_4_lut (.I0(n37502), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n37505));
    defparam n37502_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut_adj_1347 (.I0(n17370), .I1(n17358), .I2(\data_in_frame[8] [2]), 
            .I3(GND_net), .O(n17391));   // verilog/coms.v(236[9:81])
    defparam i2_2_lut_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31074 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n37496));
    defparam byte_transmit_counter_0__bdd_4_lut_31074.LUT_INIT = 16'he4aa;
    SB_LUT4 n37496_bdd_4_lut (.I0(n37496), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n37499));
    defparam n37496_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31069 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n37490));
    defparam byte_transmit_counter_0__bdd_4_lut_31069.LUT_INIT = 16'he4aa;
    SB_LUT4 i14062_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n18851));
    defparam i14062_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(n17198), .I1(\data_in_frame[13] [5]), 
            .I2(n32933), .I3(n33060), .O(n8_adj_4072));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [25]), .I3(GND_net), .O(n31958));
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1349 (.I0(n17198), .I1(\data_in_frame[13] [5]), 
            .I2(n32933), .I3(\data_in_frame[15] [7]), .O(n32731));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1349.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1350 (.I0(\data_out_frame[24] [4]), .I1(n2332), 
            .I2(\data_out_frame[24] [3]), .I3(n34610), .O(n33395));
    defparam i2_3_lut_4_lut_adj_1350.LUT_INIT = 16'h9669;
    SB_LUT4 i14063_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n18852));
    defparam i14063_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14064_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n18853));
    defparam i14064_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[4] [2]), .I3(GND_net), .O(n17237));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1352 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[4] [0]), .O(n6_adj_4100));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i14065_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n18854));
    defparam i14065_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14066_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n18855));
    defparam i14066_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14067_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n18856));
    defparam i14067_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n37490_bdd_4_lut (.I0(n37490), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n37493));
    defparam n37490_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14068_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n18857));
    defparam i14068_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1353 (.I0(n17068), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n14565), .I3(n31_adj_4099), .O(n34304));
    defparam i2_3_lut_4_lut_adj_1353.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31149 (.I0(byte_transmit_counter[3]), 
            .I1(n37367), .I2(n35907), .I3(byte_transmit_counter[4]), .O(n37484));
    defparam byte_transmit_counter_3__bdd_4_lut_31149.LUT_INIT = 16'he4aa;
    SB_LUT4 n37484_bdd_4_lut (.I0(n37484), .I1(n14_adj_4240), .I2(n7_adj_4234), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n37484_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1354 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[0] [0]), .I3(n17237), .O(n32845));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31064 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n37466));
    defparam byte_transmit_counter_0__bdd_4_lut_31064.LUT_INIT = 16'he4aa;
    SB_LUT4 n37466_bdd_4_lut (.I0(n37466), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n37469));
    defparam n37466_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1355 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [26]), .I3(GND_net), .O(n31960));
    defparam i1_2_lut_3_lut_adj_1355.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(n17751), .I1(n32638), .I2(n33017), 
            .I3(GND_net), .O(n32645));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1357 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[1] [1]), .O(n17742));   // verilog/coms.v(73[16:34])
    defparam i2_3_lut_4_lut_adj_1357.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1358 (.I0(n17589), .I1(\data_in_frame[0] [7]), 
            .I2(Kp_23__N_825), .I3(n32605), .O(n6_adj_4102));
    defparam i1_2_lut_4_lut_adj_1358.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1359 (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[5] [1]), 
            .I2(n32877), .I3(\data_in_frame[3] [1]), .O(n32863));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31044 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n37454));
    defparam byte_transmit_counter_0__bdd_4_lut_31044.LUT_INIT = 16'he4aa;
    SB_LUT4 n37454_bdd_4_lut (.I0(n37454), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n37457));
    defparam n37454_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31034 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n37448));
    defparam byte_transmit_counter_0__bdd_4_lut_31034.LUT_INIT = 16'he4aa;
    SB_LUT4 n37448_bdd_4_lut (.I0(n37448), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n37451));
    defparam n37448_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(n17370), .I1(\data_in_frame[8] [3]), 
            .I2(n32487), .I3(GND_net), .O(n17820));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31059 (.I0(byte_transmit_counter[3]), 
            .I1(n37439), .I2(n35904), .I3(byte_transmit_counter[4]), .O(n37442));
    defparam byte_transmit_counter_3__bdd_4_lut_31059.LUT_INIT = 16'he4aa;
    SB_LUT4 n37442_bdd_4_lut (.I0(n37442), .I1(n14_adj_4241), .I2(n7_adj_4227), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n37442_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n27697));
    SB_LUT4 i14069_3_lut_4_lut (.I0(n10_adj_4239), .I1(n32384), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n18858));
    defparam i14069_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n35905), .I2(n35906), .I3(byte_transmit_counter[2]), .O(n37436));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37436_bdd_4_lut (.I0(n37436), .I1(n17_adj_4242), .I2(n16_adj_4243), 
            .I3(byte_transmit_counter[2]), .O(n37439));
    defparam n37436_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31029 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n37430));
    defparam byte_transmit_counter_0__bdd_4_lut_31029.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1361 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [4]), 
            .I2(n32728), .I3(n33038), .O(n6));
    defparam i1_2_lut_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1362 (.I0(n32611), .I1(n10_adj_4038), .I2(n15478), 
            .I3(n32475), .O(n6_adj_4078));
    defparam i1_2_lut_4_lut_adj_1362.LUT_INIT = 16'h6996;
    SB_LUT4 n37430_bdd_4_lut (.I0(n37430), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n37433));
    defparam n37430_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_2_lut_3_lut (.I0(n17699), .I1(\data_in_frame[17] [7]), .I2(\data_in_frame[17] [6]), 
            .I3(GND_net), .O(n13_adj_4087));
    defparam i4_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1363 (.I0(n17466), .I1(n17222), .I2(\data_in_frame[7] [6]), 
            .I3(GND_net), .O(n17427));
    defparam i1_2_lut_3_lut_adj_1363.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31024 (.I0(byte_transmit_counter[3]), 
            .I1(n37373), .I2(n35861), .I3(byte_transmit_counter[4]), .O(n37412));
    defparam byte_transmit_counter_3__bdd_4_lut_31024.LUT_INIT = 16'he4aa;
    SB_LUT4 n37412_bdd_4_lut (.I0(n37412), .I1(n14_adj_4244), .I2(n7_adj_4224), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n37412_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_4_lut (.I0(n17246), .I1(n32942), .I2(\data_in_frame[15] [3]), 
            .I3(n17391), .O(n10_adj_4070));   // verilog/coms.v(71[16:27])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [27]), .I3(GND_net), .O(n31962));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_31014 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n37406));
    defparam byte_transmit_counter_0__bdd_4_lut_31014.LUT_INIT = 16'he4aa;
    SB_LUT4 i4_4_lut_adj_1365 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[6] [5]), 
            .I2(n17324), .I3(n6_adj_4232), .O(n32642));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 n37406_bdd_4_lut (.I0(n37406), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n37409));
    defparam n37406_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1366 (.I0(n32642), .I1(n32880), .I2(n29905), 
            .I3(\data_in_frame[1] [3]), .O(n12_adj_4245));
    defparam i5_4_lut_adj_1366.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1367 (.I0(\data_in_frame[8] [1]), .I1(n12_adj_4245), 
            .I2(n18102), .I3(\data_in_frame[3] [6]), .O(n34602));
    defparam i6_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i14046_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n18835));
    defparam i14046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14047_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n18836));
    defparam i14047_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14048_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n18837));
    defparam i14048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14049_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n18838));
    defparam i14049_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14050_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n18839));
    defparam i14050_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_31000 (.I0(byte_transmit_counter[3]), 
            .I1(n37379), .I2(n35912), .I3(byte_transmit_counter[4]), .O(n37400));
    defparam byte_transmit_counter_3__bdd_4_lut_31000.LUT_INIT = 16'he4aa;
    SB_LUT4 n37400_bdd_4_lut (.I0(n37400), .I1(n14_adj_4246), .I2(n7_adj_4223), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n37400_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30990 (.I0(byte_transmit_counter[3]), 
            .I1(n37385), .I2(n35891), .I3(byte_transmit_counter[4]), .O(n37394));
    defparam byte_transmit_counter_3__bdd_4_lut_30990.LUT_INIT = 16'he4aa;
    SB_LUT4 n37394_bdd_4_lut (.I0(n37394), .I1(n14_adj_4247), .I2(n7_adj_4219), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n37394_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14051_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n18840));
    defparam i14051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(Kp_23__N_1032), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[8] [6]), .I3(GND_net), .O(n32960));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30995 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n37388));
    defparam byte_transmit_counter_0__bdd_4_lut_30995.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [28]), .I3(GND_net), .O(n31964));
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'he0e0;
    SB_LUT4 i14052_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n18841));
    defparam i14052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .E(n18470), 
            .D(n17001), .R(n34936));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1370 (.I0(n29907), .I1(n17814), .I2(\data_in_frame[8] [0]), 
            .I3(GND_net), .O(n18_adj_4248));
    defparam i2_3_lut_adj_1370.LUT_INIT = 16'heded;
    SB_LUT4 i14053_3_lut_4_lut (.I0(n8), .I1(n32391), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n18842));
    defparam i14053_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1371 (.I0(\data_in_frame[11] [1]), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[10] [5]), .I3(n33066), .O(n32494));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_LUT4 select_413_Select_1_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4172));
    defparam select_413_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_2_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4170));
    defparam select_413_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_3_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4168));
    defparam select_413_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_4_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4166));
    defparam select_413_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_5_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4164));
    defparam select_413_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_6_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4162));
    defparam select_413_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_7_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4160));
    defparam select_413_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_8_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4158));
    defparam select_413_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i1_2_lut_4_lut_adj_1372 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(n32869), .O(n6_adj_4065));
    defparam i1_2_lut_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1373 (.I0(n17364), .I1(n17391), .I2(n10_adj_4061), 
            .I3(n18035), .O(n26_adj_4249));
    defparam i10_4_lut_adj_1373.LUT_INIT = 16'hfffe;
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n18684));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n37388_bdd_4_lut (.I0(n37388), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n37391));
    defparam n37388_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 select_413_Select_9_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4156));
    defparam select_413_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_10_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4154));
    defparam select_413_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_11_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4152));
    defparam select_413_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_12_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4150));
    defparam select_413_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_13_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4148));
    defparam select_413_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n32337), .D(n18460), 
            .R(n34324));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_413_Select_14_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4146));
    defparam select_413_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 add_43_33_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n27727), .O(n2_adj_4115)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i28607_2_lut (.I0(n17427), .I1(n17418), .I2(GND_net), .I3(GND_net), 
            .O(n35002));
    defparam i28607_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1374 (.I0(Kp_23__N_1032), .I1(n30028), .I2(\data_in_frame[8] [6]), 
            .I3(\data_in_frame[7] [7]), .O(n23_adj_4250));
    defparam i7_4_lut_adj_1374.LUT_INIT = 16'hde7b;
    SB_LUT4 i11_4_lut_adj_1375 (.I0(n30259), .I1(n34602), .I2(n29843), 
            .I3(n5_adj_4029), .O(n27_adj_4251));
    defparam i11_4_lut_adj_1375.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_4_lut_adj_1376 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_825), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [7]), .O(n17589));
    defparam i1_2_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 select_413_Select_15_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4144));
    defparam select_413_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_16_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4142));
    defparam select_413_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i2_3_lut_4_lut_adj_1377 (.I0(n17364), .I1(n10_adj_4061), .I2(n32917), 
            .I3(n17814), .O(n30777));
    defparam i2_3_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [29]), .I3(GND_net), .O(n7_adj_4111));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'he0e0;
    SB_LUT4 select_413_Select_17_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4141));
    defparam select_413_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_18_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4140));
    defparam select_413_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i13_4_lut_adj_1379 (.I0(n17820), .I1(n26_adj_4249), .I2(n18_adj_4248), 
            .I3(n8_adj_4068), .O(n29_adj_4252));
    defparam i13_4_lut_adj_1379.LUT_INIT = 16'hfffe;
    SB_LUT4 select_413_Select_19_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4139));
    defparam select_413_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_20_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4138));
    defparam select_413_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n18216), .D(n8825[5]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_413_Select_21_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4137));
    defparam select_413_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_22_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4136));
    defparam select_413_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_23_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4134));
    defparam select_413_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i5_3_lut_4_lut_adj_1380 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[16] [6]), 
            .I2(n10_adj_4059), .I3(n32571), .O(n30854));
    defparam i5_3_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n18683));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1381 (.I0(\data_in_frame[14] [7]), .I1(n10_adj_4055), 
            .I2(n15471), .I3(n32794), .O(n32602));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_4_lut_adj_1381.LUT_INIT = 16'h9669;
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n18682));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n18681));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n18216), .D(n8825[4]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_1382 (.I0(n29_adj_4252), .I1(n27_adj_4251), .I2(n23_adj_4250), 
            .I3(n35002), .O(n31_adj_4238));
    defparam i15_4_lut_adj_1382.LUT_INIT = 16'hfeff;
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n18216), .D(n8825[3]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n18680));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1383 (.I0(\data_in_frame[8] [3]), .I1(n32487), 
            .I2(n10_adj_4054), .I3(\data_in_frame[10] [4]), .O(n32972));
    defparam i5_3_lut_4_lut_adj_1383.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(n29854), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n32571));
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n18216), .D(n8825[2]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_413_Select_24_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4132));
    defparam select_413_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i1_2_lut_3_lut_adj_1385 (.I0(n17370), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[12] [6]), .I3(GND_net), .O(n6_adj_4050));
    defparam i1_2_lut_3_lut_adj_1385.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n18216), .D(n8825[1]), .R(n20456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1386 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [30]), .I3(GND_net), .O(n7_adj_4110));
    defparam i1_2_lut_3_lut_adj_1386.LUT_INIT = 16'he0e0;
    SB_LUT4 add_43_32_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n27726), .O(n2_adj_4119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_32 (.CI(n27726), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n27727));
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n18679));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_413_Select_25_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4130));
    defparam select_413_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 add_43_31_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n27725), .O(n2_adj_4121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n27725), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n27726));
    SB_LUT4 select_413_Select_26_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4128));
    defparam select_413_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n18241), .D(n5065));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_413_Select_27_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4126));
    defparam select_413_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_28_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4124));
    defparam select_413_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n18678));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_31019 (.I0(byte_transmit_counter[1]), 
            .I1(n35892), .I2(n35893), .I3(byte_transmit_counter[2]), .O(n37382));
    defparam byte_transmit_counter_1__bdd_4_lut_31019.LUT_INIT = 16'he4aa;
    SB_LUT4 select_413_Select_29_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4122));
    defparam select_413_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_30_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4120));
    defparam select_413_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 select_413_Select_31_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4116));
    defparam select_413_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(n30259), .I1(\data_in_frame[8] [0]), 
            .I2(n17358), .I3(GND_net), .O(n6_adj_4049));
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'h9696;
    SB_LUT4 select_413_Select_0_i3_2_lut_4_lut (.I0(n2236), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17089), .I3(\FRAME_MATCHER.i [0]), .O(n3));
    defparam select_413_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'h5400;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(\data_in_frame[9] [4]), .I1(n29843), 
            .I2(n17814), .I3(GND_net), .O(n30005));
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1389 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[13] [4]), 
            .I2(n33033), .I3(\data_in_frame[11] [3]), .O(n17434));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_4_lut_adj_1389.LUT_INIT = 16'h6996;
    SB_LUT4 i14030_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n18819));
    defparam i14030_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(n8_adj_4068), .I1(\data_in_frame[9] [1]), 
            .I2(n17364), .I3(GND_net), .O(n17198));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(n10_adj_4061), .I1(n17814), .I2(\data_in_frame[9] [3]), 
            .I3(n32683), .O(n32933));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1392 (.I0(n17364), .I1(n10_adj_4061), .I2(Kp_23__N_1032), 
            .I3(n32650), .O(n33033));
    defparam i1_2_lut_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(\data_in_frame[8] [1]), .I1(n17391), 
            .I2(n15471), .I3(GND_net), .O(n15478));
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1394 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4254));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_1394.LUT_INIT = 16'h7bde;
    SB_LUT4 n37382_bdd_4_lut (.I0(n37382), .I1(n17_adj_4080), .I2(n16_adj_4079), 
            .I3(byte_transmit_counter[2]), .O(n37385));
    defparam n37382_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1395 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [3]), 
            .I2(n32714), .I3(GND_net), .O(n6_adj_4034));
    defparam i1_2_lut_3_lut_adj_1395.LUT_INIT = 16'h9696;
    SB_LUT4 i14031_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n18820));
    defparam i14031_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14032_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n18821));
    defparam i14032_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14033_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n18822));
    defparam i14033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14034_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n18823));
    defparam i14034_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n18677));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n18676));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n18675));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n18674));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n18673));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n18672));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n18671));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n18670));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n18669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n18668));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n18667));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n18666));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n18665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n18664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n18663));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n37934));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n37935));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n18241), .D(n5066));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1396 (.I0(n2_adj_4010), .I1(n1_adj_4188), 
            .I2(\FRAME_MATCHER.state [31]), .I3(GND_net), .O(n7_adj_4109));
    defparam i1_2_lut_3_lut_adj_1396.LUT_INIT = 16'he0e0;
    SB_LUT4 i14035_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n18824));
    defparam i14035_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n18241), .D(n5067));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n18241), .D(n5068));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n18241), .D(n5069));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n18241), .D(n5070));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n18241), .D(n5071));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n18241), .D(n5072));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n18241), .D(n5073));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n18241), 
            .D(n5074));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n18241), 
            .D(n5075));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n18241), 
            .D(n5076));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n18241), 
            .D(n5077));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n18241), 
            .D(n5078));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n18241), 
            .D(n5079));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n18241), 
            .D(n5080));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n18241), 
            .D(n5081));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n18241), 
            .D(n5082));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n18241), 
            .D(n5083));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n18241), 
            .D(n5084));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n18241), 
            .D(n5085));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n18241), 
            .D(n5086));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n18241), 
            .D(n5087));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_30_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n27724), .O(n2_adj_4123)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_30 (.CI(n27724), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n27725));
    SB_LUT4 i2_3_lut_4_lut_adj_1397 (.I0(n33978), .I1(n14278), .I2(n1_c), 
            .I3(n4_adj_4009), .O(n5_adj_4011));
    defparam i2_3_lut_4_lut_adj_1397.LUT_INIT = 16'hfff4;
    SB_LUT4 i14036_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n18825));
    defparam i14036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1398 (.I0(n33978), .I1(n14278), .I2(n1_adj_4188), 
            .I3(\FRAME_MATCHER.state [3]), .O(n31816));
    defparam i1_3_lut_4_lut_adj_1398.LUT_INIT = 16'hf400;
    SB_LUT4 i14037_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32391), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n18826));
    defparam i14037_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14022_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n18811));
    defparam i14022_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14023_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n18812));
    defparam i14023_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i2_4_lut_adj_1399 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4255));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_1399.LUT_INIT = 16'h7bde;
    SB_LUT4 i14024_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n18813));
    defparam i14024_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i3_4_lut_adj_1400 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4256));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_1400.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1401 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_1401.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1402 (.I0(n9), .I1(n11_adj_4256), .I2(n10_adj_4255), 
            .I3(n12_adj_4254), .O(n14565));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1402.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1403 (.I0(\FRAME_MATCHER.state[0] ), .I1(n14565), 
            .I2(GND_net), .I3(GND_net), .O(n32415));
    defparam i1_2_lut_adj_1403.LUT_INIT = 16'heeee;
    SB_LUT4 i14025_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n18814));
    defparam i14025_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14026_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n18815));
    defparam i14026_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14027_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n18816));
    defparam i14027_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14028_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n18817));
    defparam i14028_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14029_3_lut_4_lut (.I0(n10_adj_4239), .I1(n33579), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n18818));
    defparam i14029_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i14014_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n18803));
    defparam i14014_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14015_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n18804));
    defparam i14015_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14016_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n18805));
    defparam i14016_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14017_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n18806));
    defparam i14017_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3362_3_lut (.I0(n31_adj_4099), .I1(n31_adj_4238), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n14047));
    defparam i3362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14018_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n18807));
    defparam i14018_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14019_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n18808));
    defparam i14019_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14020_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n18809));
    defparam i14020_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1404 (.I0(n14047), .I1(n32415), .I2(n24690), 
            .I3(n24390), .O(n10_adj_4230));
    defparam i4_4_lut_adj_1404.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n6_adj_4006));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i14021_3_lut_4_lut (.I0(n8_adj_4104), .I1(n32406), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n18810));
    defparam i14021_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[2] [7]), .I3(GND_net), .O(n32505));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1407 (.I0(n30005), .I1(n29843), .I2(n17418), 
            .I3(\data_in_frame[11] [6]), .O(n32927));
    defparam i2_3_lut_4_lut_adj_1407.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_29_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n27723), .O(n2_adj_4125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_29 (.CI(n27723), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n27724));
    SB_LUT4 add_43_28_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n27722), .O(n2_adj_4127)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_28 (.CI(n27722), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n27723));
    SB_LUT4 i1_2_lut_4_lut_adj_1408 (.I0(\data_in_frame[9] [5]), .I1(n30005), 
            .I2(n29850), .I3(\data_in_frame[11] [6]), .O(n30884));
    defparam i1_2_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1409 (.I0(\FRAME_MATCHER.state [3]), .I1(n3482), 
            .I2(n5202), .I3(GND_net), .O(n34936));
    defparam i2_3_lut_adj_1409.LUT_INIT = 16'h0101;
    SB_LUT4 i1_4_lut_adj_1410 (.I0(n3482), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n17001), .I3(n5202), .O(n18470));
    defparam i1_4_lut_adj_1410.LUT_INIT = 16'h5011;
    SB_LUT4 i2_3_lut_4_lut_adj_1411 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[8] [0]), .I3(\data_out_frame[7] [6]), .O(n32999));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i13955_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n18744));
    defparam i13955_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i5_3_lut_4_lut_adj_1412 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[10] [3]), .I3(n32580), .O(n14_adj_4000));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_4_lut_adj_1412.LUT_INIT = 16'h6996;
    SB_LUT4 i13959_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n18748));
    defparam i13959_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13960_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n18749));
    defparam i13960_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13961_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n18750));
    defparam i13961_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13962_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n18751));
    defparam i13962_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13963_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n18752));
    defparam i13963_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13964_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n18753));
    defparam i13964_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 i13965_3_lut_4_lut (.I0(n10_adj_4190), .I1(n33579), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n18754));
    defparam i13965_3_lut_4_lut.LUT_INIT = 16'hfb40;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4257));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4258));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n19173));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n19172));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n19171));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n19170));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n19169));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n19168));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n19167));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n19166));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n19165));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n19164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n19163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n19162));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n19161));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n19160));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n19159));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n19158));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n19157));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n19156));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n19155));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n19154));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n19153));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n19152));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n19151));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n19118));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n19117));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n19116));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n19115));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n19114));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n19113));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n19112));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n19111));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n19110));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n19109));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n19108));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n19107));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n19106));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n19105));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n19104));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n19103));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n19102));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n19101));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n19100));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n19099));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n19098));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n19097));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n19096));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n19095));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n19094));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n19093));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n19092));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n19091));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n19090));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n19089));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n19088));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n19087));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n19086));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n19085));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n19084));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n19083));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n19082));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n19081));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n19080));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n19079));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n19078));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n19077));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n19076));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n19075));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n19074));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n19073));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n19072));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n19071));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n19070));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n19069));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n19068));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n19067));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n19066));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n19065));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n19064));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n19063));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n19062));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n19061));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n19060));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n19059));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n19058));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk32MHz), 
           .D(n19057));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk32MHz), 
           .D(n19056));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk32MHz), 
           .D(n19055));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk32MHz), 
           .D(n19054));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk32MHz), 
           .D(n19053));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk32MHz), 
           .D(n19052));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk32MHz), 
           .D(n19051));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk32MHz), 
           .D(n19050));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n19049));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n19048));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n19047));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n19046));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n19045));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n19044));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n19043));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n19042));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n19041));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n19040));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n19039));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n19038));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n19037));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n19036));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n19035));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n19034));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n19033));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n19032));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n19031));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n19030));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n19029));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n19028));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n19027));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n19026));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n19025));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n19024));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n19023));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n19022));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n19021));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n19020));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n19019));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n19018));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n19017));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n19016));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n19015));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n19014));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n19013));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n19012));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n19011));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n19010));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n19009));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n19008));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n19007));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n19006));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n19005));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n19004));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n19003));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n19002));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n19001));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n19000));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n18999));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n18998));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n18997));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n18996));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n18994));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n18993));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n18992));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n18991));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n18990));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n18989));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n18988));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n18987));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n18986));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n18985));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n18984));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n18983));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n18982));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30975 (.I0(byte_transmit_counter[1]), 
            .I1(n35927), .I2(n35928), .I3(byte_transmit_counter[2]), .O(n37376));
    defparam byte_transmit_counter_1__bdd_4_lut_30975.LUT_INIT = 16'he4aa;
    SB_LUT4 i13998_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n18787));
    defparam i13998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13999_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n18788));
    defparam i13999_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1413 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(n32546), .O(n32860));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 i14000_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n18789));
    defparam i14000_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14001_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n18790));
    defparam i14001_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14002_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n18791));
    defparam i14002_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1414 (.I0(\FRAME_MATCHER.state[0] ), .I1(n17068), 
            .I2(n3303), .I3(n14278), .O(n4_adj_4009));
    defparam i1_3_lut_4_lut_adj_1414.LUT_INIT = 16'h0200;
    SB_LUT4 i14003_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n18792));
    defparam i14003_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14004_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n18793));
    defparam i14004_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_27_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n27721), .O(n2_adj_4129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14005_3_lut_4_lut (.I0(n10_adj_4190), .I1(n32384), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n18794));
    defparam i14005_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18929_2_lut_3_lut (.I0(n63_adj_4057), .I1(n63_c), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n123));   // verilog/coms.v(227[6] 229[9])
    defparam i18929_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i28716_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n35112));
    defparam i28716_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i28714_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35110));
    defparam i28714_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut_adj_1415 (.I0(n63_adj_4057), .I1(n63_c), .I2(n63), 
            .I3(GND_net), .O(n14278));   // verilog/coms.v(227[6] 229[9])
    defparam i2_2_lut_3_lut_adj_1415.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut_4_lut_adj_1416 (.I0(\FRAME_MATCHER.state[0] ), .I1(n17089), 
            .I2(n771), .I3(n14278), .O(n1_c));
    defparam i1_3_lut_4_lut_adj_1416.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1417 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(n32391), .I3(\FRAME_MATCHER.i [0]), .O(n32395));
    defparam i1_2_lut_3_lut_4_lut_adj_1417.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_3_lut_4_lut_adj_1418 (.I0(\FRAME_MATCHER.state[0] ), .I1(n66), 
            .I2(n4452), .I3(n14278), .O(n1_adj_4188));
    defparam i1_3_lut_4_lut_adj_1418.LUT_INIT = 16'h0200;
    SB_CARRY add_43_27 (.CI(n27721), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n27722));
    SB_LUT4 add_43_26_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n27720), .O(n2_adj_4131)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_26 (.CI(n27720), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n27721));
    SB_LUT4 i2006851_i1_3_lut (.I0(n37535), .I1(n37433), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4247));
    defparam i2006851_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29817_2_lut (.I0(n37553), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35891));
    defparam i29817_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1419 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(n32398), .I3(\FRAME_MATCHER.i [0]), .O(n32400));
    defparam i1_2_lut_3_lut_4_lut_adj_1419.LUT_INIT = 16'hfeff;
    SB_LUT4 add_43_25_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n27719), .O(n2_adj_4133)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n18981));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1420 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(n32406), .I3(\FRAME_MATCHER.i [0]), .O(n32409));
    defparam i1_2_lut_3_lut_4_lut_adj_1420.LUT_INIT = 16'hfeff;
    SB_LUT4 i28707_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n35103));
    defparam i28707_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 equal_115_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4104));
    defparam equal_115_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i28705_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35101));
    defparam i28705_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(tx_transmit_N_3350), .I1(n23655), 
            .I2(\FRAME_MATCHER.i_31__N_2460 ), .I3(GND_net), .O(n32373));   // verilog/coms.v(214[11:56])
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'he0e0;
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n18980));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n18979));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n18978));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n18977));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2007454_i1_3_lut (.I0(n37511), .I1(n37517), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4246));
    defparam i2007454_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_4_lut_adj_1422 (.I0(tx_transmit_N_3350), .I1(n23655), 
            .I2(n14278), .I3(\FRAME_MATCHER.i_31__N_2460 ), .O(n2_adj_4010));   // verilog/coms.v(214[11:56])
    defparam i1_3_lut_4_lut_adj_1422.LUT_INIT = 16'he000;
    SB_LUT4 i29826_2_lut (.I0(n37565), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35912));
    defparam i29826_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_25 (.CI(n27719), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n27720));
    SB_LUT4 i1_2_lut_3_lut_adj_1423 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [2]), .I3(GND_net), .O(n17108));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1423.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1424 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[9] [1]), .I3(n32546), .O(n32894));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 n37376_bdd_4_lut (.I0(n37376), .I1(n17_adj_4259), .I2(n16_adj_4260), 
            .I3(byte_transmit_counter[2]), .O(n37379));
    defparam n37376_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1425 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[18] [5]), 
            .I2(n32699), .I3(n29938), .O(n30867));
    defparam i2_3_lut_4_lut_adj_1425.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n18976));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13971_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n18760));
    defparam i13971_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13972_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n18761));
    defparam i13972_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i28700_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35096));
    defparam i28700_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28701_4_lut (.I0(n35096), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35097));
    defparam i28701_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i28699_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35095));
    defparam i28699_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1426 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[23] [4]), 
            .I2(\data_out_frame[23] [5]), .I3(GND_net), .O(n32737));
    defparam i1_2_lut_3_lut_adj_1426.LUT_INIT = 16'h9696;
    SB_LUT4 i13973_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n18762));
    defparam i13973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2008057_i1_3_lut (.I0(n37505), .I1(n37559), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4244));
    defparam i2008057_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13966_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n18755));
    defparam i13966_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29860_2_lut (.I0(n37571), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35861));
    defparam i29860_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13967_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n18756));
    defparam i13967_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13968_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n18757));
    defparam i13968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4243));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4242));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29831_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35906));
    defparam i29831_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29833_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35905));
    defparam i29833_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n18975));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n18974));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13969_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n18758));
    defparam i13969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30970 (.I0(byte_transmit_counter[1]), 
            .I1(n35862), .I2(n35863), .I3(byte_transmit_counter[2]), .O(n37370));
    defparam byte_transmit_counter_1__bdd_4_lut_30970.LUT_INIT = 16'he4aa;
    SB_LUT4 i13970_3_lut_4_lut (.I0(n8_adj_4253), .I1(n32406), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n18759));
    defparam i13970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_24_lut (.I0(n2236), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n27718), .O(n2_adj_4135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13982_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n18771));
    defparam i13982_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n18973));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13983_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n18772));
    defparam i13983_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n18972));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n18971));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n18970));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n18969));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n18968));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n18967));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n18966));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n18965));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13984_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n18773));
    defparam i13984_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n18964));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n18963));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n18962));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n18961));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n18960));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n18959));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n18958));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n18957));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n18956));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n18955));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n18954));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n18953));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n18952));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n18951));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n18950));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n18949));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n18948));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n18640));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n18639));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n18638));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n18637));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n18636));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n18635));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n18634));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n18947));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n18946));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n18945));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n18944));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n18943));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n18942));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n18941));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n18940));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(\data_out_frame[5] [1]), .I1(n32872), 
            .I2(n18067), .I3(GND_net), .O(n33078));
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'h9696;
    SB_LUT4 i13985_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n18774));
    defparam i13985_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n18626));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n18939));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n18938));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n18937));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n18936));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n18935));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n18934));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n18933));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n18932));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n18931));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n18930));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n18929));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n18928));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n18927));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n18926));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n18925));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n18924));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n18923));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n18922));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n18921));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n18920));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n18919));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n18918));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n18917));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n18916));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n18915));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n18914));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n18913));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n18912));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n18911));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n18910));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n18909));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n18908));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n18907));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n18906));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n18905));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n18904));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n18903));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n18902));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n18901));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n18900));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n18899));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n18898));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n18897));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n18896));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13986_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n18775));
    defparam i13986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n18895));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n18894));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n18893));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n37370_bdd_4_lut (.I0(n37370), .I1(n17_adj_4258), .I2(n16_adj_4257), 
            .I3(byte_transmit_counter[2]), .O(n37373));
    defparam n37370_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13987_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n18776));
    defparam i13987_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13988_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n18777));
    defparam i13988_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13989_3_lut_4_lut (.I0(n8), .I1(n32406), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n18778));
    defparam i13989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_24 (.CI(n27718), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n27719));
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n18892));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n18891));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1428 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n32580));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1428.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n18890));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n18889));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1429 (.I0(\data_out_frame[5] [1]), .I1(n32872), 
            .I2(\data_out_frame[9] [4]), .I3(GND_net), .O(n32561));
    defparam i1_2_lut_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n18888));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n18887));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n18886));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1430 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [2]), .I3(n32608), .O(n17678));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n18885));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n18884));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n18883));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1431 (.I0(n24219), .I1(n10_adj_4239), .I2(GND_net), 
            .I3(GND_net), .O(n32391));
    defparam i1_2_lut_adj_1431.LUT_INIT = 16'hdddd;
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n18882));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_3_lut_adj_1432 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(GND_net), .O(n10_adj_3998));   // verilog/coms.v(85[17:63])
    defparam i2_2_lut_3_lut_adj_1432.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n18881));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n18880));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n18879));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n18878));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n18877));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n18876));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n18875));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n18874));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n18873));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n18872));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n18871));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n18870));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n18869));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n18868));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n18867));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n18866));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n18865));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n18864));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n18863));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n18862));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n18861));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n18860));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n18859));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n18858));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n18857));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n18856));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n18855));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n18854));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n18853));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n18852));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n18851));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n18850));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n18849));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n18848));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n18847));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n18846));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n18845));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n18844));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n18843));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2051_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n8_adj_4221));
    defparam i2051_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n18842));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n18841));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n18840));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n18839));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n18838));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n18837));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n18836));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n18835));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28677_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n35073));
    defparam i28677_4_lut.LUT_INIT = 16'hec2c;
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n18834));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n18833));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n18832));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n18831));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n18830));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n18829));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n18828));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n18827));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n18826));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n18825));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n18824));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n18823));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28675_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35071));
    defparam i28675_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n18822));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1433 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n24219), .O(n33579));
    defparam i2_3_lut_4_lut_adj_1433.LUT_INIT = 16'h8000;
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n18821));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_117_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4253));
    defparam equal_117_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n18820));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1434 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[5] [1]), .I3(GND_net), .O(n32438));
    defparam i1_2_lut_3_lut_adj_1434.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n18819));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n18818));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_132_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4239));   // verilog/coms.v(154[7:23])
    defparam equal_132_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n18817));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n18816));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n18815));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n18814));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n18813));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n18812));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n18811));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n18810));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n18809));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n18808));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n18807));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n18806));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n18805));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n18804));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n18803));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n18802));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n18801));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_124_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4190));   // verilog/coms.v(154[7:23])
    defparam equal_124_i10_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n18800));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n18799));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n18798));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1435 (.I0(n16700), .I1(\data_out_frame[14] [2]), 
            .I2(\data_out_frame[14] [1]), .I3(n29949), .O(n29953));
    defparam i2_3_lut_4_lut_adj_1435.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n18797));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2010469_i1_3_lut (.I0(n37457), .I1(n37451), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4241));
    defparam i2010469_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n18796));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n18795));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n18794));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29835_2_lut (.I0(n37601), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35904));
    defparam i29835_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n18793));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n18792));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1436 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state_31__N_2561 [3]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n6_adj_4192));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1436.LUT_INIT = 16'h00bf;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1437 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n24776), .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n77));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1437.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1438 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n24776), .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n66));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1438.LUT_INIT = 16'hfeff;
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n18791));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n18790));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n18789));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1439 (.I0(\data_out_frame[9] [3]), .I1(n1168), 
            .I2(\data_out_frame[4] [7]), .I3(GND_net), .O(n32428));
    defparam i1_2_lut_3_lut_adj_1439.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1440 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n24776), .I2(n74), .I3(\FRAME_MATCHER.state [1]), .O(\FRAME_MATCHER.i_31__N_2460 ));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1440.LUT_INIT = 16'h1000;
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n18788));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n18787));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n18786));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1441 (.I0(\FRAME_MATCHER.state [3]), 
            .I1(n24776), .I2(\FRAME_MATCHER.state[0] ), .I3(\FRAME_MATCHER.state [1]), 
            .O(n17092));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_4_lut_adj_1441.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1442 (.I0(\FRAME_MATCHER.state [3]), .I1(n24776), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n17068));   // verilog/coms.v(212[5:16])
    defparam i2_3_lut_4_lut_adj_1442.LUT_INIT = 16'hffef;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30965 (.I0(byte_transmit_counter[1]), 
            .I1(n35908), .I2(n35909), .I3(byte_transmit_counter[2]), .O(n37364));
    defparam byte_transmit_counter_1__bdd_4_lut_30965.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1443 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[8] [1]), .O(n6_adj_3988));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n18785));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n18784));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1444 (.I0(\data_out_frame[25] [6]), .I1(n30912), 
            .I2(n29938), .I3(\data_out_frame[23] [4]), .O(n32975));
    defparam i1_2_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n18783));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[18] [4]), 
            .I2(n32831), .I3(n30803), .O(n15336));
    defparam i2_3_lut_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1446 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [5]), 
            .I2(n32561), .I3(n32805), .O(n32939));
    defparam i2_3_lut_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1447 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[11] [5]), .I3(n10_adj_3989), .O(n29949));
    defparam i5_3_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n18782));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n18781));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n18780));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1448 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[16] [4]), 
            .I2(n33517), .I3(GND_net), .O(n32831));
    defparam i1_2_lut_3_lut_adj_1448.LUT_INIT = 16'h6969;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n18779));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n18778));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n18777));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28673_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35069));
    defparam i28673_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n18776));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n18775));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n18774));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n18773));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n18772));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28674_4_lut (.I0(n35069), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35070));
    defparam i28674_4_lut.LUT_INIT = 16'ha3a0;
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n18771));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1449 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n6_adj_4017));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1449.LUT_INIT = 16'h9696;
    SB_LUT4 i28672_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35068));
    defparam i28672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n17466));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1451 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[5] [1]), 
            .I2(n32872), .I3(n18067), .O(n32802));
    defparam i1_2_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1452 (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[11] [6]), .I3(GND_net), .O(n10_adj_3993));
    defparam i2_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1453 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[4] [6]), .O(n18067));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n18770));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n18769));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2012278_i1_3_lut (.I0(n37529), .I1(n37523), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4240));
    defparam i2012278_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n18768));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1454 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[4] [5]), .I3(\data_out_frame[6] [7]), .O(n32596));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1455 (.I0(n30867), .I1(\data_out_frame[25] [4]), 
            .I2(n32825), .I3(n29938), .O(n6_adj_3986));
    defparam i1_2_lut_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 n37364_bdd_4_lut (.I0(n37364), .I1(n17_adj_4181), .I2(n16_adj_4180), 
            .I3(byte_transmit_counter[2]), .O(n37367));
    defparam n37364_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i29832_2_lut (.I0(n37331), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35907));
    defparam i29832_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_4_lut_adj_1456 (.I0(\data_out_frame[6] [6]), .I1(n1130), 
            .I2(n32596), .I3(n17610), .O(n32854));
    defparam i2_2_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i29845_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35863));
    defparam i29845_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29847_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35862));
    defparam i29847_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_4_lut_adj_1457 (.I0(\data_out_frame[6] [6]), .I1(n1130), 
            .I2(n32596), .I3(\data_out_frame[9] [2]), .O(n17886));
    defparam i2_2_lut_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n18767));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n18766));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1458 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[16] [5]), 
            .I2(n29969), .I3(GND_net), .O(n29979));
    defparam i1_2_lut_3_lut_adj_1458.LUT_INIT = 16'h9696;
    SB_LUT4 i13_3_lut_4_lut (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [7]), 
            .I2(n17711), .I3(n32529), .O(n38));
    defparam i13_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30960 (.I0(byte_transmit_counter[1]), 
            .I1(n35868), .I2(n35869), .I3(byte_transmit_counter[2]), .O(n37358));
    defparam byte_transmit_counter_1__bdd_4_lut_30960.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_4_lut_adj_1459 (.I0(n16700), .I1(n32746), .I2(n29949), 
            .I3(\data_out_frame[18] [3]), .O(n6_adj_3985));
    defparam i1_2_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n18765));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n37358_bdd_4_lut (.I0(n37358), .I1(n17_adj_4179), .I2(n16_adj_4178), 
            .I3(byte_transmit_counter[2]), .O(n37361));
    defparam n37358_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n18764));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n18763));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n18762));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1460 (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[14] [1]), .I3(n10_adj_3987), .O(n30803));
    defparam i5_3_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n18761));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1461 (.I0(n2394), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[25] [1]), .I3(n29929), .O(n34574));
    defparam i2_3_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n18760));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4260));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4259));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1462 (.I0(n2394), .I1(\data_out_frame[25] [2]), 
            .I2(n32825), .I3(GND_net), .O(n32826));
    defparam i1_2_lut_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30955 (.I0(byte_transmit_counter[1]), 
            .I1(n35902), .I2(n35903), .I3(byte_transmit_counter[2]), .O(n37352));
    defparam byte_transmit_counter_1__bdd_4_lut_30955.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1463 (.I0(\data_out_frame[20] [4]), .I1(n33521), 
            .I2(n10_adj_3982), .I3(\data_out_frame[23] [1]), .O(n2394));
    defparam i5_3_lut_4_lut_adj_1463.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1464 (.I0(\data_out_frame[4] [7]), .I1(n32438), 
            .I2(n32885), .I3(GND_net), .O(n16793));
    defparam i1_2_lut_3_lut_adj_1464.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1465 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[11] [6]), 
            .I2(\data_out_frame[14] [0]), .I3(GND_net), .O(n32690));
    defparam i1_2_lut_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 n37352_bdd_4_lut (.I0(n37352), .I1(n17_adj_4177), .I2(n16_adj_4176), 
            .I3(byte_transmit_counter[2]), .O(n36443));
    defparam n37352_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_3_lut_4_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [7]), .I3(n17731), .O(n24));   // verilog/coms.v(77[16:27])
    defparam i7_3_lut_4_lut.LUT_INIT = 16'h0096;
    SB_LUT4 i2_3_lut_4_lut_adj_1466 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [0]), .I3(Kp_23__N_825), .O(n17926));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1467 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n15437));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1467.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1468 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(76[16:27])
    defparam i2_2_lut_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30950 (.I0(byte_transmit_counter[1]), 
            .I1(n35874), .I2(n35875), .I3(byte_transmit_counter[2]), .O(n37346));
    defparam byte_transmit_counter_1__bdd_4_lut_30950.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_4_lut_adj_1469 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(\data_out_frame[8] [6]), .O(n18108));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[20] [3]), 
            .I2(n34478), .I3(GND_net), .O(n30836));
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i28694_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35090));
    defparam i28694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28695_4_lut (.I0(n35090), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35091));
    defparam i28695_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i28693_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35089));
    defparam i28693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1471 (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n33030));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i2008660_i1_3_lut (.I0(n37499), .I1(n37391), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4236));
    defparam i2008660_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29846_2_lut (.I0(n37577), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35864));
    defparam i29846_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1472 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(n32529), .I3(GND_net), .O(n30019));
    defparam i1_2_lut_3_lut_adj_1472.LUT_INIT = 16'h9696;
    SB_LUT4 i28688_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35084));
    defparam i28688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut_4_lut_adj_1473 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[2] [5]), .O(n32877));   // verilog/coms.v(76[16:27])
    defparam i2_2_lut_3_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i28689_4_lut (.I0(n35084), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n35085));
    defparam i28689_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i28687_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n35083));
    defparam i28687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut_adj_1474 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[16] [0]), 
            .I2(n10_adj_3980), .I3(n32923), .O(n32981));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1475 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[17] [4]), 
            .I2(n17207), .I3(\data_out_frame[15] [4]), .O(n32674));
    defparam i2_3_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1476 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n17664));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1476.LUT_INIT = 16'h9696;
    SB_LUT4 i2009263_i1_3_lut (.I0(n37493), .I1(n37409), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4235));
    defparam i2009263_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29843_2_lut (.I0(n37583), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n35870));
    defparam i29843_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 n37346_bdd_4_lut (.I0(n37346), .I1(n17_adj_4175), .I2(n16_adj_4174), 
            .I3(byte_transmit_counter[2]), .O(n37349));
    defparam n37346_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1477 (.I0(n17693), .I1(n30019), .I2(\data_out_frame[17] [5]), 
            .I3(GND_net), .O(n30895));
    defparam i1_2_lut_3_lut_adj_1477.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut_adj_1478 (.I0(\data_out_frame[15] [4]), .I1(n17534), 
            .I2(n32511), .I3(\data_out_frame[19] [7]), .O(n6_adj_3970));   // verilog/coms.v(71[16:27])
    defparam i2_2_lut_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1479 (.I0(n17534), .I1(\data_out_frame[15] [3]), 
            .I2(\data_out_frame[15] [2]), .I3(n29940), .O(n29942));
    defparam i2_3_lut_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i29848_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35928));
    defparam i29848_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29788_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n35927));
    defparam i29788_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1480 (.I0(\data_out_frame[23] [6]), .I1(n17693), 
            .I2(n32664), .I3(GND_net), .O(n32978));
    defparam i1_2_lut_3_lut_adj_1480.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1481 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(n24219), .O(n32384));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1481.LUT_INIT = 16'hfdff;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30980 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n37328));
    defparam byte_transmit_counter_0__bdd_4_lut_30980.LUT_INIT = 16'he4aa;
    SB_LUT4 n37328_bdd_4_lut (.I0(n37328), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n37331));
    defparam n37328_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1482 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32391), .I3(\FRAME_MATCHER.i [0]), .O(n32394));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1482.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1483 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32406), .I3(\FRAME_MATCHER.i [0]), .O(n32410));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1483.LUT_INIT = 16'hfdff;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30985 (.I0(byte_transmit_counter[3]), 
            .I1(n36443), .I2(n35901), .I3(byte_transmit_counter[4]), .O(n37322));
    defparam byte_transmit_counter_3__bdd_4_lut_30985.LUT_INIT = 16'he4aa;
    SB_LUT4 n37322_bdd_4_lut (.I0(n37322), .I1(n14_adj_4173), .I2(n7_adj_4202), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n37322_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1484 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n32398), .I3(\FRAME_MATCHER.i [0]), .O(n32402));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1484.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_4_lut_adj_1485 (.I0(n16652), .I1(n32900), .I2(\data_out_frame[20] [2]), 
            .I3(n32778), .O(n2332));
    defparam i1_2_lut_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1486 (.I0(n16767), .I1(n30832), .I2(n32837), 
            .I3(n29929), .O(n33844));
    defparam i2_3_lut_4_lut_adj_1486.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1487 (.I0(\data_in_frame[6] [5]), .I1(n10), 
            .I2(\data_in_frame[4] [4]), .I3(\data_in_frame[4] [3]), .O(n17376));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1488 (.I0(n16767), .I1(n30832), .I2(n32837), 
            .I3(n33385), .O(n33843));
    defparam i2_3_lut_4_lut_adj_1488.LUT_INIT = 16'h9669;
    SB_LUT4 i13915_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n18704));
    defparam i13915_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1489 (.I0(\FRAME_MATCHER.state_31__N_2561 [3]), .I1(n32378), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n14410));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_adj_1489.LUT_INIT = 16'h8080;
    SB_LUT4 i13916_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n18705));
    defparam i13916_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13917_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n18706));
    defparam i13917_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13918_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n18707));
    defparam i13918_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1490 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [4]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n24219), .O(n32398));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_4_lut_adj_1490.LUT_INIT = 16'hfbff;
    SB_LUT4 i13919_3_lut_4_lut (.I0(n8), .I1(n32398), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n18708));
    defparam i13919_3_lut_4_lut.LUT_INIT = 16'hfe10;
    uart_tx tx (.clk32MHz(clk32MHz), .\r_SM_Main_2__N_3453[0] (r_SM_Main_2__N_3453[0]), 
            .r_SM_Main({r_SM_Main}), .n10125(n10125), .GND_net(GND_net), 
            .tx_o(tx_o), .tx_data({tx_data}), .\r_SM_Main_2__N_3450[1] (\r_SM_Main_2__N_3450[1] ), 
            .\r_Bit_Index[0] (\r_Bit_Index[0] ), .n18336(n18336), .n18590(n18590), 
            .VCC_net(VCC_net), .n4(n4), .n18644(n18644), .tx_active(tx_active), 
            .n18660(n18660), .n37939(n37939), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n23776(n23776), .GND_net(GND_net), 
            .n4(n4_adj_3), .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_4 ), .n17079(n17079), 
            .n4_adj_1(n4_adj_5), .r_SM_Main({r_SM_Main_adj_10}), .\r_SM_Main_2__N_3379[2] (\r_SM_Main_2__N_3379[2] ), 
            .n17084(n17084), .n4_adj_2(n4_adj_9), .n31970(n31970), .VCC_net(VCC_net), 
            .rx_data_ready(rx_data_ready), .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), 
            .n33211(n33211), .n33251(n33251), .n19204(n19204), .rx_data({rx_data}), 
            .n19202(n19202), .n19201(n19201), .n19200(n19200), .n19199(n19199), 
            .n19198(n19198), .n19197(n19197), .n18696(n18696), .n18995(n18995), 
            .n32359(n32359)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk32MHz, \r_SM_Main_2__N_3453[0] , r_SM_Main, n10125, 
            GND_net, tx_o, tx_data, \r_SM_Main_2__N_3450[1] , \r_Bit_Index[0] , 
            n18336, n18590, VCC_net, n4, n18644, tx_active, n18660, 
            n37939, tx_enable) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    input \r_SM_Main_2__N_3453[0] ;
    output [2:0]r_SM_Main;
    output n10125;
    input GND_net;
    output tx_o;
    input [7:0]tx_data;
    output \r_SM_Main_2__N_3450[1] ;
    output \r_Bit_Index[0] ;
    output n18336;
    output n18590;
    input VCC_net;
    output n4;
    input n18644;
    output tx_active;
    input n18660;
    input n37939;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n18554, n3, n14341;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n12041, n3_adj_3967;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]n307;
    
    wire n24310, n12040, n37547, n37421, o_Tx_Serial_N_3481, n28465, 
        n28464, n28463, n28462, n28461, n28460, n28459, n28458, 
        n10, n33444, n37544, n37418;
    
    SB_DFFESR r_Clock_Count_1549__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n1), .D(n41[0]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n1), .D(n41[8]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n1), .D(n41[7]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n1), .D(n41[6]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n1), .D(n41[5]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n1), .D(n41[4]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n1), .D(n41[3]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n1), .D(n41[2]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1549__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n1), .D(n41[1]), .R(n18554));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i5429_2_lut (.I0(\r_SM_Main_2__N_3453[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n10125));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5429_2_lut.LUT_INIT = 16'h2222;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n12041), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i9379_2_lut_3_lut (.I0(\r_SM_Main_2__N_3450[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_3967));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i9379_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i1645_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1645_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13801_3_lut (.I0(n18336), .I1(n24310), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n18590));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13801_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1652_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1652_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n24310));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i7335_4_lut (.I0(\r_SM_Main_2__N_3453[0] ), .I1(n24310), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3450[1] ), .O(n12040));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7335_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7336_3_lut (.I0(n12040), .I1(\r_SM_Main_2__N_3450[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n12041));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7336_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2011072_i1_3_lut (.I0(n37547), .I1(n37421), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3481));
    defparam i2011072_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3481), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 r_Clock_Count_1549_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n28465), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1549_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n28464), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_9 (.CI(n28464), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n28465));
    SB_LUT4 r_Clock_Count_1549_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n28463), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_8 (.CI(n28463), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n28464));
    SB_LUT4 r_Clock_Count_1549_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n28462), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_7 (.CI(n28462), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n28463));
    SB_LUT4 r_Clock_Count_1549_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n28461), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_6 (.CI(n28461), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n28462));
    SB_LUT4 r_Clock_Count_1549_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n28460), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_5 (.CI(n28460), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n28461));
    SB_LUT4 r_Clock_Count_1549_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n28459), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_4 (.CI(n28459), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n28460));
    SB_LUT4 r_Clock_Count_1549_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n28458), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_3 (.CI(n28458), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n28459));
    SB_LUT4 r_Clock_Count_1549_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1549_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1549_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n28458));
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[3]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n33444));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n33444), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3450[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30403_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3450[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n18554));
    defparam i30403_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n37544));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n37544_bdd_4_lut (.I0(n37544), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n37547));
    defparam n37544_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3450[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_31109 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n37418));
    defparam r_Bit_Index_0__bdd_4_lut_31109.LUT_INIT = 16'he4aa;
    SB_LUT4 n37418_bdd_4_lut (.I0(n37418), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n37421));
    defparam n37418_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n18336), 
            .D(n307[2]), .R(n18590));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n18336), 
            .D(n307[1]), .R(n18590));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n14341), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3967), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n18644));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n18660));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n37939));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3450[1] ), .O(n18336));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3453[0] ), 
            .I3(r_SM_Main[1]), .O(n14341));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n23776, GND_net, n4, \r_Bit_Index[0] , n17079, 
            n4_adj_1, r_SM_Main, \r_SM_Main_2__N_3379[2] , n17084, n4_adj_2, 
            n31970, VCC_net, rx_data_ready, r_Rx_Data, RX_N_10, n33211, 
            n33251, n19204, rx_data, n19202, n19201, n19200, n19199, 
            n19198, n19197, n18696, n18995, n32359) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output n23776;
    input GND_net;
    output n4;
    output \r_Bit_Index[0] ;
    output n17079;
    output n4_adj_1;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3379[2] ;
    output n17084;
    output n4_adj_2;
    input n31970;
    input VCC_net;
    output rx_data_ready;
    output r_Rx_Data;
    input RX_N_10;
    output n33211;
    output n33251;
    input n19204;
    output [7:0]rx_data;
    input n19202;
    input n19201;
    input n19200;
    input n19199;
    input n19198;
    input n19197;
    input n18696;
    input n18995;
    input n32359;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]n37;
    
    wire n18287;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n18556;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n16882;
    wire [2:0]n326;
    
    wire n21633, r_Rx_Data_R, n24274, n22, n21627, n3, n28472, 
        n28471, n28470, n28469, n28468, n28467, n28466, n21619, 
        n24460, n21632, n31, n5, n8, n6;
    
    SB_DFFESR r_Clock_Count_1547__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n18287), .D(n37[7]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1547__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n18287), .D(n37[6]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1547__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n18287), .D(n37[5]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1547__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n18287), .D(n37[4]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1547__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n18287), .D(n37[3]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1547__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n18287), .D(n37[2]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1547__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n18287), .D(n37[0]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1547__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n18287), .D(n37[1]), .R(n18556));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i19004_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n23776));
    defparam i19004_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_143_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_143_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut (.I0(\r_Bit_Index[0] ), .I1(n16882), .I2(GND_net), 
            .I3(GND_net), .O(n17079));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_144_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_144_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3379[2] ), .O(n16882));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i3_4_lut.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_adj_836 (.I0(n16882), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n17084));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_836.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_146_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_146_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1623_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1623_2_lut.LUT_INIT = 16'h6666;
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n31970));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n21633), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 i30579_3_lut (.I0(n33211), .I1(n24274), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n33251));
    defparam i30579_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i30900_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3379[2] ), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main[1]), .O(n33211));
    defparam i30900_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1630_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1630_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1_2_lut_adj_837 (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3379[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n22));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_837.LUT_INIT = 16'h8888;
    SB_LUT4 i16850_4_lut (.I0(r_Rx_Data), .I1(n22), .I2(r_SM_Main[1]), 
            .I3(n21627), .O(n3));   // verilog/uart_rx.v(36[17:26])
    defparam i16850_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 r_Clock_Count_1547_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n28472), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1547_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n28471), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1547_add_4_8 (.CI(n28471), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n28472));
    SB_LUT4 r_Clock_Count_1547_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n28470), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1547_add_4_7 (.CI(n28470), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n28471));
    SB_LUT4 r_Clock_Count_1547_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n28469), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1547_add_4_6 (.CI(n28469), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n28470));
    SB_LUT4 r_Clock_Count_1547_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n28468), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1547_add_4_5 (.CI(n28468), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n28469));
    SB_LUT4 r_Clock_Count_1547_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n28467), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1547_add_4_4 (.CI(n28467), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n28468));
    SB_LUT4 r_Clock_Count_1547_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n28466), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1547_add_4_3 (.CI(n28466), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n28467));
    SB_LUT4 r_Clock_Count_1547_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1547_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1547_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n28466));
    SB_LUT4 i1_2_lut_adj_838 (.I0(r_SM_Main[0]), .I1(n21619), .I2(GND_net), 
            .I3(GND_net), .O(n21627));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_838.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n24274));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n24274), .I1(\r_SM_Main_2__N_3379[2] ), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n24460));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i16854_3_lut (.I0(n21632), .I1(n24460), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n21633));   // verilog/uart_rx.v(36[17:26])
    defparam i16854_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i16853_3_lut_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n21619), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n21632));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i16853_3_lut_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_LUT4 i3_4_lut_adj_839 (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[5]), 
            .I2(n31), .I3(n5), .O(n21619));
    defparam i3_4_lut_adj_839.LUT_INIT = 16'hfdff;
    SB_LUT4 i3_4_lut_adj_840 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[0]), 
            .I2(r_Clock_Count[4]), .I3(r_Clock_Count[3]), .O(n5));
    defparam i3_4_lut_adj_840.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_841 (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(GND_net), .I3(GND_net), .O(n31));   // verilog/uart_rx.v(120[34:51])
    defparam i1_2_lut_adj_841.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(n31), .I1(n5), .I2(r_Clock_Count[2]), .I3(r_Clock_Count[5]), 
            .O(\r_SM_Main_2__N_3379[2] ));
    defparam i1_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i13767_3_lut (.I0(n18287), .I1(r_SM_Main[2]), .I2(n8), .I3(GND_net), 
            .O(n18556));   // verilog/uart_rx.v(120[34:51])
    defparam i13767_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_2_lut (.I0(n21619), .I1(r_SM_Main[0]), .I2(GND_net), .I3(GND_net), 
            .O(n6));   // verilog/uart_rx.v(36[17:26])
    defparam i2_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_842 (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n6), 
            .I3(r_Rx_Data), .O(n18287));   // verilog/uart_rx.v(36[17:26])
    defparam i1_4_lut_adj_842.LUT_INIT = 16'h3233;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n33211), 
            .D(n326[2]), .R(n33251));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n33211), 
            .D(n326[1]), .R(n33251));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i19_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n21619), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3379[2] ), .O(n8));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i19_3_lut_4_lut.LUT_INIT = 16'h08f8;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n19204));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n19202));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n19201));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n19200));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n19199));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n19198));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n19197));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n18696));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n18995));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(\r_SM_Main_2__N_3379[2] ), 
            .R(n32359));   // verilog/uart_rx.v(49[10] 144[8])
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n36611, VCC_net, INHA_c, clk32MHz, n16908, pwm_counter, 
            n16906, GND_net) /* synthesis syn_module_defined=1 */ ;
    input n36611;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n16908;
    output [31:0]pwm_counter;
    input n16906;
    input GND_net;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n14, n13, n4, n33831, n8, n12, pwm_counter_31__N_648;
    wire [31:0]n133;
    
    wire n28503, n28502, n28501, n28500, n28499, n28498, n28497, 
        n28496, n28495, n28494, n28493, n28492, n28491, n28490, 
        n28489, n28488, n28487, n28486, n28485, n28484, n28483, 
        n28482, n28481, n28480, n28479, n28478, n28477, n28476, 
        n28475, n28474, n28473;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n36611), 
            .R(n16908));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i6_4_lut (.I0(pwm_counter[15]), .I1(pwm_counter[14]), .I2(pwm_counter[17]), 
            .I3(pwm_counter[22]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(pwm_counter[16]), .I1(pwm_counter[19]), .I2(n16906), 
            .I3(pwm_counter[18]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(pwm_counter[8]), .I1(pwm_counter[7]), .I2(GND_net), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut (.I0(pwm_counter[6]), .I1(pwm_counter[10]), .I2(n4), 
            .I3(pwm_counter[9]), .O(n33831));
    defparam i2_4_lut.LUT_INIT = 16'hc800;
    SB_LUT4 i1_3_lut (.I0(pwm_counter[21]), .I1(n13), .I2(n14), .I3(GND_net), 
            .O(n8));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_835 (.I0(pwm_counter[12]), .I1(pwm_counter[11]), 
            .I2(n33831), .I3(pwm_counter[20]), .O(n12));
    defparam i5_4_lut_adj_835.LUT_INIT = 16'hfffe;
    SB_LUT4 i19013_4_lut (.I0(pwm_counter[13]), .I1(pwm_counter[31]), .I2(n12), 
            .I3(n8), .O(pwm_counter_31__N_648));   // verilog/pwm.v(18[8:40])
    defparam i19013_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 pwm_counter_1545_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[31]), 
            .I3(n28503), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1545_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n28502), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_32 (.CI(n28502), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n28503));
    SB_LUT4 pwm_counter_1545_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n28501), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_31 (.CI(n28501), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n28502));
    SB_LUT4 pwm_counter_1545_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n28500), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_30 (.CI(n28500), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n28501));
    SB_LUT4 pwm_counter_1545_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n28499), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_29 (.CI(n28499), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n28500));
    SB_LUT4 pwm_counter_1545_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n28498), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_28 (.CI(n28498), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n28499));
    SB_LUT4 pwm_counter_1545_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n28497), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_27 (.CI(n28497), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n28498));
    SB_LUT4 pwm_counter_1545_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n28496), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_26 (.CI(n28496), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n28497));
    SB_LUT4 pwm_counter_1545_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n28495), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_25 (.CI(n28495), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n28496));
    SB_LUT4 pwm_counter_1545_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n28494), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_24 (.CI(n28494), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n28495));
    SB_LUT4 pwm_counter_1545_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n28493), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_23 (.CI(n28493), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n28494));
    SB_LUT4 pwm_counter_1545_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n28492), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_22 (.CI(n28492), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n28493));
    SB_LUT4 pwm_counter_1545_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n28491), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_21 (.CI(n28491), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n28492));
    SB_LUT4 pwm_counter_1545_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n28490), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_20 (.CI(n28490), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n28491));
    SB_LUT4 pwm_counter_1545_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n28489), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_19 (.CI(n28489), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n28490));
    SB_LUT4 pwm_counter_1545_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n28488), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_18 (.CI(n28488), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n28489));
    SB_LUT4 pwm_counter_1545_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n28487), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_17 (.CI(n28487), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n28488));
    SB_LUT4 pwm_counter_1545_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n28486), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_16 (.CI(n28486), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n28487));
    SB_LUT4 pwm_counter_1545_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n28485), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_15 (.CI(n28485), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n28486));
    SB_LUT4 pwm_counter_1545_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n28484), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_14 (.CI(n28484), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n28485));
    SB_LUT4 pwm_counter_1545_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n28483), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_13 (.CI(n28483), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n28484));
    SB_LUT4 pwm_counter_1545_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n28482), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_12 (.CI(n28482), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n28483));
    SB_LUT4 pwm_counter_1545_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n28481), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_11 (.CI(n28481), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n28482));
    SB_LUT4 pwm_counter_1545_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n28480), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_10 (.CI(n28480), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n28481));
    SB_LUT4 pwm_counter_1545_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n28479), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_9 (.CI(n28479), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n28480));
    SB_LUT4 pwm_counter_1545_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n28478), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_8 (.CI(n28478), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n28479));
    SB_LUT4 pwm_counter_1545_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n28477), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_7 (.CI(n28477), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n28478));
    SB_LUT4 pwm_counter_1545_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n28476), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_6 (.CI(n28476), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n28477));
    SB_LUT4 pwm_counter_1545_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n28475), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_5 (.CI(n28475), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n28476));
    SB_LUT4 pwm_counter_1545_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n28474), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_4 (.CI(n28474), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n28475));
    SB_LUT4 pwm_counter_1545_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n28473), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_3 (.CI(n28473), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n28474));
    SB_LUT4 pwm_counter_1545_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1545_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1545_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n28473));
    SB_DFFSR pwm_counter_1545__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n133[10]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n133[11]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n133[12]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n133[13]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n133[14]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n133[15]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n133[16]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n133[17]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n133[18]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n133[19]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n133[20]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n133[21]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n133[22]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1545__i31 (.Q(pwm_counter[31]), .C(clk32MHz), .D(n133[31]), 
            .R(pwm_counter_31__N_648));   // verilog/pwm.v(17[20:33])
    
endmodule
